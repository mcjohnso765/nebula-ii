* NGSPICE file created from team_09.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_1 abstract view
.subckt sky130_fd_sc_hd__o221ai_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_1 abstract view
.subckt sky130_fd_sc_hd__a311oi_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_8 abstract view
.subckt sky130_fd_sc_hd__inv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_8 abstract view
.subckt sky130_fd_sc_hd__clkinv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__bufinv_16 abstract view
.subckt sky130_fd_sc_hd__bufinv_16 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_1 abstract view
.subckt sky130_fd_sc_hd__o2111ai_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_4 abstract view
.subckt sky130_fd_sc_hd__a21boi_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_2 abstract view
.subckt sky130_fd_sc_hd__o21ba_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_1 abstract view
.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_2 abstract view
.subckt sky130_fd_sc_hd__nand4b_2 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_16 abstract view
.subckt sky130_fd_sc_hd__inv_16 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_12 abstract view
.subckt sky130_fd_sc_hd__inv_12 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_4 abstract view
.subckt sky130_fd_sc_hd__o21bai_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_2 abstract view
.subckt sky130_fd_sc_hd__or4bb_2 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_2 abstract view
.subckt sky130_fd_sc_hd__o311a_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_4 abstract view
.subckt sky130_fd_sc_hd__a2111o_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinvlp_4 abstract view
.subckt sky130_fd_sc_hd__clkinvlp_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_4 abstract view
.subckt sky130_fd_sc_hd__o22ai_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_4 abstract view
.subckt sky130_fd_sc_hd__o31a_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_4 abstract view
.subckt sky130_fd_sc_hd__o221ai_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_4 abstract view
.subckt sky130_fd_sc_hd__or4bb_4 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_1 abstract view
.subckt sky130_fd_sc_hd__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_4 abstract view
.subckt sky130_fd_sc_hd__nand3b_4 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_2 abstract view
.subckt sky130_fd_sc_hd__o32a_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_2 abstract view
.subckt sky130_fd_sc_hd__o41a_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_4 abstract view
.subckt sky130_fd_sc_hd__nand2b_4 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_2 abstract view
.subckt sky130_fd_sc_hd__o2111a_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_4 abstract view
.subckt sky130_fd_sc_hd__dfstp_4 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_4 abstract view
.subckt sky130_fd_sc_hd__a31o_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_2 abstract view
.subckt sky130_fd_sc_hd__and4bb_2 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_16 abstract view
.subckt sky130_fd_sc_hd__clkinv_16 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_4 abstract view
.subckt sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_2 abstract view
.subckt sky130_fd_sc_hd__a311o_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_4 abstract view
.subckt sky130_fd_sc_hd__o2111a_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_1 abstract view
.subckt sky130_fd_sc_hd__nand4b_1 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2oi_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2oi_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_2 abstract view
.subckt sky130_fd_sc_hd__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_1 abstract view
.subckt sky130_fd_sc_hd__nor4b_1 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_4 abstract view
.subckt sky130_fd_sc_hd__and4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_2 abstract view
.subckt sky130_fd_sc_hd__a2111oi_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_2 abstract view
.subckt sky130_fd_sc_hd__a221oi_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_2 abstract view
.subckt sky130_fd_sc_hd__a311oi_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_4 abstract view
.subckt sky130_fd_sc_hd__a211o_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_4 abstract view
.subckt sky130_fd_sc_hd__o41a_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_4 abstract view
.subckt sky130_fd_sc_hd__o2111ai_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_2 abstract view
.subckt sky130_fd_sc_hd__dfstp_2 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_2 abstract view
.subckt sky130_fd_sc_hd__o221a_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_2 abstract view
.subckt sky130_fd_sc_hd__nand3b_2 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

.subckt team_09 clk en gpio_in[0] gpio_in[10] gpio_in[11] gpio_in[12] gpio_in[13]
+ gpio_in[14] gpio_in[15] gpio_in[16] gpio_in[17] gpio_in[18] gpio_in[19] gpio_in[1]
+ gpio_in[20] gpio_in[21] gpio_in[22] gpio_in[23] gpio_in[24] gpio_in[25] gpio_in[26]
+ gpio_in[27] gpio_in[28] gpio_in[29] gpio_in[2] gpio_in[30] gpio_in[31] gpio_in[32]
+ gpio_in[33] gpio_in[3] gpio_in[4] gpio_in[5] gpio_in[6] gpio_in[7] gpio_in[8] gpio_in[9]
+ gpio_oeb[0] gpio_oeb[10] gpio_oeb[11] gpio_oeb[12] gpio_oeb[13] gpio_oeb[14] gpio_oeb[15]
+ gpio_oeb[16] gpio_oeb[17] gpio_oeb[18] gpio_oeb[19] gpio_oeb[1] gpio_oeb[20] gpio_oeb[21]
+ gpio_oeb[22] gpio_oeb[23] gpio_oeb[24] gpio_oeb[25] gpio_oeb[26] gpio_oeb[27] gpio_oeb[28]
+ gpio_oeb[29] gpio_oeb[2] gpio_oeb[30] gpio_oeb[31] gpio_oeb[32] gpio_oeb[33] gpio_oeb[3]
+ gpio_oeb[4] gpio_oeb[5] gpio_oeb[6] gpio_oeb[7] gpio_oeb[8] gpio_oeb[9] gpio_out[0]
+ gpio_out[10] gpio_out[11] gpio_out[12] gpio_out[13] gpio_out[14] gpio_out[15] gpio_out[16]
+ gpio_out[17] gpio_out[18] gpio_out[19] gpio_out[1] gpio_out[20] gpio_out[21] gpio_out[22]
+ gpio_out[23] gpio_out[24] gpio_out[25] gpio_out[26] gpio_out[27] gpio_out[28] gpio_out[29]
+ gpio_out[2] gpio_out[30] gpio_out[31] gpio_out[32] gpio_out[33] gpio_out[3] gpio_out[4]
+ gpio_out[5] gpio_out[6] gpio_out[7] gpio_out[8] gpio_out[9] nrst vccd1 vssd1
XFILLER_0_20_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18243__B1 net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10669__A1 net1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10669__B2 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09671_ _04635_ _04639_ _04642_ vssd1 vssd1 vccd1 vccd1 _04644_ sky130_fd_sc_hd__a21oi_2
X_18869_ clknet_leaf_26_clk img_gen.tracker.next_frame\[307\] net1342 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[307\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_74_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10958__B net1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14804__B1 ag2.body\[291\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10310__Y _05283_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14280__A1 net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout162_A net183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14280__B2 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_3999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10974__A net1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1071_A net1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14446__A net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout427_A net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1169_A net1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12043__B1 net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_227 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10693__B net1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__20228__CLK clknet_leaf_66_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_884 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09105_ ag2.body\[365\] vssd1 vssd1 vccd1 vccd1 _04130_ sky130_fd_sc_hd__inv_2
XFILLER_0_115_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09036_ ag2.body\[195\] vssd1 vssd1 vccd1 vccd1 _04061_ sky130_fd_sc_hd__inv_2
XFILLER_0_32_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17476__B net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_107_Left_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout796_A net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1556 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold340 img_gen.tracker.frame\[269\] vssd1 vssd1 vccd1 vccd1 net1902 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1503_A net1504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold351 img_gen.tracker.frame\[252\] vssd1 vssd1 vccd1 vccd1 net1913 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold362 img_gen.tracker.frame\[551\] vssd1 vssd1 vccd1 vccd1 net1924 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold373 img_gen.tracker.frame\[431\] vssd1 vssd1 vccd1 vccd1 net1935 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_51_clk_X clknet_leaf_51_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold384 img_gen.tracker.frame\[317\] vssd1 vssd1 vccd1 vccd1 net1946 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout963_A net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold395 img_gen.tracker.frame\[436\] vssd1 vssd1 vccd1 vccd1 net1957 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout820 net823 vssd1 vssd1 vccd1 vccd1 net820 sky130_fd_sc_hd__buf_4
XANTENNA_fanout584_X net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout831 _03966_ vssd1 vssd1 vccd1 vccd1 net831 sky130_fd_sc_hd__buf_4
XFILLER_0_99_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20127_ clknet_leaf_81_clk _01071_ net1485 vssd1 vssd1 vccd1 vccd1 ag2.body\[269\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__15835__A2 net204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout842 net847 vssd1 vssd1 vccd1 vccd1 net842 sky130_fd_sc_hd__buf_4
X_09938_ ag2.body\[26\] net774 _04904_ _04905_ _04907_ vssd1 vssd1 vccd1 vccd1 _04911_
+ sky130_fd_sc_hd__a2111o_1
XFILLER_0_99_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout853 net857 vssd1 vssd1 vccd1 vccd1 net853 sky130_fd_sc_hd__buf_4
XANTENNA__10214__A net1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13846__B2 ag2.body\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout864 net867 vssd1 vssd1 vccd1 vccd1 net864 sky130_fd_sc_hd__buf_4
Xfanout875 net878 vssd1 vssd1 vccd1 vccd1 net875 sky130_fd_sc_hd__buf_2
X_20058_ clknet_leaf_72_clk _01002_ net1501 vssd1 vssd1 vccd1 vccd1 ag2.body\[328\]
+ sky130_fd_sc_hd__dfrtp_4
Xfanout886 net889 vssd1 vssd1 vccd1 vccd1 net886 sky130_fd_sc_hd__clkbuf_8
XANTENNA__11857__B1 net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09869_ ag2.body\[153\] net1209 vssd1 vssd1 vccd1 vccd1 _04842_ sky130_fd_sc_hd__xor2_1
XANTENNA_fanout751_X net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout897 net898 vssd1 vssd1 vccd1 vccd1 net897 sky130_fd_sc_hd__clkbuf_2
XANTENNA__14415__A1_N net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1040 control.body\[908\] vssd1 vssd1 vccd1 vccd1 net2602 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1493_X net1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_66_clk_X clknet_leaf_66_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout849_X net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1051 control.body\[939\] vssd1 vssd1 vccd1 vccd1 net2613 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11321__A2 net1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1364 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11900_ img_gen.tracker.frame\[52\] net596 net541 img_gen.tracker.frame\[55\] _06871_
+ vssd1 vssd1 vccd1 vccd1 _06872_ sky130_fd_sc_hd__o221a_1
Xhold1062 control.body\[655\] vssd1 vssd1 vccd1 vccd1 net2624 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1073 control.body\[817\] vssd1 vssd1 vccd1 vccd1 net2635 sky130_fd_sc_hd__dlygate4sd3_1
X_12880_ net292 _07425_ _07638_ _07640_ net1875 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[197\]
+ sky130_fd_sc_hd__a32o_1
XPHY_EDGE_ROW_116_Left_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1084 control.body\[814\] vssd1 vssd1 vccd1 vccd1 net2646 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_96_910 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1095 control.body\[892\] vssd1 vssd1 vccd1 vccd1 net2657 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10868__B net1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11609__B1 net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11831_ img_gen.tracker.frame\[551\] net579 net541 img_gen.tracker.frame\[548\] _06802_
+ vssd1 vssd1 vccd1 vccd1 _06803_ sky130_fd_sc_hd__o221a_1
XFILLER_0_16_1602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15740__A _05253_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14550_ _08707_ _08708_ _08710_ _08706_ vssd1 vssd1 vccd1 vccd1 _08711_ sky130_fd_sc_hd__a211o_1
XFILLER_0_67_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11762_ img_gen.tracker.frame\[266\] net622 net550 img_gen.tracker.frame\[272\] _06733_
+ vssd1 vssd1 vccd1 vccd1 _06734_ sky130_fd_sc_hd__o221a_1
XFILLER_0_138_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13501_ net666 _07912_ vssd1 vssd1 vccd1 vccd1 _07913_ sky130_fd_sc_hd__nor2_1
X_10713_ _04600_ _05346_ _05685_ vssd1 vssd1 vccd1 vccd1 _05686_ sky130_fd_sc_hd__a21oi_4
X_14481_ net842 ag2.body\[440\] ag2.body\[447\] net792 _08639_ vssd1 vssd1 vccd1 vccd1
+ _08642_ sky130_fd_sc_hd__a221o_1
X_11693_ img_gen.tracker.frame\[110\] net619 net602 img_gen.tracker.frame\[113\] vssd1
+ vssd1 vccd1 vccd1 _06665_ sky130_fd_sc_hd__o22a_1
XFILLER_0_67_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_124_clk_X clknet_leaf_124_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16220_ net537 _01889_ _01897_ _01737_ vssd1 vssd1 vccd1 vccd1 _01899_ sky130_fd_sc_hd__a22o_1
XFILLER_0_10_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12034__B1 net557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13432_ net236 _07884_ _07885_ net1588 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[504\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__20508__D net2301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10644_ _04573_ _05615_ _05616_ vssd1 vssd1 vccd1 vccd1 _05617_ sky130_fd_sc_hd__or3_1
XANTENNA__16036__D_N net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12585__A1 net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16151_ obsg2.obstacleArray\[22\] obsg2.obstacleArray\[23\] net429 vssd1 vssd1 vccd1
+ vccd1 _01830_ sky130_fd_sc_hd__mux2_1
X_10575_ ag2.body\[190\] net1080 vssd1 vssd1 vccd1 vccd1 _05548_ sky130_fd_sc_hd__or2_1
X_13363_ net670 _07858_ vssd1 vssd1 vccd1 vccd1 _07859_ sky130_fd_sc_hd__nor2_1
XFILLER_0_88_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_125_Left_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15102_ _04557_ net58 vssd1 vssd1 vccd1 vccd1 _01564_ sky130_fd_sc_hd__nor2_2
XANTENNA__10060__A2 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12314_ _07221_ _07274_ _07278_ _07280_ _07268_ vssd1 vssd1 vccd1 vccd1 _07281_ sky130_fd_sc_hd__a2111o_1
XANTENNA__17386__B net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16082_ obsg2.obstacleArray\[98\] net421 vssd1 vssd1 vccd1 vccd1 _01761_ sky130_fd_sc_hd__or2_1
XANTENNA__16720__B1 net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13294_ net671 _07831_ vssd1 vssd1 vccd1 vccd1 _07832_ sky130_fd_sc_hd__nor2_1
XFILLER_0_126_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18768__CLK clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19910_ clknet_leaf_56_clk _00854_ net1457 vssd1 vssd1 vccd1 vccd1 ag2.body\[484\]
+ sky130_fd_sc_hd__dfrtp_4
X_15033_ control.body\[969\] net165 _01557_ control.body\[961\] vssd1 vssd1 vccd1
+ vccd1 _00363_ sky130_fd_sc_hd__a22o_1
XFILLER_0_20_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12245_ img_gen.updater.commands.cmd_num\[0\] _07207_ vssd1 vssd1 vccd1 vccd1 _07215_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_62_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09456__Y _04429_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14091__A net1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12176_ _07039_ _07093_ _07145_ _07146_ vssd1 vssd1 vccd1 vccd1 _07148_ sky130_fd_sc_hd__a22o_1
X_19841_ clknet_leaf_122_clk _00785_ net1414 vssd1 vssd1 vccd1 vccd1 ag2.body\[559\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_62_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11127_ net1131 control.body\[868\] vssd1 vssd1 vccd1 vccd1 _06100_ sky130_fd_sc_hd__and2b_1
XANTENNA__16510__S net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16984_ _04016_ net885 net735 ag2.body\[89\] vssd1 vssd1 vccd1 vccd1 _02663_ sky130_fd_sc_hd__a22o_1
XFILLER_0_78_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10124__A net1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19772_ clknet_leaf_127_clk _00716_ net1331 vssd1 vssd1 vccd1 vccd1 ag2.body\[618\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_120_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13837__B2 net1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11058_ ag2.body\[436\] net1127 vssd1 vssd1 vccd1 vccd1 _06031_ sky130_fd_sc_hd__xnor2_1
X_15935_ ag2.body\[173\] net138 _01655_ ag2.body\[165\] vssd1 vssd1 vccd1 vccd1 _01167_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_120_1288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18723_ clknet_leaf_142_clk img_gen.tracker.next_frame\[161\] net1254 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[161\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_120_1299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_1431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_134_Left_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09992__A1_N net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13435__A _07572_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10009_ net891 _04239_ _04980_ vssd1 vssd1 vccd1 vccd1 _04982_ sky130_fd_sc_hd__or3b_2
X_18654_ clknet_leaf_131_clk img_gen.tracker.next_frame\[92\] net1312 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[92\] sky130_fd_sc_hd__dfrtp_1
X_15866_ ag2.body\[224\] net161 _01647_ ag2.body\[216\] vssd1 vssd1 vccd1 vccd1 _01106_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_133_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17605_ _04148_ net872 net714 ag2.body\[420\] _03278_ vssd1 vssd1 vccd1 vccd1 _03284_
+ sky130_fd_sc_hd__a221o_1
X_14817_ net793 ag2.body\[383\] _01483_ _01487_ vssd1 vssd1 vccd1 vccd1 _01488_ sky130_fd_sc_hd__a211o_1
XANTENNA__13154__B net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18585_ clknet_leaf_15_clk img_gen.tracker.next_frame\[23\] net1277 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[23\] sky130_fd_sc_hd__dfrtp_1
X_15797_ ag2.body\[290\] net207 _01640_ ag2.body\[282\] vssd1 vssd1 vccd1 vccd1 _01044_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__14818__X _01489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_280 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15650__A _05152_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17536_ ag2.body\[272\] net740 net699 ag2.body\[278\] _03214_ vssd1 vssd1 vccd1 vccd1
+ _03215_ sky130_fd_sc_hd__a221o_1
X_14748_ net1003 ag2.body\[104\] vssd1 vssd1 vccd1 vccd1 _08909_ sky130_fd_sc_hd__xor2_1
XANTENNA__17736__C1 _03206_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10823__A1 net1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17467_ ag2.body\[528\] net886 vssd1 vssd1 vccd1 vccd1 _03146_ sky130_fd_sc_hd__xor2_1
X_14679_ net1037 ag2.body\[388\] vssd1 vssd1 vccd1 vccd1 _08840_ sky130_fd_sc_hd__xor2_1
XFILLER_0_104_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14266__A net999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16418_ obsg2.obstacleArray\[114\] obsg2.obstacleArray\[115\] net455 vssd1 vssd1
+ vccd1 vccd1 _02097_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_1257 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19206_ clknet_leaf_86_clk _00150_ net1461 vssd1 vssd1 vccd1 vccd1 ag2.body\[69\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__19543__CLK clknet_leaf_118_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12025__B1 net557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17398_ ag2.body\[506\] net727 net932 _04187_ _03072_ vssd1 vssd1 vccd1 vccd1 _03077_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_73_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11379__A2 net1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19137_ clknet_leaf_140_clk img_gen.tracker.next_frame\[575\] net1297 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[575\] sky130_fd_sc_hd__dfrtp_1
X_16349_ _02016_ _02020_ _02027_ _01912_ _01918_ vssd1 vssd1 vccd1 vccd1 _02028_ sky130_fd_sc_hd__a221o_1
XANTENNA__11402__B net1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17503__A2 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__20173__RESET_B net1480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20520__CLK clknet_leaf_93_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19068_ clknet_leaf_29_clk img_gen.tracker.next_frame\[506\] net1335 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[506\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__17296__B net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_114_3792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18019_ net45 _03628_ vssd1 vssd1 vccd1 vccd1 _03629_ sky130_fd_sc_hd__nor2_1
XFILLER_0_113_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12514__A net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12879__A2 _07425_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_3667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09095__A ag2.body\[340\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_3678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20504__Q ag2.goodColl vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_3689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout105 net107 vssd1 vssd1 vccd1 vccd1 net105 sky130_fd_sc_hd__buf_2
Xfanout116 net117 vssd1 vssd1 vccd1 vccd1 net116 sky130_fd_sc_hd__buf_2
Xfanout127 net128 vssd1 vssd1 vccd1 vccd1 net127 sky130_fd_sc_hd__clkbuf_4
Xfanout138 net139 vssd1 vssd1 vccd1 vccd1 net138 sky130_fd_sc_hd__clkbuf_4
Xfanout149 net154 vssd1 vssd1 vccd1 vccd1 net149 sky130_fd_sc_hd__buf_2
XANTENNA__13048__C _07638_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09823__A net1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09723_ net909 _04637_ vssd1 vssd1 vccd1 vccd1 _04696_ sky130_fd_sc_hd__nand2_1
XFILLER_0_38_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11839__B1 net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10969__A net1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout377_A net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09654_ net1150 control.body\[747\] vssd1 vssd1 vccd1 vccd1 _04627_ sky130_fd_sc_hd__xor2_1
XANTENNA__16778__B1 net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10688__B net1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14253__A1 net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09585_ net1131 control.body\[908\] vssd1 vssd1 vccd1 vccd1 _04558_ sky130_fd_sc_hd__xor2_1
XANTENNA_fanout544_A net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14253__B2 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15450__B1 _01601_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1286_A net1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16375__B net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout332_X net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout711_A net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14176__A net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1453_A net1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15202__B1 _01574_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16943__X _02622_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout809_A net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1074_X net1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_1508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12016__B1 net557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16950__B1 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_93_clk_A clknet_4_11__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_810 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11312__B net1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10209__A net1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10360_ ag2.body\[294\] net752 _05330_ _05331_ _05332_ vssd1 vssd1 vccd1 vccd1 _05333_
+ sky130_fd_sc_hd__a2111o_1
XFILLER_0_5_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16702__B1 net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_230 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout799_X net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09019_ ag2.body\[153\] vssd1 vssd1 vccd1 vccd1 _04044_ sky130_fd_sc_hd__inv_2
XANTENNA__17774__X _03453_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10291_ ag2.body\[334\] net1090 vssd1 vssd1 vccd1 vccd1 _05264_ sky130_fd_sc_hd__nand2_1
XANTENNA__11527__C1 net1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12030_ img_gen.tracker.frame\[24\] net629 net594 img_gen.tracker.frame\[33\] vssd1
+ vssd1 vccd1 vccd1 _07002_ sky130_fd_sc_hd__a22o_1
XANTENNA__09735__A2 net1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold170 img_gen.tracker.frame\[95\] vssd1 vssd1 vccd1 vccd1 net1732 sky130_fd_sc_hd__dlygate4sd3_1
Xhold181 img_gen.tracker.frame\[132\] vssd1 vssd1 vccd1 vccd1 net1743 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout966_X net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12143__B net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold192 img_gen.tracker.frame\[135\] vssd1 vssd1 vccd1 vccd1 net1754 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__16330__S net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18111__A net44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_31_clk_A clknet_4_4__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout650 net651 vssd1 vssd1 vccd1 vccd1 net650 sky130_fd_sc_hd__buf_1
Xfanout661 _04394_ vssd1 vssd1 vccd1 vccd1 net661 sky130_fd_sc_hd__clkbuf_2
Xfanout672 net674 vssd1 vssd1 vccd1 vccd1 net672 sky130_fd_sc_hd__buf_2
X_13981_ ag2.body\[119\] net203 _08158_ ag2.body\[111\] vssd1 vssd1 vccd1 vccd1 _00200_
+ sky130_fd_sc_hd__a22o_1
Xfanout683 net684 vssd1 vssd1 vccd1 vccd1 net683 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09499__A1 _04427_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14492__A1 net1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout694 net695 vssd1 vssd1 vccd1 vccd1 net694 sky130_fd_sc_hd__buf_4
XANTENNA__19416__CLK clknet_leaf_103_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14492__B2 net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15720_ ag2.body\[367\] net193 _01630_ ag2.body\[359\] vssd1 vssd1 vccd1 vccd1 _00977_
+ sky130_fd_sc_hd__a22o_1
X_12932_ img_gen.tracker.frame\[226\] net660 vssd1 vssd1 vccd1 vccd1 _07664_ sky130_fd_sc_hd__and2_1
XANTENNA__16769__B1 net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15651_ ag2.body\[416\] net139 _01624_ ag2.body\[408\] vssd1 vssd1 vccd1 vccd1 _00914_
+ sky130_fd_sc_hd__a22o_1
X_12863_ net286 _07631_ _07632_ net1702 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[188\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_46_clk_A clknet_4_7__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14602_ net829 ag2.body\[130\] ag2.body\[134\] net803 vssd1 vssd1 vccd1 vccd1 _08763_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_9_1566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15470__A _05133_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18370_ _08138_ _03860_ vssd1 vssd1 vccd1 vccd1 _03863_ sky130_fd_sc_hd__nor2_1
X_11814_ img_gen.tracker.frame\[470\] net616 net600 img_gen.tracker.frame\[473\] _06785_
+ vssd1 vssd1 vccd1 vccd1 _06786_ sky130_fd_sc_hd__o221a_1
XFILLER_0_115_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15582_ ag2.body\[482\] net130 _01617_ ag2.body\[474\] vssd1 vssd1 vccd1 vccd1 _00852_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__19566__CLK clknet_leaf_115_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12794_ net252 _07599_ _07600_ net1995 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[151\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_51_1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17321_ ag2.body\[218\] net727 net719 ag2.body\[219\] vssd1 vssd1 vccd1 vccd1 _03000_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_84_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14533_ net1001 _04079_ ag2.body\[251\] net820 vssd1 vssd1 vccd1 vccd1 _08694_ sky130_fd_sc_hd__a22o_1
XFILLER_0_138_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17949__X _03577_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11745_ net565 _06707_ _06710_ net470 vssd1 vssd1 vccd1 vccd1 _06717_ sky130_fd_sc_hd__a211o_1
XANTENNA__14086__A net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_137_4493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20543__CLK clknet_leaf_105_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12007__B1 net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17252_ ag2.body\[544\] net881 vssd1 vssd1 vccd1 vccd1 _02931_ sky130_fd_sc_hd__xor2_1
XANTENNA__15744__A1 ag2.body\[339\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_467 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14464_ net1001 ag2.body\[264\] vssd1 vssd1 vccd1 vccd1 _08625_ sky130_fd_sc_hd__nand2_1
X_11676_ _06639_ _06640_ vssd1 vssd1 vccd1 vccd1 _06648_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_43_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16941__B1 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_133_4368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16203_ obsg2.obstacleArray\[56\] obsg2.obstacleArray\[57\] obsg2.obstacleArray\[58\]
+ obsg2.obstacleArray\[59\] net424 net377 vssd1 vssd1 vccd1 vccd1 _01882_ sky130_fd_sc_hd__mux4_1
XFILLER_0_128_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18590__CLK clknet_leaf_13_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13415_ _07561_ net302 vssd1 vssd1 vccd1 vccd1 _07878_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_133_4379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10627_ _05590_ _05591_ _05595_ _05599_ vssd1 vssd1 vccd1 vccd1 _05600_ sky130_fd_sc_hd__or4_1
X_17183_ ag2.body\[570\] net859 vssd1 vssd1 vccd1 vccd1 _02862_ sky130_fd_sc_hd__nand2_1
X_14395_ net993 _04029_ ag2.body\[124\] net815 vssd1 vssd1 vccd1 vccd1 _08556_ sky130_fd_sc_hd__a22o_1
XANTENNA__16505__S net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10119__A net1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_104_clk_A clknet_4_10__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14814__A net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_1290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_12_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11766__C1 net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16134_ _01777_ _01812_ _01724_ vssd1 vssd1 vccd1 vccd1 _01813_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_12_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13346_ net274 _07850_ _07851_ net1825 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[452\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_45_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_1420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10558_ ag2.body\[513\] net1203 vssd1 vssd1 vccd1 vccd1 _05531_ sky130_fd_sc_hd__xor2_1
XFILLER_0_24_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11781__A2 net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16065_ obsg2.obstacleArray\[105\] net430 vssd1 vssd1 vccd1 vccd1 _01744_ sky130_fd_sc_hd__or2_1
X_13277_ net280 _07823_ _07824_ net1787 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[410\]
+ sky130_fd_sc_hd__a22o_1
X_10489_ _05458_ _05459_ _05461_ vssd1 vssd1 vccd1 vccd1 _05462_ sky130_fd_sc_hd__and3_1
XFILLER_0_126_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15016_ control.body\[988\] net152 _01553_ net2384 vssd1 vssd1 vccd1 vccd1 _00350_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__09726__A2 net1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12228_ img_gen.updater.commands.cmd_num\[3\] _07197_ vssd1 vssd1 vccd1 vccd1 _07198_
+ sky130_fd_sc_hd__nand2_1
XANTENNA_clkbuf_leaf_119_clk_A clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16457__C1 _02075_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12730__A1 net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19824_ clknet_4_9__leaf_clk _00768_ net1411 vssd1 vssd1 vccd1 vccd1 ag2.body\[574\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_120_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12159_ _07127_ _07128_ _07130_ net558 vssd1 vssd1 vccd1 vccd1 _07131_ sky130_fd_sc_hd__a22o_1
XFILLER_0_75_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19755_ clknet_leaf_130_clk _00699_ net1315 vssd1 vssd1 vccd1 vccd1 control.body\[633\]
+ sky130_fd_sc_hd__dfrtp_1
X_16967_ ag2.body\[409\] net872 vssd1 vssd1 vccd1 vccd1 _02646_ sky130_fd_sc_hd__xor2_1
XANTENNA__13286__A2 _07827_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10789__A net1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15680__B1 _01627_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18706_ clknet_leaf_144_clk img_gen.tracker.next_frame\[144\] net1255 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[144\] sky130_fd_sc_hd__dfrtp_1
X_15918_ ag2.body\[191\] net131 _01652_ ag2.body\[183\] vssd1 vssd1 vccd1 vccd1 _01153_
+ sky130_fd_sc_hd__a22o_1
X_16898_ _02573_ _02574_ _02576_ vssd1 vssd1 vccd1 vccd1 _02577_ sky130_fd_sc_hd__and3_1
X_19686_ clknet_leaf_135_clk _00630_ net1302 vssd1 vssd1 vccd1 vccd1 control.body\[708\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_56_1223 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__20073__CLK clknet_leaf_73_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18637_ clknet_leaf_131_clk img_gen.tracker.next_frame\[75\] net1297 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[75\] sky130_fd_sc_hd__dfrtp_1
X_15849_ ag2.body\[241\] net173 _01645_ ag2.body\[233\] vssd1 vssd1 vccd1 vccd1 _01091_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__14235__A1 net1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_103_3460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14235__B2 net1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_3471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09370_ net271 _04369_ _04370_ vssd1 vssd1 vccd1 vccd1 _01419_ sky130_fd_sc_hd__and3_1
XFILLER_0_73_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18568_ clknet_leaf_15_clk img_gen.tracker.next_frame\[6\] net1313 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[6\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_75_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17519_ ag2.body\[481\] net869 vssd1 vssd1 vccd1 vccd1 _03198_ sky130_fd_sc_hd__xor2_1
XFILLER_0_46_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18499_ net1514 net1508 vssd1 vssd1 vccd1 vccd1 _00030_ sky130_fd_sc_hd__or2_1
XFILLER_0_30_1418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11413__A net1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20530_ clknet_leaf_112_clk _01395_ net1424 vssd1 vssd1 vccd1 vccd1 toggle1.bcd_ones\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_28_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15735__B2 ag2.body\[339\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16923__B net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkload64_A clknet_leaf_53_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20461_ clknet_leaf_31_clk _01348_ net1338 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[97\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_116_3854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout125_A net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_116_3865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14724__A net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_116_3876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_3729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10024__A2 _04968_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20392_ clknet_leaf_38_clk _01279_ net1354 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[28\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_28_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11772__A2 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1034_A net1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09717__A2 net1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17754__B _03429_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout494_A _01736_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16448__C1 net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_2482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1201_A net1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_71_2493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09553__A net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout282_X net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout661_A _04394_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout759_A net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09706_ _04665_ _04666_ _04675_ _04678_ vssd1 vssd1 vccd1 vccd1 _04679_ sky130_fd_sc_hd__a211o_1
XFILLER_0_138_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19589__CLK clknet_leaf_118_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09637_ net787 control.body\[1016\] control.body\[1019\] net771 _04609_ vssd1 vssd1
+ vccd1 vccd1 _04610_ sky130_fd_sc_hd__o221ai_1
XANTENNA__11307__B net1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14226__A1 net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16386__A net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1191_X net1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout547_X net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14226__B2 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_2876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__20566__CLK clknet_leaf_43_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_2887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15974__A1 net223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_2898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09568_ ag2.body\[206\] net1089 vssd1 vssd1 vccd1 vccd1 _04541_ sky130_fd_sc_hd__xor2_1
XFILLER_0_116_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1632 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout38_A net39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_710 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_2297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12788__A1 net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12419__A net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout714_X net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09499_ _04427_ _04471_ net642 vssd1 vssd1 vccd1 vccd1 _04472_ sky130_fd_sc_hd__a21o_1
XANTENNA__20095__RESET_B net1492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10865__C _05812_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11530_ _06489_ _06502_ _06497_ vssd1 vssd1 vccd1 vccd1 _06503_ sky130_fd_sc_hd__or3b_1
XFILLER_0_33_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17929__B net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16833__B net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_137_Right_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11461_ ag2.body\[262\] net1091 vssd1 vssd1 vccd1 vccd1 _06434_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_22_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13200_ _07790_ net263 _07788_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[367\]
+ sky130_fd_sc_hd__mux2_1
X_10412_ _05379_ _05380_ _05383_ _05384_ vssd1 vssd1 vccd1 vccd1 _05385_ sky130_fd_sc_hd__or4_1
XFILLER_0_85_1463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14180_ _08337_ _08338_ _08340_ _08334_ vssd1 vssd1 vccd1 vccd1 _08341_ sky130_fd_sc_hd__a211o_1
X_11392_ net1195 control.body\[641\] vssd1 vssd1 vccd1 vccd1 _06365_ sky130_fd_sc_hd__xor2_1
XANTENNA__09810__D1 _04711_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18140__A2 _03558_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16687__C1 net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13131_ _07757_ net265 _07755_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[331\]
+ sky130_fd_sc_hd__mux2_1
XANTENNA__12960__A1 net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10343_ ag2.body\[521\] net780 net775 ag2.body\[522\] vssd1 vssd1 vccd1 vccd1 _05316_
+ sky130_fd_sc_hd__o22ai_1
XFILLER_0_131_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14921__X _01543_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09708__A2 net1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10274_ ag2.body\[136\] net1235 vssd1 vssd1 vccd1 vccd1 _05247_ sky130_fd_sc_hd__nand2_1
X_13062_ img_gen.tracker.frame\[295\] net660 vssd1 vssd1 vccd1 vccd1 _07725_ sky130_fd_sc_hd__and2_1
XFILLER_0_29_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12712__A1 net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12013_ net385 _06958_ _06984_ _06724_ net382 vssd1 vssd1 vccd1 vccd1 _06985_ sky130_fd_sc_hd__o2111a_1
XANTENNA__17678__A2_N net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17870_ net2263 _03504_ vssd1 vssd1 vccd1 vccd1 _01242_ sky130_fd_sc_hd__xor2_1
Xfanout1401 net1402 vssd1 vssd1 vccd1 vccd1 net1401 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_40_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1412 net1413 vssd1 vssd1 vccd1 vccd1 net1412 sky130_fd_sc_hd__clkbuf_4
Xfanout1423 net1435 vssd1 vssd1 vccd1 vccd1 net1423 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_TAPCELL_ROW_126_4161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1434 net1435 vssd1 vssd1 vccd1 vccd1 net1434 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_40_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1445 net1448 vssd1 vssd1 vccd1 vccd1 net1445 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_126_4172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16821_ _02492_ _02495_ _02499_ vssd1 vssd1 vccd1 vccd1 _02500_ sky130_fd_sc_hd__and3_1
XANTENNA__18549__Q ag2.y\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1456 net1458 vssd1 vssd1 vccd1 vccd1 net1456 sky130_fd_sc_hd__clkbuf_4
Xfanout1467 net1468 vssd1 vssd1 vccd1 vccd1 net1467 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_50_1843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_122_4036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1478 net1505 vssd1 vssd1 vccd1 vccd1 net1478 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_50_1854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_4047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout491 net492 vssd1 vssd1 vccd1 vccd1 net491 sky130_fd_sc_hd__clkbuf_4
Xfanout1489 net1493 vssd1 vssd1 vccd1 vccd1 net1489 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_6_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16752_ obsg2.obstacleArray\[43\] net500 net486 obsg2.obstacleArray\[42\] vssd1 vssd1
+ vccd1 vccd1 _02431_ sky130_fd_sc_hd__a22o_1
X_19540_ clknet_leaf_113_clk _00484_ net1396 vssd1 vssd1 vccd1 vccd1 control.body\[850\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_122_4058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13964_ _05347_ net67 vssd1 vssd1 vccd1 vccd1 _08157_ sky130_fd_sc_hd__and2_2
XFILLER_0_92_1412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_31_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09750__X _04723_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15703_ _04434_ net63 vssd1 vssd1 vccd1 vccd1 _01629_ sky130_fd_sc_hd__and2_2
X_12915_ net265 _07654_ _07655_ net1728 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[217\]
+ sky130_fd_sc_hd__a22o_1
X_16683_ _02244_ _02356_ _02357_ _02361_ _02262_ vssd1 vssd1 vccd1 vccd1 _02362_ sky130_fd_sc_hd__a311oi_1
X_19471_ clknet_leaf_110_clk net2197 net1419 vssd1 vssd1 vccd1 vccd1 control.body\[925\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10896__X _05869_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13895_ ag2.body\[42\] net118 _08149_ ag2.body\[34\] vssd1 vssd1 vccd1 vccd1 _00123_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__18956__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15634_ ag2.body\[433\] net126 _01622_ ag2.body\[425\] vssd1 vssd1 vccd1 vccd1 _00899_
+ sky130_fd_sc_hd__a22o_1
X_18422_ track.nextHighScore\[1\] _03782_ _03807_ vssd1 vssd1 vccd1 vccd1 _03911_
+ sky130_fd_sc_hd__a21boi_1
XFILLER_0_69_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09910__B net1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12846_ net388 _07535_ vssd1 vssd1 vccd1 vccd1 _07624_ sky130_fd_sc_hd__nand2_2
XFILLER_0_61_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18353_ _03846_ _03848_ _03819_ vssd1 vssd1 vccd1 vccd1 _03849_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_31_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_48_1783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15565_ ag2.body\[500\] net185 _01614_ ag2.body\[492\] vssd1 vssd1 vccd1 vccd1 _00838_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_51_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09644__A1 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17167__B1 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12777_ net1907 net648 _07590_ _07591_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[143\]
+ sky130_fd_sc_hd__a31o_1
XANTENNA__09644__B2 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_968 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17304_ ag2.body\[350\] net701 _02981_ _02982_ vssd1 vssd1 vccd1 vccd1 _02983_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_29_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14516_ net1041 ag2.body\[316\] vssd1 vssd1 vccd1 vccd1 _08677_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_44_1658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18284_ net319 _03587_ obsg2.obstacleArray\[139\] vssd1 vssd1 vccd1 vccd1 _03781_
+ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_44_1669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11728_ img_gen.tracker.frame\[206\] net624 vssd1 vssd1 vccd1 vccd1 _06700_ sky130_fd_sc_hd__or2_1
X_15496_ ag2.body\[567\] net110 _01606_ ag2.body\[559\] vssd1 vssd1 vccd1 vccd1 _00777_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_71_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17235_ ag2.body\[442\] net724 net709 ag2.body\[444\] vssd1 vssd1 vccd1 vccd1 _02914_
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_9_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_104_Right_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14447_ net992 ag2.body\[225\] vssd1 vssd1 vccd1 vccd1 _08608_ sky130_fd_sc_hd__xor2_1
X_11659_ _06628_ _06629_ vssd1 vssd1 vccd1 vccd1 _06632_ sky130_fd_sc_hd__nor2_1
XFILLER_0_25_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14246__A1_N net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17166_ ag2.body\[597\] net946 vssd1 vssd1 vccd1 vccd1 _02845_ sky130_fd_sc_hd__xor2_1
X_14378_ net1017 ag2.body\[422\] vssd1 vssd1 vccd1 vccd1 _08539_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_94_3183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_3194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold906 control.body\[1060\] vssd1 vssd1 vccd1 vccd1 net2468 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16117_ obsg2.obstacleArray\[94\] obsg2.obstacleArray\[95\] net425 vssd1 vssd1 vccd1
+ vccd1 _01796_ sky130_fd_sc_hd__mux2_1
Xhold917 control.body\[928\] vssd1 vssd1 vccd1 vccd1 net2479 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11754__A2 net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12951__A1 net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold928 control.body\[677\] vssd1 vssd1 vccd1 vccd1 net2490 sky130_fd_sc_hd__dlygate4sd3_1
X_13329_ net228 _07844_ _07845_ net1751 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[441\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_110_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_3058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17097_ _04099_ net965 obsg2.randCord\[6\] _04100_ vssd1 vssd1 vccd1 vccd1 _02776_
+ sky130_fd_sc_hd__a22o_1
Xhold939 control.body\[1050\] vssd1 vssd1 vccd1 vccd1 net2501 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_126_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_90_3069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20054__Q ag2.body\[340\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_3_1_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_3_1_0_clk sky130_fd_sc_hd__clkbuf_8
X_16048_ net497 _01726_ vssd1 vssd1 vccd1 vccd1 _01727_ sky130_fd_sc_hd__nand2_4
XFILLER_0_126_1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19807_ clknet_leaf_124_clk _00751_ net1405 vssd1 vssd1 vccd1 vccd1 ag2.body\[589\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__17642__B2 ag2.body\[167\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14456__A1 net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17999_ net299 _03613_ vssd1 vssd1 vccd1 vccd1 _03614_ sky130_fd_sc_hd__nand2_1
XANTENNA__14456__B2 net1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_3511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_105_3522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_3533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19738_ clknet_leaf_128_clk _00682_ net1329 vssd1 vssd1 vccd1 vccd1 control.body\[648\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14861__D1 _08181_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_3408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19669_ clknet_leaf_118_clk _00613_ net1301 vssd1 vssd1 vccd1 vccd1 control.body\[723\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09883__A1 ag2.body\[160\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15405__B1 _01581_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09422_ obsg2.obsNeeded\[2\] _04399_ _04400_ net1712 vssd1 vssd1 vccd1 vccd1 _00001_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_87_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09353_ sound_gen.osc1.stayCount\[10\] sound_gen.osc1.stayCount\[9\] _04354_ vssd1
+ vssd1 vccd1 vccd1 _04355_ sky130_fd_sc_hd__and3_1
XANTENNA__13342__B net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09635__A1 net1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09635__B2 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout242_A net247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_118_3916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_118_3927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20229__Q ag2.body\[163\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19111__CLK clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_2150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09284_ _04303_ _04305_ vssd1 vssd1 vccd1 vccd1 _04307_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_60_2161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1636 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20513_ clknet_leaf_113_clk track.nextHighScore\[3\] net1403 vssd1 vssd1 vccd1 vccd1
+ track.highScore\[3\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__11993__A2 net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10982__A net1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1151_A net1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12526__X _07460_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout128_X net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout507_A net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13195__A1 net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1249_A net1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20444_ clknet_leaf_42_clk _01331_ net1371 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[80\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_132_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09938__A2 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19261__CLK clknet_leaf_73_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12942__A1 net246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_2680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20375_ clknet_leaf_23_clk _01262_ net1359 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[11\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA_fanout1037_X net1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_2544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_2090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18829__CLK clknet_leaf_141_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload90 clknet_leaf_108_clk vssd1 vssd1 vccd1 vccd1 clkload90/Y sky130_fd_sc_hd__inv_8
XFILLER_0_30_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14695__A1 net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout876_A net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14695__B2 net1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout497_X net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11110__A_N net1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1204_X net1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12702__A net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09571__B1 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12170__A2 net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13517__B net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08999_ ag2.body\[99\] vssd1 vssd1 vccd1 vccd1 _04024_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout664_X net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18979__CLK clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15644__B1 _01623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17704__S net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_2359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout831_X net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10961_ ag2.body\[168\] net1224 vssd1 vssd1 vccd1 vccd1 _05934_ sky130_fd_sc_hd__xor2_1
XFILLER_0_39_1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14629__A net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout929_X net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12700_ net258 net310 _07553_ _07554_ net1624 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[103\]
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_116_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09730__B net1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13680_ _04238_ net639 vssd1 vssd1 vccd1 vccd1 _08025_ sky130_fd_sc_hd__xnor2_4
XANTENNA__10484__A2 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10892_ net1195 control.body\[649\] vssd1 vssd1 vccd1 vccd1 _05865_ sky130_fd_sc_hd__xor2_1
X_12631_ net225 _07516_ _07517_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[71\]
+ sky130_fd_sc_hd__o21bai_1
XANTENNA__13252__B net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11969__C1 net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15350_ net2559 net75 _01591_ control.body\[684\] vssd1 vssd1 vccd1 vccd1 _00646_
+ sky130_fd_sc_hd__a22o_1
X_12562_ net306 _07480_ vssd1 vssd1 vccd1 vccd1 _07481_ sky130_fd_sc_hd__nor2_1
XANTENNA__17659__B net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_264 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14301_ net838 ag2.body\[217\] ag2.body\[216\] net844 vssd1 vssd1 vccd1 vccd1 _08462_
+ sky130_fd_sc_hd__a2bb2o_1
X_11513_ obsg2.obstacleArray\[113\] obsg2.obstacleArray\[117\] net512 vssd1 vssd1
+ vccd1 vccd1 _06486_ sky130_fd_sc_hd__mux2_1
XANTENNA__11984__A2 net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15281_ net2238 net88 _01583_ control.body\[751\] vssd1 vssd1 vccd1 vccd1 _00585_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__10892__A net1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12493_ net1731 _07441_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[9\] sky130_fd_sc_hd__and2_1
XANTENNA__14364__A net1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17020_ ag2.body\[330\] net728 net935 _04117_ _02698_ vssd1 vssd1 vccd1 vccd1 _02699_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_108_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14232_ net996 _04173_ _04175_ net971 _08392_ vssd1 vssd1 vccd1 vccd1 _08393_ sky130_fd_sc_hd__a221o_1
X_11444_ net1229 control.body\[952\] vssd1 vssd1 vccd1 vccd1 _06417_ sky130_fd_sc_hd__or2_1
XFILLER_0_106_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11500__B net1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14163_ _08320_ _08321_ _08323_ vssd1 vssd1 vccd1 vccd1 _08324_ sky130_fd_sc_hd__nand3b_1
X_11375_ ag2.body\[472\] net1223 vssd1 vssd1 vccd1 vccd1 _06348_ sky130_fd_sc_hd__xor2_1
XANTENNA__17321__B1 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10944__B1 net1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_128_4212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13114_ img_gen.tracker.frame\[323\] net652 _07748_ vssd1 vssd1 vccd1 vccd1 _07749_
+ sky130_fd_sc_hd__and3_1
XANTENNA__19754__CLK clknet_leaf_127_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10326_ _05295_ _05296_ _05297_ _05298_ vssd1 vssd1 vccd1 vccd1 _05299_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_128_4223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14094_ _08247_ _08248_ _08251_ _08252_ _08254_ vssd1 vssd1 vccd1 vccd1 _08255_ sky130_fd_sc_hd__a221o_1
X_18971_ clknet_leaf_6_clk img_gen.tracker.next_frame\[409\] net1265 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[409\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_128_4234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14686__A1 net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13489__A2 net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14370__Y _08531_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14686__B2 net1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17922_ net318 _03555_ obsg2.obstacleArray\[2\] vssd1 vssd1 vccd1 vccd1 _03556_ sky130_fd_sc_hd__a21oi_1
Xclkbuf_4_2__f_clk clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_2__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_24_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13045_ net2124 net646 _07716_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[286\]
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_37_1462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09905__B net1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_4109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10257_ control.body\[789\] net1099 vssd1 vssd1 vccd1 vccd1 _05230_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_33_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10358__A_N net1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1220 net1221 vssd1 vssd1 vccd1 vccd1 net1220 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09562__B1 _04522_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12161__A2 net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1231 net1232 vssd1 vssd1 vccd1 vccd1 net1231 sky130_fd_sc_hd__buf_4
XFILLER_0_98_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17853_ img_gen.updater.commands.rR1.rainbowRNG\[15\] img_gen.updater.commands.rR1.rainbowRNG\[14\]
+ _03506_ _03508_ _07321_ vssd1 vssd1 vccd1 vccd1 _01231_ sky130_fd_sc_hd__a311o_1
Xfanout1242 net1243 vssd1 vssd1 vccd1 vccd1 net1242 sky130_fd_sc_hd__clkbuf_4
X_10188_ net912 net920 net916 net908 net900 vssd1 vssd1 vccd1 vccd1 _05161_ sky130_fd_sc_hd__a311o_1
Xfanout1253 net1254 vssd1 vssd1 vccd1 vccd1 net1253 sky130_fd_sc_hd__clkbuf_4
Xfanout1264 net1267 vssd1 vssd1 vccd1 vccd1 net1264 sky130_fd_sc_hd__clkbuf_4
X_16804_ ag2.body\[68\] net963 vssd1 vssd1 vccd1 vccd1 _02483_ sky130_fd_sc_hd__xor2_1
Xfanout1275 net1287 vssd1 vssd1 vccd1 vccd1 net1275 sky130_fd_sc_hd__buf_2
XFILLER_0_59_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10132__A net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1286 net1287 vssd1 vssd1 vccd1 vccd1 net1286 sky130_fd_sc_hd__clkbuf_2
X_17784_ obsg2.obstacleFlag _03461_ _03460_ vssd1 vssd1 vccd1 vccd1 _03462_ sky130_fd_sc_hd__o21ai_1
Xfanout1297 net1311 vssd1 vssd1 vccd1 vccd1 net1297 sky130_fd_sc_hd__clkbuf_4
X_14996_ net2656 net151 _01551_ control.body\[994\] vssd1 vssd1 vccd1 vccd1 _00332_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__13110__A1 net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19523_ clknet_leaf_121_clk _00467_ net1401 vssd1 vssd1 vccd1 vccd1 control.body\[865\]
+ sky130_fd_sc_hd__dfrtp_1
X_13947_ ag2.body\[88\] net190 _08155_ ag2.body\[80\] vssd1 vssd1 vccd1 vccd1 _00169_
+ sky130_fd_sc_hd__a22o_1
X_16735_ _02411_ _02413_ net499 vssd1 vssd1 vccd1 vccd1 _02414_ sky130_fd_sc_hd__mux2_1
XANTENNA__17388__B1 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14539__A net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12985__C _07508_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15938__A1 ag2.body\[160\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16666_ net396 _02342_ _02344_ net360 vssd1 vssd1 vccd1 vccd1 _02345_ sky130_fd_sc_hd__a211o_1
X_19454_ clknet_leaf_110_clk _00398_ net1419 vssd1 vssd1 vccd1 vccd1 control.body\[940\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11672__A1 net1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13878_ ag2.body\[27\] net121 _08147_ ag2.body\[19\] vssd1 vssd1 vccd1 vccd1 _00108_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_53_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15617_ ag2.body\[450\] net123 _01613_ ag2.body\[442\] vssd1 vssd1 vccd1 vccd1 _00884_
+ sky130_fd_sc_hd__a22o_1
X_18405_ _03890_ _03828_ vssd1 vssd1 vccd1 vccd1 _03895_ sky130_fd_sc_hd__nand2b_1
X_12829_ _07431_ _07615_ vssd1 vssd1 vccd1 vccd1 _07616_ sky130_fd_sc_hd__nor2_1
XFILLER_0_5_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16597_ obsg2.obstacleArray\[76\] obsg2.obstacleArray\[77\] _02214_ vssd1 vssd1 vccd1
+ vccd1 _02276_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19385_ clknet_leaf_93_clk _00329_ net1436 vssd1 vssd1 vccd1 vccd1 control.body\[1015\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09617__B2 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14610__B2 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18336_ _08139_ _03830_ vssd1 vssd1 vccd1 vccd1 _03832_ sky130_fd_sc_hd__nand2_1
X_15548_ ag2.body\[518\] net188 _01580_ ag2.body\[510\] vssd1 vssd1 vccd1 vccd1 _00824_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_127_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_96_3245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11975__A2 net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19284__CLK clknet_leaf_98_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_96_3256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18267_ net516 _03772_ vssd1 vssd1 vccd1 vccd1 _01381_ sky130_fd_sc_hd__nor2_1
XFILLER_0_115_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16363__A1 net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15479_ _06371_ net54 vssd1 vssd1 vccd1 vccd1 _01605_ sky130_fd_sc_hd__nor2_2
XFILLER_0_21_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17218_ _02893_ _02896_ _02884_ vssd1 vssd1 vccd1 vccd1 _02897_ sky130_fd_sc_hd__o21a_1
XFILLER_0_112_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18198_ _03543_ net36 vssd1 vssd1 vccd1 vccd1 _03738_ sky130_fd_sc_hd__nor2_1
XFILLER_0_31_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14913__A2 net171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20261__CLK clknet_leaf_43_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12506__B net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold703 control.body\[702\] vssd1 vssd1 vccd1 vccd1 net2265 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11727__A2 net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16115__A1 _01742_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold714 control.body\[856\] vssd1 vssd1 vccd1 vccd1 net2276 sky130_fd_sc_hd__dlygate4sd3_1
X_17149_ ag2.body\[609\] net868 vssd1 vssd1 vccd1 vccd1 _02828_ sky130_fd_sc_hd__nand2_1
XANTENNA__10307__A net1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold725 control.body\[782\] vssd1 vssd1 vccd1 vccd1 net2287 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_879 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold736 control.body\[1054\] vssd1 vssd1 vccd1 vccd1 net2298 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10935__B1 _05907_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold747 control.body\[635\] vssd1 vssd1 vccd1 vccd1 net2309 sky130_fd_sc_hd__dlygate4sd3_1
Xhold758 _00269_ vssd1 vssd1 vccd1 vccd1 net2320 sky130_fd_sc_hd__dlygate4sd3_1
X_20160_ clknet_leaf_101_clk _01104_ net1439 vssd1 vssd1 vccd1 vccd1 ag2.body\[238\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_126_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold769 control.body\[837\] vssd1 vssd1 vccd1 vccd1 net2331 sky130_fd_sc_hd__dlygate4sd3_1
X_09971_ net639 _04427_ vssd1 vssd1 vccd1 vccd1 _04944_ sky130_fd_sc_hd__nand2_2
XANTENNA__19882__RESET_B net1480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10026__B net1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkload27_A clknet_leaf_132_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20091_ clknet_leaf_78_clk _01035_ net1490 vssd1 vssd1 vccd1 vccd1 ag2.body\[297\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_42_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12152__A2 net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13337__B _07508_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout192_A net218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15626__B1 _01621_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_1115 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11138__A _05152_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17091__A2 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09831__A net1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_323 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10977__A net1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14449__A net975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout457_A net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_2802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1199_A net1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13353__A net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_2201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_2212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_2223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09405_ net272 _04342_ _04386_ vssd1 vssd1 vccd1 vccd1 _01400_ sky130_fd_sc_hd__nor3_1
XANTENNA_fanout245_X net245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout624_A net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1366_A net1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09336_ _04334_ net1889 vssd1 vssd1 vccd1 vccd1 _01428_ sky130_fd_sc_hd__nor2_1
XFILLER_0_34_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17479__B net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_510 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_2720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout412_X net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_2731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09267_ sound_gen.osc1.stayCount\[8\] _04289_ sound_gen.osc1.stayCount\[10\] sound_gen.osc1.stayCount\[9\]
+ vssd1 vssd1 vccd1 vccd1 _04290_ sky130_fd_sc_hd__o211a_1
XFILLER_0_84_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_79_2742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_141_clk clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_141_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_63_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1154_X net1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_2606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_2617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09198_ ag2.body\[618\] vssd1 vssd1 vccd1 vccd1 _04223_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout993_A net994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_2016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12915__A1 net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11320__B net1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_2027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20427_ clknet_leaf_37_clk _01314_ net1353 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[63\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__16106__A1 net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_2038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17303__B1 net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_120 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17926__C _03558_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16657__A2 net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11160_ ag2.body\[601\] net1196 vssd1 vssd1 vccd1 vccd1 _06133_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout781_X net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20358_ clknet_leaf_18_clk _01249_ net1324 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleCount\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14668__A1 net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14668__B2 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout879_X net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10111_ net1180 control.body\[938\] vssd1 vssd1 vccd1 vccd1 _05084_ sky130_fd_sc_hd__or2_1
XFILLER_0_105_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_8_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11091_ _06052_ _06057_ _06059_ _06063_ vssd1 vssd1 vccd1 vccd1 _06064_ sky130_fd_sc_hd__nor4_1
X_20289_ clknet_leaf_35_clk control.divider.next_count\[10\] net1350 vssd1 vssd1 vccd1
+ vccd1 control.divider.count\[10\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_105_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09725__B net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16409__A2 _02059_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10042_ _05011_ _05012_ _05013_ _05014_ vssd1 vssd1 vccd1 vccd1 _05015_ sky130_fd_sc_hd__or4_1
XANTENNA__13340__A1 net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09544__B1 net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13247__B net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold30 img_gen.tracker.frame\[520\] vssd1 vssd1 vccd1 vccd1 net1592 sky130_fd_sc_hd__dlygate4sd3_1
Xhold41 sound_gen.osc1.stayCount\[2\] vssd1 vssd1 vccd1 vccd1 net1603 sky130_fd_sc_hd__dlygate4sd3_1
X_14850_ _08784_ _08787_ _08792_ _08292_ _08191_ vssd1 vssd1 vccd1 vccd1 _01521_ sky130_fd_sc_hd__o311a_1
Xhold52 img_gen.tracker.frame\[190\] vssd1 vssd1 vccd1 vccd1 net1614 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout60_X net60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold63 img_gen.tracker.frame\[88\] vssd1 vssd1 vccd1 vccd1 net1625 sky130_fd_sc_hd__dlygate4sd3_1
Xhold74 img_gen.tracker.frame\[124\] vssd1 vssd1 vccd1 vccd1 net1636 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_610 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold85 img_gen.tracker.frame\[330\] vssd1 vssd1 vccd1 vccd1 net1647 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_118_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13801_ net677 _08104_ vssd1 vssd1 vccd1 vccd1 _08105_ sky130_fd_sc_hd__nor2_1
Xhold96 img_gen.tracker.frame\[10\] vssd1 vssd1 vccd1 vccd1 net1658 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14781_ net1020 ag2.body\[278\] vssd1 vssd1 vccd1 vccd1 _01452_ sky130_fd_sc_hd__or2_1
XANTENNA__11103__B1 net1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10887__A net1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11993_ img_gen.tracker.frame\[409\] net616 net545 img_gen.tracker.frame\[415\] vssd1
+ vssd1 vccd1 vccd1 _06965_ sky130_fd_sc_hd__o22a_1
X_16520_ _02152_ _02169_ _02057_ vssd1 vssd1 vccd1 vccd1 _02199_ sky130_fd_sc_hd__mux2_1
XANTENNA__13263__A net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13732_ img_gen.updater.commands.mode\[1\] _07224_ vssd1 vssd1 vccd1 vccd1 _08056_
+ sky130_fd_sc_hd__nand2_1
Xclkbuf_4_10__f_clk clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_10__leaf_clk
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__09460__B net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10944_ _04098_ net1164 net1091 _04100_ _05911_ vssd1 vssd1 vccd1 vccd1 _05917_ sky130_fd_sc_hd__a221o_1
X_16451_ obsg2.obstacleArray\[82\] obsg2.obstacleArray\[83\] net458 vssd1 vssd1 vccd1
+ vccd1 _02130_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13663_ net972 _08014_ vssd1 vssd1 vccd1 vccd1 _08017_ sky130_fd_sc_hd__or2_1
XFILLER_0_38_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10875_ ag2.body\[531\] net1158 vssd1 vssd1 vccd1 vccd1 _05848_ sky130_fd_sc_hd__or2_1
X_15402_ control.body\[643\] net82 _01581_ net2309 vssd1 vssd1 vccd1 vccd1 _00693_
+ sky130_fd_sc_hd__a22o_1
X_19170_ clknet_leaf_53_clk _00114_ net1365 vssd1 vssd1 vccd1 vccd1 ag2.body\[33\]
+ sky130_fd_sc_hd__dfrtp_4
X_12614_ net341 net332 net308 _07508_ vssd1 vssd1 vccd1 vccd1 _07509_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_26_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16382_ net493 _02053_ vssd1 vssd1 vccd1 vccd1 _02061_ sky130_fd_sc_hd__nand2_2
XFILLER_0_27_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13594_ control.divider.count\[10\] _07954_ _07967_ _07968_ vssd1 vssd1 vccd1 vccd1
+ _07969_ sky130_fd_sc_hd__a211o_1
XFILLER_0_87_1300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18121_ net352 _03635_ vssd1 vssd1 vccd1 vccd1 _03696_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_22_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15333_ net2222 net72 _01587_ control.body\[701\] vssd1 vssd1 vccd1 vccd1 _00631_
+ sky130_fd_sc_hd__a22o_1
X_12545_ net1934 net652 _07469_ _07470_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[32\]
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_54_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_132_clk clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_132_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__12607__A net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13159__A1 net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18052_ net301 _03566_ net39 obsg2.obstacleArray\[37\] vssd1 vssd1 vccd1 vccd1 _03651_
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_48_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15264_ _04604_ net54 vssd1 vssd1 vccd1 vccd1 _01582_ sky130_fd_sc_hd__nor2_2
X_12476_ net382 net308 vssd1 vssd1 vccd1 vccd1 _07431_ sky130_fd_sc_hd__nand2_8
XFILLER_0_22_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17003_ ag2.body\[141\] net708 net944 _04039_ _02681_ vssd1 vssd1 vccd1 vccd1 _02682_
+ sky130_fd_sc_hd__o221a_1
XANTENNA__12906__A1 net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14215_ net973 ag2.body\[411\] vssd1 vssd1 vccd1 vccd1 _08376_ sky130_fd_sc_hd__xnor2_1
X_11427_ ag2.body\[399\] net1056 vssd1 vssd1 vccd1 vccd1 _06400_ sky130_fd_sc_hd__nand2_1
XFILLER_0_111_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_5 _03442_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_1502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14381__X _08542_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15195_ net2531 net94 _01573_ control.body\[819\] vssd1 vssd1 vccd1 vccd1 _00509_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_39_1513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10127__A net1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14146_ net970 ag2.body\[595\] vssd1 vssd1 vccd1 vccd1 _08307_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_1_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11358_ net900 _04238_ _04554_ _05075_ _04491_ vssd1 vssd1 vccd1 vccd1 _06331_ sky130_fd_sc_hd__a41o_1
XFILLER_0_123_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18013__B net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10309_ net1218 control.body\[696\] vssd1 vssd1 vccd1 vccd1 _05282_ sky130_fd_sc_hd__xor2_1
XANTENNA__10414__X _05387_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18954_ clknet_leaf_5_clk img_gen.tracker.next_frame\[392\] net1276 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[392\] sky130_fd_sc_hd__dfrtp_1
X_14077_ net1025 ag2.body\[565\] vssd1 vssd1 vccd1 vccd1 _08238_ sky130_fd_sc_hd__xor2_1
XANTENNA__12342__A net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11289_ net1137 control.body\[1108\] vssd1 vssd1 vccd1 vccd1 _06262_ sky130_fd_sc_hd__or2_1
XFILLER_0_67_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12134__A2 net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17905_ _03533_ _03538_ vssd1 vssd1 vccd1 vccd1 _03540_ sky130_fd_sc_hd__nor2_2
X_13028_ net238 _07708_ _07709_ net1975 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[276\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__10145__A1 _04238_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18885_ clknet_leaf_11_clk img_gen.tracker.next_frame\[323\] net1283 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[323\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__15608__B1 _01620_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1050 net1051 vssd1 vssd1 vccd1 vccd1 net1050 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__13725__X toggle1.nextDisplayOut\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1061 net1062 vssd1 vssd1 vccd1 vccd1 net1061 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10696__A2 _05657_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17836_ net1026 ag2.apple_cord\[5\] _03489_ vssd1 vssd1 vccd1 vccd1 _03495_ sky130_fd_sc_hd__mux2_1
Xfanout1072 net1074 vssd1 vssd1 vccd1 vccd1 net1072 sky130_fd_sc_hd__clkbuf_4
XANTENNA__16101__X _01780_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1083 net1084 vssd1 vssd1 vccd1 vccd1 net1083 sky130_fd_sc_hd__clkbuf_4
Xfanout1094 net1095 vssd1 vssd1 vccd1 vccd1 net1094 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_83_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09651__A net1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16820__A2 net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15372__B _01581_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17767_ _02902_ _02907_ _03187_ vssd1 vssd1 vccd1 vccd1 _03446_ sky130_fd_sc_hd__o21a_2
XANTENNA__14269__A net1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14979_ control.body\[1018\] net151 _01550_ net2371 vssd1 vssd1 vccd1 vccd1 _00316_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_117_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19506_ clknet_leaf_121_clk _00450_ net1402 vssd1 vssd1 vccd1 vccd1 control.body\[880\]
+ sky130_fd_sc_hd__dfrtp_1
X_16718_ _02394_ _02396_ net495 vssd1 vssd1 vccd1 vccd1 _02397_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_1068 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17698_ obsg2.obstacleArray\[130\] obsg2.obstacleArray\[131\] obsg2.obstacleArray\[134\]
+ obsg2.obstacleArray\[135\] net410 net370 vssd1 vssd1 vccd1 vccd1 _03377_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_18_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19437_ clknet_leaf_108_clk _00381_ net1422 vssd1 vssd1 vccd1 vccd1 control.body\[955\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11405__B net1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_98_3307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16649_ _02326_ _02327_ net396 vssd1 vssd1 vccd1 vccd1 _02328_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_18_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_3318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17781__B1 _03457_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13398__A1 net238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17299__B net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19368_ clknet_leaf_94_clk net2555 net1439 vssd1 vssd1 vccd1 vccd1 control.body\[1030\]
+ sky130_fd_sc_hd__dfrtp_1
X_09121_ ag2.body\[406\] vssd1 vssd1 vccd1 vccd1 _04146_ sky130_fd_sc_hd__inv_2
XANTENNA__14716__B ag2.body\[339\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11948__A2 net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18319_ _08138_ _03814_ vssd1 vssd1 vccd1 vccd1 _03815_ sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_123_clk clknet_4_9__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_123_clk
+ sky130_fd_sc_hd__clkbuf_8
X_19299_ clknet_leaf_99_clk _00243_ net1445 vssd1 vssd1 vccd1 vccd1 control.body\[1089\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__17533__B1 net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11421__A net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09052_ ag2.body\[245\] vssd1 vssd1 vccd1 vccd1 _04077_ sky130_fd_sc_hd__inv_2
XFILLER_0_72_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_854 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11140__B net1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold500 img_gen.tracker.frame\[166\] vssd1 vssd1 vccd1 vccd1 net2062 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_114_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14732__A net993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold511 img_gen.tracker.frame\[33\] vssd1 vssd1 vccd1 vccd1 net2073 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout205_A net210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold522 img_gen.tracker.frame\[27\] vssd1 vssd1 vccd1 vccd1 net2084 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold533 img_gen.tracker.frame\[538\] vssd1 vssd1 vccd1 vccd1 net2095 sky130_fd_sc_hd__dlygate4sd3_1
X_20212_ clknet_leaf_60_clk _01156_ net1466 vssd1 vssd1 vccd1 vccd1 ag2.body\[178\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__09826__A net1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold544 img_gen.tracker.frame\[559\] vssd1 vssd1 vccd1 vccd1 net2106 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold555 sound_gen.dac1.dacCount\[4\] vssd1 vssd1 vccd1 vccd1 net2117 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold566 img_gen.tracker.frame\[555\] vssd1 vssd1 vccd1 vccd1 net2128 sky130_fd_sc_hd__dlygate4sd3_1
Xhold577 img_gen.updater.commands.rR1.rainbowRNG\[7\] vssd1 vssd1 vccd1 vccd1 net2139
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold588 control.body\[904\] vssd1 vssd1 vccd1 vccd1 net2150 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13348__A net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20143_ clknet_leaf_96_clk _01087_ net1451 vssd1 vssd1 vccd1 vccd1 ag2.body\[253\]
+ sky130_fd_sc_hd__dfrtp_4
X_09954_ net777 control.body\[737\] control.body\[742\] net748 vssd1 vssd1 vccd1 vccd1
+ _04927_ sky130_fd_sc_hd__o22ai_1
Xhold599 control.body\[770\] vssd1 vssd1 vccd1 vccd1 net2161 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1114_A net1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12125__A2 net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20074_ clknet_leaf_77_clk _01018_ net1491 vssd1 vssd1 vccd1 vccd1 ag2.body\[312\]
+ sky130_fd_sc_hd__dfrtp_2
X_09885_ _04847_ _04853_ _04855_ _04857_ vssd1 vssd1 vccd1 vccd1 _04858_ sky130_fd_sc_hd__or4b_2
XANTENNA_fanout574_A net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout195_X net195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_2410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16498__S1 net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16811__A2 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15282__B net55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout741_A _04262_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout362_X net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout839_A _03965_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14822__A1 net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1483_A net1484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14822__B2 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13083__A net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11636__A1 _06485_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_808 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout627_X net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1369_X net1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10660_ net640 _05051_ net636 vssd1 vssd1 vccd1 vccd1 _05633_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_119_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_1620 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11939__A2 net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09319_ _04319_ _04322_ _04333_ net272 sound_gen.osc1.count\[2\] vssd1 vssd1 vccd1
+ vccd1 _01437_ sky130_fd_sc_hd__a32o_1
XANTENNA__17524__B1 net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_114_clk clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_114_clk
+ sky130_fd_sc_hd__clkbuf_8
X_10591_ net1076 control.body\[830\] vssd1 vssd1 vccd1 vccd1 _05564_ sky130_fd_sc_hd__or2_1
XFILLER_0_49_1604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11331__A net1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12330_ _07256_ _07292_ _07296_ _07290_ vssd1 vssd1 vccd1 vccd1 _07297_ sky130_fd_sc_hd__a22o_1
XFILLER_0_49_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17496__Y _03175_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout996_X net996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16841__B net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12261_ img_gen.updater.commands.mode\[2\] img_gen.updater.commands.mode\[0\] img_gen.updater.commands.mode\[1\]
+ vssd1 vssd1 vccd1 vccd1 _07231_ sky130_fd_sc_hd__nor3b_1
XANTENNA__12714__X _07561_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15550__A2 _04944_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18114__A net44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14642__A net1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14000_ net844 ag2.body\[504\] ag2.body\[506\] net828 vssd1 vssd1 vccd1 vccd1 _08161_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_47_1361 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11212_ net1226 control.body\[840\] vssd1 vssd1 vccd1 vccd1 _06185_ sky130_fd_sc_hd__xnor2_1
X_12192_ net1054 ag2.apple_cord\[7\] vssd1 vssd1 vccd1 vccd1 _07164_ sky130_fd_sc_hd__or2_1
Xoutput20 net20 vssd1 vssd1 vccd1 vccd1 gpio_out[19] sky130_fd_sc_hd__buf_2
Xoutput31 net31 vssd1 vssd1 vccd1 vccd1 gpio_out[6] sky130_fd_sc_hd__buf_2
X_11143_ ag2.body\[413\] net1105 vssd1 vssd1 vccd1 vccd1 _06116_ sky130_fd_sc_hd__xor2_1
XANTENNA__09455__B net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12116__A2 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15951_ ag2.body\[156\] net196 _01656_ ag2.body\[148\] vssd1 vssd1 vccd1 vccd1 _01182_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_120_1459 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17672__B net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11074_ ag2.body\[362\] net776 net763 ag2.body\[364\] _06043_ vssd1 vssd1 vccd1 vccd1
+ _06047_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_37_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17055__A2 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10025_ ag2.body\[508\] net1138 vssd1 vssd1 vccd1 vccd1 _04998_ sky130_fd_sc_hd__xor2_1
X_14902_ net2199 net178 _01540_ control.body\[1087\] vssd1 vssd1 vccd1 vccd1 _00249_
+ sky130_fd_sc_hd__a22o_1
X_15882_ ag2.body\[223\] net188 _01648_ ag2.body\[215\] vssd1 vssd1 vccd1 vccd1 _01121_
+ sky130_fd_sc_hd__a22o_1
X_18670_ clknet_leaf_26_clk img_gen.tracker.next_frame\[108\] net1339 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[108\] sky130_fd_sc_hd__dfrtp_1
X_17621_ ag2.body\[191\] net929 vssd1 vssd1 vccd1 vccd1 _03300_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_95_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14833_ _08802_ _08804_ _08810_ _08315_ vssd1 vssd1 vccd1 vccd1 _01504_ sky130_fd_sc_hd__o31a_1
XANTENNA__14089__A net1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11627__A1 net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11506__A net1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17552_ ag2.body\[352\] net888 vssd1 vssd1 vccd1 vccd1 _03231_ sky130_fd_sc_hd__xor2_1
X_14764_ net1039 ag2.body\[100\] vssd1 vssd1 vccd1 vccd1 _08925_ sky130_fd_sc_hd__xor2_1
X_11976_ img_gen.tracker.frame\[565\] net622 net605 img_gen.tracker.frame\[568\] _06946_
+ vssd1 vssd1 vccd1 vccd1 _06948_ sky130_fd_sc_hd__o221a_1
XANTENNA__10410__A net1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16503_ obsg2.obstacleArray\[2\] obsg2.obstacleArray\[3\] net457 vssd1 vssd1 vccd1
+ vccd1 _02182_ sky130_fd_sc_hd__mux2_1
X_13715_ track.highScore\[4\] _08025_ net356 vssd1 vssd1 vccd1 vccd1 track.nextHighScore\[4\]
+ sky130_fd_sc_hd__mux2_1
X_17483_ ag2.body\[130\] net728 net934 _04035_ _03161_ vssd1 vssd1 vccd1 vccd1 _03162_
+ sky130_fd_sc_hd__a221o_1
XANTENNA__15920__B net57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10927_ net775 control.body\[1034\] _05899_ _04235_ vssd1 vssd1 vccd1 vccd1 _05900_
+ sky130_fd_sc_hd__a211oi_1
X_14695_ net845 ag2.body\[320\] _04111_ net1040 _08855_ vssd1 vssd1 vccd1 vccd1 _08856_
+ sky130_fd_sc_hd__a221o_1
XANTENNA__17763__B1 _03441_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19222_ clknet_leaf_67_clk _00166_ net1494 vssd1 vssd1 vccd1 vccd1 ag2.body\[85\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_89_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13721__A net26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13646_ control.divider.count\[15\] control.divider.count\[16\] _08001_ vssd1 vssd1
+ vccd1 vccd1 _08005_ sky130_fd_sc_hd__and3_1
X_16434_ obsg2.obstacleArray\[76\] obsg2.obstacleArray\[77\] net453 vssd1 vssd1 vccd1
+ vccd1 _02113_ sky130_fd_sc_hd__mux2_1
X_10858_ _05825_ _05828_ _05829_ _05830_ vssd1 vssd1 vccd1 vccd1 _05831_ sky130_fd_sc_hd__or4_1
XFILLER_0_39_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10850__A2 net1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11512__Y _06485_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16365_ obsg2.obstacleArray\[12\] net409 vssd1 vssd1 vccd1 vccd1 _02044_ sky130_fd_sc_hd__or2_1
X_19153_ clknet_leaf_52_clk _00097_ net1367 vssd1 vssd1 vccd1 vccd1 ag2.body\[17\]
+ sky130_fd_sc_hd__dfrtp_4
X_13577_ control.divider.count\[19\] control.divider.count\[18\] _07949_ vssd1 vssd1
+ vccd1 vccd1 _07952_ sky130_fd_sc_hd__and3_1
XFILLER_0_82_852 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_105_clk clknet_4_10__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_105_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_13_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12337__A _07301_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10789_ net1120 control.body\[628\] vssd1 vssd1 vccd1 vccd1 _05762_ sky130_fd_sc_hd__xor2_1
XANTENNA__17515__B1 net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18104_ net345 _03545_ _03573_ vssd1 vssd1 vccd1 vccd1 _03685_ sky130_fd_sc_hd__and3_1
X_15316_ net2626 net74 _01588_ net2421 vssd1 vssd1 vccd1 vccd1 _00615_ sky130_fd_sc_hd__a22o_1
XFILLER_0_48_1103 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12528_ net2165 net651 _07461_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[24\]
+ sky130_fd_sc_hd__and3_1
X_16296_ obsg2.obstacleArray\[115\] net413 _01974_ net415 vssd1 vssd1 vccd1 vccd1
+ _01975_ sky130_fd_sc_hd__o211a_1
XFILLER_0_54_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19084_ clknet_leaf_29_clk img_gen.tracker.next_frame\[522\] net1334 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[522\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_124_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18035_ _01714_ net345 net299 vssd1 vssd1 vccd1 vccd1 _03640_ sky130_fd_sc_hd__and3_1
X_15247_ net2594 net97 _01579_ net2243 vssd1 vssd1 vccd1 vccd1 _00555_ sky130_fd_sc_hd__a22o_1
X_20597__1529 vssd1 vssd1 vccd1 vccd1 _20597__1529/HI net1529 sky130_fd_sc_hd__conb_1
XANTENNA__16243__S net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12459_ _07223_ _07263_ _07270_ _07280_ _07275_ vssd1 vssd1 vccd1 vccd1 _07418_ sky130_fd_sc_hd__a221o_1
XANTENNA__14552__A net1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09646__A net1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15178_ net2588 net102 _01571_ control.body\[836\] vssd1 vssd1 vccd1 vccd1 _00494_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_61_1314 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15829__B1 _01643_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14129_ net843 ag2.body\[368\] _08281_ _08282_ _08289_ vssd1 vssd1 vccd1 vccd1 _08290_
+ sky130_fd_sc_hd__a221o_1
X_19986_ clknet_leaf_64_clk _00930_ net1474 vssd1 vssd1 vccd1 vccd1 ag2.body\[400\]
+ sky130_fd_sc_hd__dfrtp_4
Xfanout309 _07429_ vssd1 vssd1 vccd1 vccd1 net309 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09508__B1 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12107__A2 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18937_ clknet_leaf_139_clk img_gen.tracker.next_frame\[375\] net1288 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[375\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_103_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17046__A2 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09670_ _04635_ _04639_ _04642_ vssd1 vssd1 vccd1 vccd1 _04643_ sky130_fd_sc_hd__and3_1
X_18868_ clknet_leaf_26_clk img_gen.tracker.next_frame\[306\] net1342 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[306\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_118_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17819_ _03476_ _03485_ net924 _03475_ vssd1 vssd1 vccd1 vccd1 _01221_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_55_1107 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18799_ clknet_leaf_18_clk img_gen.tracker.next_frame\[237\] net1319 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[237\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14804__B2 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11416__A net1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11618__A1 net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16422__B1_N _02057_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16926__B net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16557__A1 net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14286__X _08447_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14727__A net1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout155_A net162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1151 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17506__B1 net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1064_A net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_239 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09104_ ag2.body\[360\] vssd1 vssd1 vccd1 vccd1 _04129_ sky130_fd_sc_hd__inv_2
XANTENNA__13791__A1 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09035_ ag2.body\[193\] vssd1 vssd1 vccd1 vccd1 _04060_ sky130_fd_sc_hd__inv_2
XFILLER_0_5_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1231_A net1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_445 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold330 img_gen.tracker.frame\[341\] vssd1 vssd1 vccd1 vccd1 net1892 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__19144__RESET_B net1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold341 img_gen.tracker.frame\[55\] vssd1 vssd1 vccd1 vccd1 net1903 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout691_A net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold352 img_gen.tracker.frame\[505\] vssd1 vssd1 vccd1 vccd1 net1914 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold363 img_gen.tracker.frame\[200\] vssd1 vssd1 vccd1 vccd1 net1925 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold374 img_gen.tracker.frame\[29\] vssd1 vssd1 vccd1 vccd1 net1936 sky130_fd_sc_hd__dlygate4sd3_1
Xhold385 img_gen.tracker.frame\[506\] vssd1 vssd1 vccd1 vccd1 net1947 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold396 img_gen.tracker.frame\[313\] vssd1 vssd1 vccd1 vccd1 net1958 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout810 _03971_ vssd1 vssd1 vccd1 vccd1 net810 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_111_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1117_X net1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout821 net822 vssd1 vssd1 vccd1 vccd1 net821 sky130_fd_sc_hd__clkbuf_4
XANTENNA__20049__RESET_B net1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09937_ ag2.body\[29\] net1102 vssd1 vssd1 vccd1 vccd1 _04910_ sky130_fd_sc_hd__and2b_1
X_20126_ clknet_leaf_81_clk _01070_ net1486 vssd1 vssd1 vccd1 vccd1 ag2.body\[268\]
+ sky130_fd_sc_hd__dfrtp_4
Xfanout832 net836 vssd1 vssd1 vccd1 vccd1 net832 sky130_fd_sc_hd__clkbuf_4
Xfanout843 net847 vssd1 vssd1 vccd1 vccd1 net843 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout956_A net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout854 net857 vssd1 vssd1 vccd1 vccd1 net854 sky130_fd_sc_hd__buf_4
XANTENNA_fanout577_X net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout865 net867 vssd1 vssd1 vccd1 vccd1 net865 sky130_fd_sc_hd__buf_4
XFILLER_0_99_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout876 net877 vssd1 vssd1 vccd1 vccd1 net876 sky130_fd_sc_hd__buf_4
XANTENNA__17037__A2 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20057_ clknet_leaf_72_clk _01001_ net1502 vssd1 vssd1 vccd1 vccd1 ag2.body\[343\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__13806__A net1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout887 net888 vssd1 vssd1 vccd1 vccd1 net887 sky130_fd_sc_hd__clkbuf_4
X_09868_ ag2.body\[152\] net1234 vssd1 vssd1 vccd1 vccd1 _04841_ sky130_fd_sc_hd__xor2_1
XANTENNA__12710__A net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1030 control.body\[907\] vssd1 vssd1 vccd1 vccd1 net2592 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout898 net899 vssd1 vssd1 vccd1 vccd1 net898 sky130_fd_sc_hd__buf_2
Xhold1041 control.body\[915\] vssd1 vssd1 vccd1 vccd1 net2603 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1052 control.body\[885\] vssd1 vssd1 vccd1 vccd1 net2614 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_77_1376 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1063 control.body\[640\] vssd1 vssd1 vccd1 vccd1 net2625 sky130_fd_sc_hd__dlygate4sd3_1
X_09799_ net893 _04519_ net636 vssd1 vssd1 vccd1 vccd1 _04772_ sky130_fd_sc_hd__o21a_2
Xhold1074 control.body\[657\] vssd1 vssd1 vccd1 vccd1 net2636 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout744_X net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17993__B1 net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1085 control.body\[652\] vssd1 vssd1 vccd1 vccd1 net2647 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11609__A1 net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11830_ img_gen.tracker.frame\[542\] net613 net596 img_gen.tracker.frame\[545\] vssd1
+ vssd1 vccd1 vccd1 _06802_ sky130_fd_sc_hd__o22a_1
Xhold1096 control.body\[695\] vssd1 vssd1 vccd1 vccd1 net2658 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16836__B net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15740__B net60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11761_ img_gen.tracker.frame\[269\] net604 net587 img_gen.tracker.frame\[275\] vssd1
+ vssd1 vccd1 vccd1 _06733_ sky130_fd_sc_hd__o22a_1
XANTENNA__16328__S net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13500_ _07607_ net304 vssd1 vssd1 vccd1 vccd1 _07912_ sky130_fd_sc_hd__nor2_1
XFILLER_0_95_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10712_ net898 _05161_ net891 vssd1 vssd1 vccd1 vccd1 _05685_ sky130_fd_sc_hd__a21o_2
XFILLER_0_138_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14480_ net972 ag2.body\[443\] vssd1 vssd1 vccd1 vccd1 _08641_ sky130_fd_sc_hd__xor2_1
X_11692_ img_gen.tracker.frame\[104\] net546 _06663_ net562 vssd1 vssd1 vccd1 vccd1
+ _06664_ sky130_fd_sc_hd__o211a_1
XFILLER_0_126_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_3__f_clk_X clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13431_ net682 _07884_ vssd1 vssd1 vccd1 vccd1 _07885_ sky130_fd_sc_hd__nor2_1
XFILLER_0_10_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10643_ _04603_ _04791_ vssd1 vssd1 vccd1 vccd1 _05616_ sky130_fd_sc_hd__nor2_1
XFILLER_0_125_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15771__A2 net210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16150_ obsg2.obstacleArray\[20\] net429 net375 _01828_ vssd1 vssd1 vccd1 vccd1 _01829_
+ sky130_fd_sc_hd__o211a_1
X_13362_ net314 _07528_ vssd1 vssd1 vccd1 vccd1 _07858_ sky130_fd_sc_hd__and2_1
XANTENNA__17667__B net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10574_ ag2.body\[190\] net1080 vssd1 vssd1 vccd1 vccd1 _05547_ sky130_fd_sc_hd__nand2_1
XFILLER_0_107_976 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_5_clk_A clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11793__B1 net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15101_ control.body\[919\] net145 _01563_ net2110 vssd1 vssd1 vccd1 vccd1 _00425_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_2_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12313_ _07279_ vssd1 vssd1 vccd1 vccd1 _07280_ sky130_fd_sc_hd__inv_2
X_16081_ obsg2.obstacleArray\[96\] obsg2.obstacleArray\[97\] net421 vssd1 vssd1 vccd1
+ vccd1 _01760_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13293_ _07476_ net303 vssd1 vssd1 vccd1 vccd1 _07831_ sky130_fd_sc_hd__nor2_1
XANTENNA__14372__A net1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20322__CLK clknet_leaf_43_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15032_ net2236 net163 _01557_ net2312 vssd1 vssd1 vccd1 vccd1 _00362_ sky130_fd_sc_hd__a22o_1
XFILLER_0_121_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12244_ img_gen.updater.commands.count\[16\] _07213_ vssd1 vssd1 vccd1 vccd1 _07214_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_82_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11545__B1 net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19495__CLK clknet_leaf_113_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19840_ clknet_leaf_122_clk _00784_ net1414 vssd1 vssd1 vccd1 vccd1 ag2.body\[558\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_48_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12175_ _07039_ _07093_ _07145_ _07146_ vssd1 vssd1 vccd1 vccd1 _07147_ sky130_fd_sc_hd__a22oi_4
XANTENNA__18131__X _03702_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10405__A net1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16484__B1 net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1234 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__20401__RESET_B net1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11126_ control.body\[868\] net1131 vssd1 vssd1 vccd1 vccd1 _06099_ sky130_fd_sc_hd__and2b_1
X_19771_ clknet_leaf_19_clk _00715_ net1322 vssd1 vssd1 vccd1 vccd1 ag2.body\[617\]
+ sky130_fd_sc_hd__dfrtp_4
X_16983_ _02659_ _02660_ _02661_ vssd1 vssd1 vccd1 vccd1 _02662_ sky130_fd_sc_hd__and3_1
XFILLER_0_120_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18722_ clknet_leaf_142_clk img_gen.tracker.next_frame\[160\] net1253 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[160\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__09472__Y _04445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09913__B net1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11057_ ag2.body\[432\] net1224 vssd1 vssd1 vccd1 vccd1 _06030_ sky130_fd_sc_hd__xnor2_1
X_15934_ ag2.body\[172\] net136 _01655_ ag2.body\[164\] vssd1 vssd1 vccd1 vccd1 _01166_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12620__A net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_1454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10008_ net742 net923 _04980_ vssd1 vssd1 vccd1 vccd1 _04981_ sky130_fd_sc_hd__and3_1
X_18653_ clknet_leaf_131_clk img_gen.tracker.next_frame\[91\] net1317 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[91\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__10520__A1 _04421_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15865_ _05517_ net66 vssd1 vssd1 vccd1 vccd1 _01647_ sky130_fd_sc_hd__and2_2
X_17604_ _04150_ net961 net697 ag2.body\[422\] _03282_ vssd1 vssd1 vccd1 vccd1 _03283_
+ sky130_fd_sc_hd__a221o_1
X_14816_ net982 _04134_ _01485_ _01486_ _01484_ vssd1 vssd1 vccd1 vccd1 _01487_ sky130_fd_sc_hd__a221o_1
XANTENNA__10140__A net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18584_ clknet_leaf_14_clk img_gen.tracker.next_frame\[22\] net1278 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[22\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15796_ ag2.body\[289\] net205 _01640_ ag2.body\[281\] vssd1 vssd1 vccd1 vccd1 _01043_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_86_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15650__B net57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11076__A2 net1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_292 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17535_ ag2.body\[272\] net740 net864 _04093_ vssd1 vssd1 vccd1 vccd1 _03214_ sky130_fd_sc_hd__a2bb2o_1
X_14747_ net1023 ag2.body\[110\] vssd1 vssd1 vccd1 vccd1 _08908_ sky130_fd_sc_hd__xor2_1
X_11959_ _06876_ _06930_ net387 vssd1 vssd1 vccd1 vccd1 _06931_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17736__B1 _02703_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14547__A net975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18019__A net45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13451__A net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17200__A2 net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14678_ net818 ag2.body\[387\] ag2.body\[390\] net801 vssd1 vssd1 vccd1 vccd1 _08839_
+ sky130_fd_sc_hd__a22o_1
X_17466_ _03141_ _03142_ _03143_ _03144_ vssd1 vssd1 vccd1 vccd1 _03145_ sky130_fd_sc_hd__or4_1
XANTENNA__10794__B net1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19205_ clknet_leaf_86_clk _00149_ net1459 vssd1 vssd1 vccd1 vccd1 ag2.body\[68\]
+ sky130_fd_sc_hd__dfrtp_4
X_13629_ control.divider.count\[10\] _07992_ net222 vssd1 vssd1 vccd1 vccd1 _07994_
+ sky130_fd_sc_hd__o21ai_1
X_16417_ net398 _02095_ vssd1 vssd1 vccd1 vccd1 _02096_ sky130_fd_sc_hd__or2_1
XFILLER_0_89_1269 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17397_ ag2.body\[509\] net952 vssd1 vssd1 vccd1 vccd1 _03076_ sky130_fd_sc_hd__xor2_1
XFILLER_0_82_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19136_ clknet_leaf_132_clk img_gen.tracker.next_frame\[574\] net1297 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[574\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__09928__X _04901_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16348_ _02023_ _02026_ net371 vssd1 vssd1 vccd1 vccd1 _02027_ sky130_fd_sc_hd__mux2_1
XANTENNA__14970__B1 net51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11784__B1 net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_1545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18712__CLK clknet_leaf_144_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16279_ obsg2.obstacleArray\[16\] obsg2.obstacleArray\[17\] net412 vssd1 vssd1 vccd1
+ vccd1 _01958_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19067_ clknet_leaf_29_clk img_gen.tracker.next_frame\[505\] net1334 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[505\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_120_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18018_ net299 _03627_ vssd1 vssd1 vccd1 vccd1 _03628_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_114_3793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12514__B net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12879__A3 _07638_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_3668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_3679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17267__A2 net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout106 net107 vssd1 vssd1 vccd1 vccd1 net106 sky130_fd_sc_hd__clkbuf_2
Xfanout117 net128 vssd1 vssd1 vccd1 vccd1 net117 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__16475__B1 net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19988__CLK clknet_leaf_66_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20142__RESET_B net1451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout128 net219 vssd1 vssd1 vccd1 vccd1 net128 sky130_fd_sc_hd__buf_2
XFILLER_0_129_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_487 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout139 net144 vssd1 vssd1 vccd1 vccd1 net139 sky130_fd_sc_hd__buf_2
X_19969_ clknet_leaf_62_clk _00913_ net1469 vssd1 vssd1 vccd1 vccd1 ag2.body\[431\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA_clkbuf_4_14__f_clk_X clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09722_ net909 _04637_ vssd1 vssd1 vccd1 vccd1 _04695_ sky130_fd_sc_hd__and2_4
XFILLER_0_39_1603 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09653_ net1098 control.body\[749\] vssd1 vssd1 vccd1 vccd1 _04626_ sky130_fd_sc_hd__xor2_1
XFILLER_0_39_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_2_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_1095 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10050__A _04931_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09584_ _04555_ _04556_ _04553_ vssd1 vssd1 vccd1 vccd1 _04557_ sky130_fd_sc_hd__o21a_1
XFILLER_0_132_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_118_Right_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16656__B net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15560__B net61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10985__A net1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout537_A _01707_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1181_A net1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1279_A net1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09680__A2 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_446 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout704_A net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10049__X _05022_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1067_X net1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14961__B1 _01547_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11775__B1 net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1618 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14192__A net1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15505__A2 net113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1234_X net1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09018_ ag2.body\[149\] vssd1 vssd1 vccd1 vccd1 _04043_ sky130_fd_sc_hd__inv_2
XFILLER_0_20_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14713__B1 ag2.body\[340\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10290_ ag2.body\[334\] net1090 vssd1 vssd1 vccd1 vccd1 _05263_ sky130_fd_sc_hd__or2_1
XFILLER_0_130_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout694_X net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20495__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold160 img_gen.tracker.frame\[78\] vssd1 vssd1 vccd1 vccd1 net1722 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__16611__S net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold171 img_gen.tracker.frame\[435\] vssd1 vssd1 vccd1 vccd1 net1733 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold182 img_gen.tracker.frame\[391\] vssd1 vssd1 vccd1 vccd1 net1744 sky130_fd_sc_hd__dlygate4sd3_1
Xhold193 control.fsm.temp\[0\] vssd1 vssd1 vccd1 vccd1 net1755 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout861_X net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout959_X net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout640 _04426_ vssd1 vssd1 vccd1 vccd1 net640 sky130_fd_sc_hd__clkbuf_4
Xfanout651 net653 vssd1 vssd1 vccd1 vccd1 net651 sky130_fd_sc_hd__buf_2
Xfanout662 net663 vssd1 vssd1 vccd1 vccd1 net662 sky130_fd_sc_hd__clkbuf_4
X_20109_ clknet_leaf_79_clk _01053_ net1487 vssd1 vssd1 vccd1 vccd1 ag2.body\[283\]
+ sky130_fd_sc_hd__dfrtp_4
X_13980_ ag2.body\[118\] net203 _08158_ ag2.body\[110\] vssd1 vssd1 vccd1 vccd1 _00199_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__09733__B net1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout673 net674 vssd1 vssd1 vccd1 vccd1 net673 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10879__B net1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout684 _04393_ vssd1 vssd1 vccd1 vccd1 net684 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09499__A2 _04471_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout695 _04269_ vssd1 vssd1 vccd1 vccd1 net695 sky130_fd_sc_hd__buf_6
X_12931_ net244 _07662_ _07663_ net1598 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[225\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__09452__C net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15650_ _05152_ net57 vssd1 vssd1 vccd1 vccd1 _01624_ sky130_fd_sc_hd__nor2_2
X_12862_ net261 _07631_ _07632_ net1771 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[187\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_34_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20596__1528 vssd1 vssd1 vccd1 vccd1 _20596__1528/HI net1528 sky130_fd_sc_hd__conb_1
XFILLER_0_38_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14601_ _08759_ _08760_ _08761_ vssd1 vssd1 vccd1 vccd1 _08762_ sky130_fd_sc_hd__or3_1
X_11813_ img_gen.tracker.frame\[479\] net578 net540 img_gen.tracker.frame\[476\] vssd1
+ vssd1 vccd1 vccd1 _06785_ sky130_fd_sc_hd__o22a_1
X_15581_ ag2.body\[481\] net130 _01617_ ag2.body\[473\] vssd1 vssd1 vccd1 vccd1 _00851_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__15470__B net54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12793_ net231 _07599_ _07600_ net1920 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[150\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_69_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14532_ _08689_ _08690_ _08691_ _08692_ vssd1 vssd1 vccd1 vccd1 _08693_ sky130_fd_sc_hd__a22o_1
X_17320_ ag2.body\[216\] net886 vssd1 vssd1 vccd1 vccd1 _02999_ sky130_fd_sc_hd__xor2_1
X_11744_ img_gen.tracker.frame\[2\] net623 net565 _06715_ vssd1 vssd1 vccd1 vccd1
+ _06716_ sky130_fd_sc_hd__o211a_1
XFILLER_0_68_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_4494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14463_ net1038 ag2.body\[268\] vssd1 vssd1 vccd1 vccd1 _08624_ sky130_fd_sc_hd__xor2_1
XANTENNA__11503__B net1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17251_ ag2.body\[549\] net947 vssd1 vssd1 vccd1 vccd1 _02930_ sky130_fd_sc_hd__xor2_1
X_11675_ _06638_ _06640_ vssd1 vssd1 vccd1 vccd1 _06647_ sky130_fd_sc_hd__xnor2_4
XANTENNA__16582__A _01700_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10018__B1 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16202_ _01879_ _01880_ net376 vssd1 vssd1 vccd1 vccd1 _01881_ sky130_fd_sc_hd__mux2_1
X_13414_ net280 _07876_ _07877_ net2041 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[494\]
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_133_4369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17182_ _02856_ _02858_ _02859_ _02860_ vssd1 vssd1 vccd1 vccd1 _02861_ sky130_fd_sc_hd__or4_1
XANTENNA__14952__B1 _01546_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10626_ _05593_ _05594_ _05596_ _05597_ vssd1 vssd1 vccd1 vccd1 _05599_ sky130_fd_sc_hd__a22o_1
X_14394_ net1003 _04028_ ag2.body\[122\] net829 _08553_ vssd1 vssd1 vccd1 vccd1 _08555_
+ sky130_fd_sc_hd__a221o_1
XANTENNA__17397__B net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16133_ _01785_ _01794_ _01802_ _01811_ vssd1 vssd1 vccd1 vccd1 _01812_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_12_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13345_ net249 _07850_ _07851_ net1762 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[451\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_64_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10557_ ag2.body\[517\] net1108 vssd1 vssd1 vccd1 vccd1 _05530_ sky130_fd_sc_hd__xor2_1
XANTENNA__09908__B net1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12615__A net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13507__A1 net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16064_ _01727_ _01741_ vssd1 vssd1 vccd1 vccd1 _01743_ sky130_fd_sc_hd__nand2_4
XFILLER_0_49_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13276_ net255 _07823_ _07824_ net1807 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[409\]
+ sky130_fd_sc_hd__a22o_1
X_10488_ ag2.body\[586\] net773 net1101 _04216_ _05460_ vssd1 vssd1 vccd1 vccd1 _05461_
+ sky130_fd_sc_hd__o221a_1
X_15015_ control.body\[987\] net167 _01553_ control.body\[979\] vssd1 vssd1 vccd1
+ vccd1 _00349_ sky130_fd_sc_hd__a22o_1
X_12227_ _04274_ _07196_ vssd1 vssd1 vccd1 vccd1 _07197_ sky130_fd_sc_hd__nor2_1
XANTENNA__11613__S0 net1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10135__A net1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18302__A track.nextHighScore\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19823_ clknet_leaf_89_clk _00767_ net1411 vssd1 vssd1 vccd1 vccd1 ag2.body\[573\]
+ sky130_fd_sc_hd__dfrtp_4
X_12158_ img_gen.tracker.frame\[456\] net614 net540 img_gen.tracker.frame\[462\] _07129_
+ vssd1 vssd1 vccd1 vccd1 _07130_ sky130_fd_sc_hd__o221a_1
XANTENNA__13446__A net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11109_ net1137 control.body\[1100\] vssd1 vssd1 vccd1 vccd1 _06082_ sky130_fd_sc_hd__nand2b_1
X_19754_ clknet_leaf_127_clk _00698_ net1326 vssd1 vssd1 vccd1 vccd1 control.body\[632\]
+ sky130_fd_sc_hd__dfrtp_1
X_16966_ ag2.body\[410\] net725 net709 ag2.body\[412\] vssd1 vssd1 vccd1 vccd1 _02645_
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_75_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12089_ img_gen.tracker.frame\[288\] net630 net557 img_gen.tracker.frame\[294\] vssd1
+ vssd1 vccd1 vccd1 _07061_ sky130_fd_sc_hd__a22o_1
X_18705_ clknet_leaf_10_clk img_gen.tracker.next_frame\[143\] net1275 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[143\] sky130_fd_sc_hd__dfrtp_1
X_15917_ ag2.body\[190\] net131 _01652_ ag2.body\[182\] vssd1 vssd1 vccd1 vccd1 _01152_
+ sky130_fd_sc_hd__a22o_1
X_19685_ clknet_leaf_136_clk _00629_ net1384 vssd1 vssd1 vccd1 vccd1 control.body\[707\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14829__X _01500_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16897_ ag2.body\[208\] net739 net719 ag2.body\[211\] _02575_ vssd1 vssd1 vccd1 vccd1
+ _02576_ sky130_fd_sc_hd__o221a_1
XANTENNA__16757__A net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17421__A2 net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18636_ clknet_leaf_131_clk img_gen.tracker.next_frame\[74\] net1295 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[74\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__09930__Y _04903_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15848_ ag2.body\[240\] net173 _01645_ ag2.body\[232\] vssd1 vssd1 vccd1 vccd1 _01090_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_103_3450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19510__CLK clknet_leaf_113_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_103_3461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_3472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18567_ clknet_leaf_14_clk img_gen.tracker.next_frame\[5\] net1278 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[5\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__14277__A net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15779_ ag2.body\[306\] net208 _01638_ ag2.body\[298\] vssd1 vssd1 vccd1 vccd1 _01028_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_75_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19836__RESET_B net1414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11253__X _06226_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17518_ ag2.body\[485\] net947 vssd1 vssd1 vccd1 vccd1 _03197_ sky130_fd_sc_hd__xor2_1
XFILLER_0_86_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13994__B2 ag2.body\[122\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18498_ net1515 net1509 vssd1 vssd1 vccd1 vccd1 _00029_ sky130_fd_sc_hd__or2_1
XFILLER_0_74_446 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15196__B1 _01573_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17449_ ag2.body\[378\] net724 net931 _04138_ _03121_ vssd1 vssd1 vccd1 vccd1 _03128_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_28_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20460_ clknet_leaf_30_clk _01347_ net1357 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[96\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_83_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_116_3855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_3866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11757__B1 net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkload57_A clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19119_ clknet_leaf_141_clk img_gen.tracker.next_frame\[557\] net1295 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[557\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10024__A3 _04978_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20391_ clknet_leaf_40_clk _01278_ net1374 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[27\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__16696__B1 net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_12_Right_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14171__A1 net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14171__B2 net1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16431__S net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10045__A net1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1027_A net1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09834__A net1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_2483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout487_A net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_2494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10699__B net1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09705_ _04662_ _04674_ _04676_ _04677_ vssd1 vssd1 vccd1 vccd1 _04678_ sky130_fd_sc_hd__or4_1
XFILLER_0_4_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout654_A _04394_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_94_clk clknet_4_11__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_94_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_138_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09636_ net1108 control.body\[1021\] vssd1 vssd1 vccd1 vccd1 _04609_ sky130_fd_sc_hd__xnor2_1
XANTENNA__19190__CLK clknet_leaf_53_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_21_Right_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_84_2877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_1499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_84_2888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18758__CLK clknet_leaf_15_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09567_ _04538_ _04539_ vssd1 vssd1 vccd1 vccd1 _04540_ sky130_fd_sc_hd__nor2_1
XANTENNA__14187__A net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout821_A net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_2899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16954__X _02633_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1184_X net1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout919_A net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13985__A1 ag2.body\[122\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_402 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_2298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09498_ net911 net919 net915 vssd1 vssd1 vccd1 vccd1 _04471_ sky130_fd_sc_hd__or3_4
XFILLER_0_110_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18373__B1 net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11996__B1 net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11323__B net1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10865__D _05837_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1351_X net1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15726__A2 net200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16606__S net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout707_X net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1449_X net1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11460_ _06429_ _06430_ _06431_ _06432_ _06428_ vssd1 vssd1 vccd1 vccd1 _06433_ sky130_fd_sc_hd__a221o_1
XFILLER_0_110_1288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_3_5_0_clk_X clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10411_ net1135 control.body\[1076\] vssd1 vssd1 vccd1 vccd1 _05384_ sky130_fd_sc_hd__xor2_1
XFILLER_0_46_1404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09728__B net1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11391_ net1120 control.body\[644\] vssd1 vssd1 vccd1 vccd1 _06364_ sky130_fd_sc_hd__xor2_1
X_20589_ net1521 vssd1 vssd1 vccd1 vccd1 gpio_oeb[1] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_30_Right_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13130_ img_gen.tracker.frame\[331\] net663 vssd1 vssd1 vccd1 vccd1 _07757_ sky130_fd_sc_hd__and2_1
XFILLER_0_33_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20064__RESET_B net1502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10342_ ag2.body\[521\] net780 net745 ag2.body\[527\] vssd1 vssd1 vccd1 vccd1 _05315_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_123_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14162__A1 net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13061_ net246 _07723_ _07724_ net2042 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[294\]
+ sky130_fd_sc_hd__a22o_1
X_10273_ ag2.body\[141\] net1113 vssd1 vssd1 vccd1 vccd1 _05246_ sky130_fd_sc_hd__xor2_1
XANTENNA__14162__B2 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18122__A net46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14650__A net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout90_X net90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16439__B1 net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12012_ net388 _06983_ vssd1 vssd1 vccd1 vccd1 _06984_ sky130_fd_sc_hd__or2_1
Xfanout1402 net1403 vssd1 vssd1 vccd1 vccd1 net1402 sky130_fd_sc_hd__clkbuf_4
Xfanout1413 net1414 vssd1 vssd1 vccd1 vccd1 net1413 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10723__A1 _05686_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_4151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11920__B1 net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1424 net1430 vssd1 vssd1 vccd1 vccd1 net1424 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10723__B2 _05671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_4162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16820_ _04012_ net876 net706 ag2.body\[85\] _02496_ vssd1 vssd1 vccd1 vccd1 _02499_
+ sky130_fd_sc_hd__o221a_1
XANTENNA__15111__B1 _01554_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1435 net1453 vssd1 vssd1 vccd1 vccd1 net1435 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_54_1980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09463__B net1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17651__A2 net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1446 net1448 vssd1 vssd1 vccd1 vccd1 net1446 sky130_fd_sc_hd__clkbuf_4
Xfanout1457 net1458 vssd1 vssd1 vccd1 vccd1 net1457 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_50_1833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1468 net1478 vssd1 vssd1 vccd1 vccd1 net1468 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_22_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_50_1844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout470 _06648_ vssd1 vssd1 vccd1 vccd1 net470 sky130_fd_sc_hd__buf_2
Xfanout481 net483 vssd1 vssd1 vccd1 vccd1 net481 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_35_1390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_4037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1479 net1480 vssd1 vssd1 vccd1 vccd1 net1479 sky130_fd_sc_hd__clkbuf_4
X_16751_ _02428_ _02429_ vssd1 vssd1 vccd1 vccd1 _02430_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_122_4048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout492 _01736_ vssd1 vssd1 vccd1 vccd1 net492 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_122_4059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13963_ ag2.body\[103\] net189 _08156_ ag2.body\[95\] vssd1 vssd1 vccd1 vccd1 _00184_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_31_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10402__B _04758_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_85_clk clknet_4_12__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_85_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_31_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15702_ ag2.body\[383\] net137 _01628_ ag2.body\[375\] vssd1 vssd1 vccd1 vccd1 _00961_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_134_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_1506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19470_ clknet_leaf_110_clk net2389 net1418 vssd1 vssd1 vccd1 vccd1 control.body\[924\]
+ sky130_fd_sc_hd__dfrtp_1
X_12914_ net244 _07654_ _07655_ net1808 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[216\]
+ sky130_fd_sc_hd__a22o_1
X_16682_ _02212_ _02333_ _02341_ _02360_ _02243_ vssd1 vssd1 vccd1 vccd1 _02361_ sky130_fd_sc_hd__o311a_1
X_13894_ ag2.body\[41\] net118 _08149_ ag2.body\[33\] vssd1 vssd1 vccd1 vccd1 _00122_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__09511__D_N _04472_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18421_ _03910_ _03889_ _08024_ net2058 vssd1 vssd1 vccd1 vccd1 _01397_ sky130_fd_sc_hd__o2bb2a_1
X_15633_ ag2.body\[432\] net125 _01622_ ag2.body\[424\] vssd1 vssd1 vccd1 vccd1 _00898_
+ sky130_fd_sc_hd__a22o_1
X_12845_ net286 _07622_ _07623_ net1781 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[179\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_57_1599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1170 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18352_ _04646_ _08032_ vssd1 vssd1 vccd1 vccd1 _03848_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_48_1773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15564_ ag2.body\[499\] net185 _01614_ ag2.body\[491\] vssd1 vssd1 vccd1 vccd1 _00837_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_48_1784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12776_ net225 _07590_ vssd1 vssd1 vccd1 vccd1 _07591_ sky130_fd_sc_hd__nor2_1
XANTENNA__19247__RESET_B net1482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11987__B1 net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17303_ ag2.body\[345\] net734 net934 _04125_ _02972_ vssd1 vssd1 vccd1 vccd1 _02982_
+ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_29_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14515_ net993 ag2.body\[313\] vssd1 vssd1 vccd1 vccd1 _08676_ sky130_fd_sc_hd__xor2_1
XFILLER_0_72_906 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11727_ img_gen.tracker.frame\[197\] net607 net552 img_gen.tracker.frame\[200\] _06698_
+ vssd1 vssd1 vccd1 vccd1 _06699_ sky130_fd_sc_hd__o221a_1
X_18283_ net517 _03780_ vssd1 vssd1 vccd1 vccd1 _01389_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_44_1659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15495_ ag2.body\[566\] net110 _01606_ ag2.body\[558\] vssd1 vssd1 vccd1 vccd1 _00776_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__16516__S net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17234_ ag2.body\[442\] net724 net930 _04159_ vssd1 vssd1 vccd1 vccd1 _02913_ sky130_fd_sc_hd__a22o_1
XFILLER_0_86_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14925__B1 _01543_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11658_ net1071 net1045 vssd1 vssd1 vccd1 vccd1 _06631_ sky130_fd_sc_hd__and2_1
X_14446_ net983 ag2.body\[226\] vssd1 vssd1 vccd1 vccd1 _08607_ sky130_fd_sc_hd__xor2_1
XFILLER_0_9_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10609_ net1204 control.body\[985\] vssd1 vssd1 vccd1 vccd1 _05582_ sky130_fd_sc_hd__xor2_1
X_14377_ net1029 ag2.body\[421\] vssd1 vssd1 vccd1 vccd1 _08538_ sky130_fd_sc_hd__xnor2_1
XANTENNA__16127__C1 net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17165_ _04218_ net868 net722 ag2.body\[594\] _02841_ vssd1 vssd1 vccd1 vccd1 _02844_
+ sky130_fd_sc_hd__a221o_1
X_11589_ _06527_ _06561_ vssd1 vssd1 vccd1 vccd1 _06562_ sky130_fd_sc_hd__xnor2_1
XANTENNA__12345__A _07306_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_94_3184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_94_3195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold907 _00278_ vssd1 vssd1 vccd1 vccd1 net2469 sky130_fd_sc_hd__dlygate4sd3_1
X_16116_ obsg2.obstacleArray\[92\] obsg2.obstacleArray\[93\] net424 vssd1 vssd1 vccd1
+ vccd1 _01795_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13328_ net664 _07844_ vssd1 vssd1 vccd1 vccd1 _07845_ sky130_fd_sc_hd__nor2_1
Xhold918 control.body\[637\] vssd1 vssd1 vccd1 vccd1 net2480 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17096_ ag2.body\[296\] net886 vssd1 vssd1 vccd1 vccd1 _02775_ sky130_fd_sc_hd__or2_1
Xhold929 control.body\[624\] vssd1 vssd1 vccd1 vccd1 net2491 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_90_3059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19063__CLK clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18419__A1 _04646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16047_ net502 _01716_ _01717_ vssd1 vssd1 vccd1 vccd1 _01726_ sky130_fd_sc_hd__and3_1
X_13259_ net670 _07817_ vssd1 vssd1 vccd1 vccd1 _07818_ sky130_fd_sc_hd__nor2_1
XANTENNA__18032__A net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12164__B1 net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09654__A net1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11911__B1 net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09580__A1 _04471_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19806_ clknet_leaf_125_clk _00750_ net1410 vssd1 vssd1 vccd1 vccd1 ag2.body\[588\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__17642__A2 net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17998_ net484 net345 _03561_ vssd1 vssd1 vccd1 vccd1 _03613_ sky130_fd_sc_hd__and3_1
XFILLER_0_97_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16850__B1 net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_3512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19737_ clknet_leaf_132_clk _00681_ net1304 vssd1 vssd1 vccd1 vccd1 control.body\[663\]
+ sky130_fd_sc_hd__dfrtp_1
X_16949_ ag2.body\[384\] net884 vssd1 vssd1 vccd1 vccd1 _02628_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_105_3523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12011__S0 net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_92_clk_A clknet_4_9__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11408__B net1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_3534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14861__C1 _01531_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_76_clk clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_76_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_79_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18900__CLK clknet_leaf_144_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__20190__CLK clknet_leaf_88_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09660__Y _04633_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19668_ clknet_leaf_118_clk _00612_ net1390 vssd1 vssd1 vccd1 vccd1 control.body\[722\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_101_3409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09883__A2 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09421_ ag2.goodColl _04398_ net516 vssd1 vssd1 vccd1 vccd1 _04400_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_17_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18619_ clknet_leaf_144_clk img_gen.tracker.next_frame\[57\] net1241 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[57\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_133_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19599_ clknet_leaf_118_clk _00543_ net1390 vssd1 vssd1 vccd1 vccd1 control.body\[797\]
+ sky130_fd_sc_hd__dfrtp_1
X_09352_ sound_gen.osc1.stayCount\[8\] sound_gen.osc1.stayCount\[7\] _04345_ vssd1
+ vssd1 vccd1 vccd1 _04354_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_118_3917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11978__B1 net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16934__B net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11143__B net1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_118_3928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_60_2140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09283_ _04303_ _04305_ vssd1 vssd1 vccd1 vccd1 _04306_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_60_2151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16366__C1 net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14735__A net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_2162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout235_A net236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20512_ clknet_leaf_113_clk track.nextHighScore\[2\] net1402 vssd1 vssd1 vccd1 vccd1
+ track.highScore\[2\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__09829__A net1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1648 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_30_clk_A clknet_4_4__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14392__A1 net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19406__CLK clknet_leaf_103_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20443_ clknet_leaf_25_clk _01330_ net1343 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[79\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__14392__B2 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout402_A net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10327__X _05300_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1144_A net1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_2670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_2681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20374_ clknet_leaf_23_clk _01261_ net1358 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[10\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_28_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_58_2080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20595__1527 vssd1 vssd1 vccd1 vccd1 _20595__1527/HI net1527 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_73_2545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_2091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload80 clknet_leaf_89_clk vssd1 vssd1 vccd1 vccd1 clkload80/Y sky130_fd_sc_hd__clkinv_8
XANTENNA_clkbuf_leaf_45_clk_A clknet_4_7__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_2556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15341__B1 _01590_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload91 clknet_leaf_109_clk vssd1 vssd1 vccd1 vccd1 clkload91/Y sky130_fd_sc_hd__bufinv_16
XFILLER_0_28_1178 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16161__S net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1311_A net1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18552__RESET_B net1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12155__B1 net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1409_A net1415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09564__A net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout392_X net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout771_A _04230_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11902__B1 net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout869_A obsg2.randCord\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10062__X _05035_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08998_ ag2.body\[97\] vssd1 vssd1 vccd1 vccd1 _04023_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_3_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12458__A1 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11318__B net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_86_2939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_67_clk clknet_4_13__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_67_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__14852__C1 _01522_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16397__A net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout657_X net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10222__B net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_302 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_103_clk_A clknet_4_10__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10960_ ag2.body\[169\] net1209 vssd1 vssd1 vccd1 vccd1 _05933_ sky130_fd_sc_hd__xor2_1
XFILLER_0_138_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09619_ net1075 control.body\[806\] vssd1 vssd1 vccd1 vccd1 _04592_ sky130_fd_sc_hd__xor2_1
XANTENNA__17005__B net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout824_X net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10891_ net1173 control.body\[650\] vssd1 vssd1 vccd1 vccd1 _05864_ sky130_fd_sc_hd__xor2_1
XANTENNA__11681__A2 net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15947__A2 net195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17720__S net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12630_ img_gen.tracker.frame\[71\] net644 _07516_ vssd1 vssd1 vccd1 vccd1 _07517_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_17_1572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16844__B net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_118_clk_A clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_134_4420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11053__B net1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12561_ net334 _07479_ vssd1 vssd1 vccd1 vccd1 _07480_ sky130_fd_sc_hd__nand2_2
XFILLER_0_93_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_1504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_1496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16336__S net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18117__A net44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11512_ _06482_ _06483_ vssd1 vssd1 vccd1 vccd1 _06485_ sky130_fd_sc_hd__nand2_8
X_14300_ net1021 ag2.body\[222\] vssd1 vssd1 vccd1 vccd1 _08461_ sky130_fd_sc_hd__xor2_1
XFILLER_0_19_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_980 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15280_ net2257 net89 _01583_ control.body\[750\] vssd1 vssd1 vccd1 vccd1 _00584_
+ sky130_fd_sc_hd__a22o_1
X_12492_ net678 _07440_ vssd1 vssd1 vccd1 vccd1 _07441_ sky130_fd_sc_hd__nor2_1
XANTENNA__11988__B net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_1559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14231_ net824 ag2.body\[482\] ag2.body\[484\] net813 vssd1 vssd1 vccd1 vccd1 _08392_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__14383__A1 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11443_ net1229 control.body\[952\] vssd1 vssd1 vccd1 vccd1 _06416_ sky130_fd_sc_hd__nand2_1
XANTENNA__14383__B2 net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09458__B _04421_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11197__A1 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11197__B2 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14162_ net832 ag2.body\[617\] ag2.body\[621\] net806 _08322_ vssd1 vssd1 vccd1 vccd1
+ _08323_ sky130_fd_sc_hd__o221a_1
XFILLER_0_132_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11374_ _04170_ net1104 net749 ag2.body\[478\] _06346_ vssd1 vssd1 vccd1 vccd1 _06347_
+ sky130_fd_sc_hd__a221o_1
XANTENNA__20063__CLK clknet_leaf_73_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13113_ net1905 net652 _07748_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[322\]
+ sky130_fd_sc_hd__and3_1
X_10325_ ag2.body\[613\] net1097 vssd1 vssd1 vccd1 vccd1 _05298_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_128_4213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16071__S net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14093_ net820 ag2.body\[283\] ag2.body\[284\] net816 _08253_ vssd1 vssd1 vccd1 vccd1
+ _08254_ sky130_fd_sc_hd__a221o_1
X_18970_ clknet_leaf_7_clk img_gen.tracker.next_frame\[408\] net1266 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[408\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_128_4224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_128_4235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17921_ net48 net296 _03554_ vssd1 vssd1 vccd1 vccd1 _03555_ sky130_fd_sc_hd__and3_1
X_13044_ net2109 net651 _07716_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[285\]
+ sky130_fd_sc_hd__and3_1
X_10256_ net1201 control.body\[785\] vssd1 vssd1 vccd1 vccd1 _05229_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_37_1452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1210 net1212 vssd1 vssd1 vccd1 vccd1 net1210 sky130_fd_sc_hd__buf_4
XANTENNA__17085__B1 net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11068__X _06041_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09562__A1 _04512_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1221 ag2.y\[0\] vssd1 vssd1 vccd1 vccd1 net1221 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_33_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17852_ img_gen.updater.commands.rR1.rainbowRNG\[0\] net248 vssd1 vssd1 vccd1 vccd1
+ _03508_ sky130_fd_sc_hd__nor2_1
XANTENNA__09562__B2 _04534_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1232 net1238 vssd1 vssd1 vccd1 vccd1 net1232 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_33_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10187_ _05152_ _05157_ _05158_ _05159_ vssd1 vssd1 vccd1 vccd1 _05160_ sky130_fd_sc_hd__or4_2
XANTENNA__10413__A net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1243 net1333 vssd1 vssd1 vccd1 vccd1 net1243 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_98_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1254 net1263 vssd1 vssd1 vccd1 vccd1 net1254 sky130_fd_sc_hd__clkbuf_2
X_16803_ ag2.body\[64\] net888 vssd1 vssd1 vccd1 vccd1 _02482_ sky130_fd_sc_hd__xor2_1
Xfanout1265 net1267 vssd1 vssd1 vccd1 vccd1 net1265 sky130_fd_sc_hd__clkbuf_4
Xfanout1276 net1280 vssd1 vssd1 vccd1 vccd1 net1276 sky130_fd_sc_hd__clkbuf_4
X_17783_ net807 net800 net792 vssd1 vssd1 vccd1 vccd1 _03461_ sky130_fd_sc_hd__or3_1
Xfanout1287 net1333 vssd1 vssd1 vccd1 vccd1 net1287 sky130_fd_sc_hd__buf_2
Xclkbuf_leaf_58_clk clknet_4_13__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_58_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_89_814 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14995_ control.body\[1001\] net153 _01551_ control.body\[993\] vssd1 vssd1 vccd1
+ vccd1 _00331_ sky130_fd_sc_hd__a22o_1
Xfanout1298 net1310 vssd1 vssd1 vccd1 vccd1 net1298 sky130_fd_sc_hd__clkbuf_4
X_19522_ clknet_leaf_120_clk net2277 net1401 vssd1 vssd1 vccd1 vccd1 control.body\[864\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_92_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16734_ obsg2.obstacleArray\[100\] net490 net486 obsg2.obstacleArray\[102\] _02412_
+ vssd1 vssd1 vccd1 vccd1 _02413_ sky130_fd_sc_hd__a221o_1
XFILLER_0_57_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13946_ _04698_ net67 vssd1 vssd1 vccd1 vccd1 _08155_ sky130_fd_sc_hd__and2_2
XFILLER_0_72_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19453_ clknet_leaf_111_clk _00397_ net1427 vssd1 vssd1 vccd1 vccd1 control.body\[939\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__15399__B1 _01581_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16665_ obsg2.obstacleArray\[23\] net451 net393 _02343_ vssd1 vssd1 vccd1 vccd1 _02344_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_9_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15938__A2 net196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13877_ ag2.body\[26\] net115 _08147_ ag2.body\[18\] vssd1 vssd1 vccd1 vccd1 _00107_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11672__A2 net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18404_ _04638_ _03832_ _03893_ _03828_ vssd1 vssd1 vccd1 vccd1 _03894_ sky130_fd_sc_hd__a211o_1
X_15616_ ag2.body\[449\] net123 _01613_ ag2.body\[441\] vssd1 vssd1 vccd1 vccd1 _00883_
+ sky130_fd_sc_hd__a22o_1
X_12828_ _06672_ _07522_ vssd1 vssd1 vccd1 vccd1 _07615_ sky130_fd_sc_hd__or2_1
X_19384_ clknet_leaf_112_clk _00328_ net1426 vssd1 vssd1 vccd1 vccd1 control.body\[1014\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16596_ obsg2.obstacleArray\[79\] net449 net390 _02274_ vssd1 vssd1 vccd1 vccd1 _02275_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_118_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18335_ _08139_ _03830_ vssd1 vssd1 vccd1 vccd1 _03831_ sky130_fd_sc_hd__and2_1
X_15547_ ag2.body\[517\] net162 _01580_ ag2.body\[509\] vssd1 vssd1 vccd1 vccd1 _00823_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__16246__S net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12759_ net258 _07582_ _07583_ net1684 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[133\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_122_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_96_3246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09649__A net1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_96_3257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18266_ net319 _03555_ obsg2.obstacleArray\[130\] vssd1 vssd1 vccd1 vccd1 _03772_
+ sky130_fd_sc_hd__a21oi_1
X_15478_ ag2.body\[583\] net108 _01604_ ag2.body\[575\] vssd1 vssd1 vccd1 vccd1 _00761_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_112_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_175 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17217_ _02890_ _02892_ _02894_ _02895_ vssd1 vssd1 vccd1 vccd1 _02896_ sky130_fd_sc_hd__or4_1
X_14429_ net997 ag2.body\[552\] vssd1 vssd1 vccd1 vccd1 _08590_ sky130_fd_sc_hd__xor2_1
X_18197_ net519 _03737_ vssd1 vssd1 vccd1 vccd1 _01346_ sky130_fd_sc_hd__nor2_1
XFILLER_0_126_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_1443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold704 _00632_ vssd1 vssd1 vccd1 vccd1 net2266 sky130_fd_sc_hd__dlygate4sd3_1
X_17148_ ag2.body\[608\] net879 vssd1 vssd1 vccd1 vccd1 _02827_ sky130_fd_sc_hd__xor2_1
Xhold715 _00466_ vssd1 vssd1 vccd1 vccd1 net2277 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1611 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold726 _00552_ vssd1 vssd1 vccd1 vccd1 net2288 sky130_fd_sc_hd__dlygate4sd3_1
Xhold737 _00280_ vssd1 vssd1 vccd1 vccd1 net2299 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10935__B2 _04646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14126__A1 net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14126__B2 net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09970_ _04862_ _04942_ vssd1 vssd1 vccd1 vccd1 _04943_ sky130_fd_sc_hd__or2_1
Xhold748 _00693_ vssd1 vssd1 vccd1 vccd1 net2310 sky130_fd_sc_hd__dlygate4sd3_1
X_17079_ ag2.body\[196\] net962 vssd1 vssd1 vccd1 vccd1 _02758_ sky130_fd_sc_hd__nand2_1
Xhold759 control.body\[913\] vssd1 vssd1 vccd1 vccd1 net2321 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__20556__CLK clknet_leaf_105_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20090_ clknet_leaf_78_clk _01034_ net1490 vssd1 vssd1 vccd1 vccd1 ag2.body\[296\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_42_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11419__A net1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13337__C _07813_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11360__B2 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11138__B _06110_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout185_A net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11112__A1 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11112__B2 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17878__A_N _04903_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_2803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout352_A net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16587__C1 net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_62_2202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1604 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_62_2213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09404_ sound_gen.osc1.stayCount\[0\] _04305_ net2399 vssd1 vssd1 vccd1 vccd1 _04386_
+ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout1094_A net1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_2224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16664__B net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09335_ sound_gen.at_max sound_gen.dac1.dacCount\[0\] net1888 vssd1 vssd1 vccd1 vccd1
+ _04341_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12612__A1 net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10993__A ag2.body\[340\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout617_A net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14465__A net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17000__B1 net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout238_X net238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1359_A net1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_79_2721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09266_ sound_gen.osc1.stayCount\[6\] _04288_ sound_gen.osc1.stayCount\[7\] vssd1
+ vssd1 vccd1 vccd1 _04289_ sky130_fd_sc_hd__o21a_1
XANTENNA__09559__A net1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_2732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13800__C net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_2743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15995__S net223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_2607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09197_ ag2.body\[616\] vssd1 vssd1 vccd1 vccd1 _04222_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_75_2618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1147_X net1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_2017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20426_ clknet_leaf_38_clk _01313_ net1353 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[62\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__17839__C1 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16106__A2 _01780_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_2028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10926__A1 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_2039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout986_A ag2.randCord\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14912__B net51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10926__B2 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14117__A1 net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18946__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14117__B2 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20357_ clknet_leaf_18_clk _01248_ net1323 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleCount\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_101_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10110_ net1179 control.body\[938\] vssd1 vssd1 vccd1 vccd1 _05083_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout98_A net100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12679__A1 net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11090_ _04198_ net1084 _06060_ _06061_ _06062_ vssd1 vssd1 vccd1 vccd1 _06063_ sky130_fd_sc_hd__a2111o_1
X_20288_ clknet_leaf_35_clk control.divider.next_count\[9\] net1350 vssd1 vssd1 vccd1
+ vccd1 control.divider.count\[9\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_101_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_8_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout774_X net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09544__A1 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17715__S net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10041_ net1058 control.body\[903\] vssd1 vssd1 vccd1 vccd1 _05014_ sky130_fd_sc_hd__xor2_1
XANTENNA__11329__A net1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17606__A2 net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11887__C1 net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold20 control.detect2.Q\[0\] vssd1 vssd1 vccd1 vccd1 net1582 sky130_fd_sc_hd__dlygate4sd3_1
Xhold31 img_gen.tracker.frame\[101\] vssd1 vssd1 vccd1 vccd1 net1593 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__16814__B1 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold42 img_gen.tracker.frame\[236\] vssd1 vssd1 vccd1 vccd1 net1604 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11048__B net1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold53 img_gen.tracker.frame\[413\] vssd1 vssd1 vccd1 vccd1 net1615 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout941_X net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16871__A2_N net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold64 img_gen.tracker.frame\[524\] vssd1 vssd1 vccd1 vccd1 net1626 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__19592__RESET_B net1404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11763__S net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold75 img_gen.tracker.frame\[474\] vssd1 vssd1 vccd1 vccd1 net1637 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_118_1515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13800_ _06632_ _07178_ net465 vssd1 vssd1 vccd1 vccd1 _08104_ sky130_fd_sc_hd__and3_1
Xhold86 img_gen.tracker.frame\[466\] vssd1 vssd1 vccd1 vccd1 net1648 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09741__B net1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_622 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold97 img_gen.tracker.frame\[189\] vssd1 vssd1 vccd1 vccd1 net1659 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_19_1601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11992_ _06959_ _06961_ _06963_ net560 vssd1 vssd1 vccd1 vccd1 _06964_ sky130_fd_sc_hd__a22o_1
X_14780_ net1020 ag2.body\[278\] vssd1 vssd1 vccd1 vccd1 _01451_ sky130_fd_sc_hd__nand2_1
XFILLER_0_19_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout53_X net53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10943_ ag2.body\[299\] _04230_ net752 ag2.body\[302\] _05912_ vssd1 vssd1 vccd1
+ vccd1 _05916_ sky130_fd_sc_hd__a221o_1
X_13731_ _04391_ _07210_ _07244_ _07259_ vssd1 vssd1 vccd1 vccd1 _08055_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__09460__C net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_919 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16450_ net399 _02128_ vssd1 vssd1 vccd1 vccd1 _02129_ sky130_fd_sc_hd__or2_1
XFILLER_0_116_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13662_ net998 net835 _08014_ _08015_ vssd1 vssd1 vccd1 vccd1 _08016_ sky130_fd_sc_hd__o22a_1
XFILLER_0_42_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_3_0_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_3_0_0_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_45_1710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10874_ ag2.body\[531\] net1158 vssd1 vssd1 vccd1 vccd1 _05847_ sky130_fd_sc_hd__nand2_1
XFILLER_0_112_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16574__B net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15401_ net2583 net80 _01581_ net2289 vssd1 vssd1 vccd1 vccd1 _00692_ sky130_fd_sc_hd__a22o_1
XFILLER_0_112_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12613_ net609 _06639_ net438 net569 vssd1 vssd1 vccd1 vccd1 _07508_ sky130_fd_sc_hd__and4_2
XTAP_TAPCELL_ROW_26_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13593_ _03960_ control.divider.count\[12\] _07953_ control.divider.count\[13\] control.divider.count\[11\]
+ vssd1 vssd1 vccd1 vccd1 _07968_ sky130_fd_sc_hd__a221o_1
X_16381_ _01900_ _02058_ vssd1 vssd1 vccd1 vccd1 _02060_ sky130_fd_sc_hd__nand2_1
XANTENNA__14375__A net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18120_ net526 _03695_ vssd1 vssd1 vccd1 vccd1 _01311_ sky130_fd_sc_hd__and2_1
XFILLER_0_66_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15332_ net2247 net74 _01587_ net2307 vssd1 vssd1 vccd1 vccd1 _00630_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_22_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12544_ net225 _07469_ vssd1 vssd1 vccd1 vccd1 _07470_ sky130_fd_sc_hd__nor2_1
XFILLER_0_108_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09480__B1 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19721__CLK clknet_leaf_132_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10090__A1 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12607__B net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14356__A1 net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18051_ obsg2.obstacleArray\[36\] _03650_ net522 vssd1 vssd1 vccd1 vccd1 _01287_
+ sky130_fd_sc_hd__o21a_1
XANTENNA__10090__B2 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14356__B2 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12475_ _06821_ net315 vssd1 vssd1 vccd1 vccd1 _07430_ sky130_fd_sc_hd__nor2_1
X_15263_ _04573_ net52 vssd1 vssd1 vccd1 vccd1 _01581_ sky130_fd_sc_hd__nor2_4
XFILLER_0_48_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10408__A net1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1610 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_3110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17002_ _04037_ net865 net702 ag2.body\[142\] vssd1 vssd1 vccd1 vccd1 _02681_ sky130_fd_sc_hd__o22a_1
X_14214_ net801 ag2.body\[414\] ag2.body\[415\] net793 _08374_ vssd1 vssd1 vccd1 vccd1
+ _08375_ sky130_fd_sc_hd__a221o_1
X_11426_ _04556_ _04982_ _04472_ vssd1 vssd1 vccd1 vccd1 _06399_ sky130_fd_sc_hd__o21ba_1
XANTENNA_6 _03442_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15194_ control.body\[826\] net94 _01573_ net2551 vssd1 vssd1 vccd1 vccd1 _00508_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_39_1503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_1514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_39_1525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14145_ net996 ag2.body\[592\] vssd1 vssd1 vccd1 vccd1 _08306_ sky130_fd_sc_hd__xnor2_1
X_11357_ net1201 control.body\[809\] vssd1 vssd1 vccd1 vccd1 _06330_ sky130_fd_sc_hd__nand2_1
XFILLER_0_22_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12119__B1 net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18013__C net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10308_ net1072 control.body\[702\] vssd1 vssd1 vccd1 vccd1 _05281_ sky130_fd_sc_hd__nand2_1
X_18953_ clknet_leaf_5_clk img_gen.tracker.next_frame\[391\] net1276 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[391\] sky130_fd_sc_hd__dfrtp_1
X_14076_ net813 ag2.body\[564\] ag2.body\[566\] net799 vssd1 vssd1 vccd1 vccd1 _08237_
+ sky130_fd_sc_hd__o22a_1
X_11288_ net1136 control.body\[1108\] vssd1 vssd1 vccd1 vccd1 _06261_ sky130_fd_sc_hd__nand2_1
XANTENNA__17058__B1 net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17904_ net381 _02054_ vssd1 vssd1 vccd1 vccd1 _03539_ sky130_fd_sc_hd__nor2_2
X_13027_ net673 _07708_ vssd1 vssd1 vccd1 vccd1 _07709_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_89_3050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10239_ net903 _04493_ _04417_ vssd1 vssd1 vccd1 vccd1 _05212_ sky130_fd_sc_hd__a21oi_4
XANTENNA__10143__A net1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18884_ clknet_leaf_12_clk img_gen.tracker.next_frame\[322\] net1281 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[322\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__10145__A2 _04759_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1040 net1042 vssd1 vssd1 vccd1 vccd1 net1040 sky130_fd_sc_hd__clkbuf_8
XANTENNA__16805__B1 net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1248 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1051 net1052 vssd1 vssd1 vccd1 vccd1 net1051 sky130_fd_sc_hd__clkbuf_4
X_17835_ net662 _03494_ vssd1 vssd1 vccd1 vccd1 _01227_ sky130_fd_sc_hd__and2_1
Xfanout1062 net1063 vssd1 vssd1 vccd1 vccd1 net1062 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_98_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1073 net1074 vssd1 vssd1 vccd1 vccd1 net1073 sky130_fd_sc_hd__buf_4
Xfanout1084 net1093 vssd1 vssd1 vccd1 vccd1 net1084 sky130_fd_sc_hd__buf_4
Xfanout1095 net1096 vssd1 vssd1 vccd1 vccd1 net1095 sky130_fd_sc_hd__clkbuf_4
X_17766_ _02662_ _03230_ _03443_ _03444_ vssd1 vssd1 vccd1 vccd1 _03445_ sky130_fd_sc_hd__and4b_1
XFILLER_0_83_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19262__RESET_B net1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14978_ control.body\[1017\] net153 _01550_ net2368 vssd1 vssd1 vccd1 vccd1 _00315_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_88_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16005__A_N net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1040 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19505_ clknet_leaf_113_clk _00449_ net1404 vssd1 vssd1 vccd1 vccd1 control.body\[895\]
+ sky130_fd_sc_hd__dfrtp_1
X_16717_ obsg2.obstacleArray\[120\] net491 net482 obsg2.obstacleArray\[121\] _02395_
+ vssd1 vssd1 vccd1 vccd1 _02396_ sky130_fd_sc_hd__a221o_1
X_13929_ ag2.body\[72\] net193 _08153_ ag2.body\[64\] vssd1 vssd1 vccd1 vccd1 _00153_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__19251__CLK clknet_leaf_75_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17697_ _03372_ _03373_ _03375_ vssd1 vssd1 vccd1 vccd1 _03376_ sky130_fd_sc_hd__or3_1
XANTENNA__16569__C1 net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17230__B1 net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20594__1526 vssd1 vssd1 vccd1 vccd1 _20594__1526/HI net1526 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_18_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19436_ clknet_leaf_108_clk _00380_ net1421 vssd1 vssd1 vccd1 vccd1 control.body\[954\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_130_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16648_ obsg2.obstacleArray\[0\] obsg2.obstacleArray\[1\] net446 vssd1 vssd1 vccd1
+ vccd1 _02327_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_18_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_3308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_3319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19367_ clknet_leaf_93_clk net2224 net1438 vssd1 vssd1 vccd1 vccd1 control.body\[1029\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13901__B net52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16579_ obsg2.obstacleArray\[115\] net449 net390 _02257_ vssd1 vssd1 vccd1 vccd1
+ _02258_ sky130_fd_sc_hd__o211a_1
X_09120_ ag2.body\[405\] vssd1 vssd1 vccd1 vccd1 _04145_ sky130_fd_sc_hd__inv_2
XFILLER_0_44_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18318_ net322 _03813_ _03793_ vssd1 vssd1 vccd1 vccd1 _03814_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_17_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19298_ clknet_leaf_100_clk _00242_ net1444 vssd1 vssd1 vccd1 vccd1 control.body\[1088\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12070__A2 net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09051_ ag2.body\[241\] vssd1 vssd1 vccd1 vccd1 _04076_ sky130_fd_sc_hd__inv_2
X_18249_ obsg2.obstacleArray\[121\] _03763_ net525 vssd1 vssd1 vccd1 vccd1 _01372_
+ sky130_fd_sc_hd__o21a_1
XPHY_EDGE_ROW_6_Right_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16704__S net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold501 img_gen.tracker.frame\[169\] vssd1 vssd1 vccd1 vccd1 net2063 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold512 img_gen.tracker.frame\[12\] vssd1 vssd1 vccd1 vccd1 net2074 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__17297__B1 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20211_ clknet_leaf_60_clk _01155_ net1466 vssd1 vssd1 vccd1 vccd1 ag2.body\[177\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__18204__B net40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold523 control.body\[1036\] vssd1 vssd1 vccd1 vccd1 net2085 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11848__S net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17883__X _03523_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold534 img_gen.tracker.frame\[214\] vssd1 vssd1 vccd1 vccd1 net2096 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout100_A net114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold545 img_gen.tracker.frame\[106\] vssd1 vssd1 vccd1 vccd1 net2107 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold556 sound_gen.dac1.dacCount\[5\] vssd1 vssd1 vccd1 vccd1 net2118 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12533__A net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold567 img_gen.tracker.frame\[558\] vssd1 vssd1 vccd1 vccd1 net2129 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__20523__Q control.body_update.curr_length\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold578 img_gen.tracker.frame\[63\] vssd1 vssd1 vccd1 vccd1 net2140 sky130_fd_sc_hd__dlygate4sd3_1
X_20142_ clknet_leaf_96_clk _01086_ net1451 vssd1 vssd1 vccd1 vccd1 ag2.body\[252\]
+ sky130_fd_sc_hd__dfrtp_2
Xhold589 _00418_ vssd1 vssd1 vccd1 vccd1 net2151 sky130_fd_sc_hd__dlygate4sd3_1
X_09953_ net783 control.body\[736\] _04923_ _04924_ _04925_ vssd1 vssd1 vccd1 vccd1
+ _04926_ sky130_fd_sc_hd__o2111ai_1
Xmax_cap297 _07835_ vssd1 vssd1 vccd1 vccd1 net297 sky130_fd_sc_hd__buf_1
XANTENNA__13858__B1 _08134_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17049__B1 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20073_ clknet_leaf_73_clk _01017_ net1501 vssd1 vssd1 vccd1 vccd1 ag2.body\[327\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__10053__A _04429_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09884_ ag2.body\[161\] net778 net763 ag2.body\[164\] _04856_ vssd1 vssd1 vccd1 vccd1
+ _04857_ sky130_fd_sc_hd__o221a_1
XANTENNA__18220__A _03662_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1107_A net1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_2400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_2411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1095 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13086__A1 net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12833__A1 net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17757__D1 net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout734_A net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1476_A net1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1097_X net1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10844__B1 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16575__A2 net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_1445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14586__A1 net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14586__B2 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout901_A control.body_update.curr_length\[5\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_48_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12708__A net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09318_ sound_gen.osc1.count\[1\] sound_gen.osc1.count\[0\] sound_gen.osc1.count\[2\]
+ vssd1 vssd1 vccd1 vccd1 _04333_ sky130_fd_sc_hd__a21o_1
XFILLER_0_88_1632 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12061__A2 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10590_ net1076 control.body\[830\] vssd1 vssd1 vccd1 vccd1 _05563_ sky130_fd_sc_hd__nand2_1
XFILLER_0_118_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16327__A2 net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09249_ img_gen.updater.commands.cmd_num\[2\] vssd1 vssd1 vccd1 vccd1 _04274_ sky130_fd_sc_hd__inv_2
XFILLER_0_90_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12260_ _07224_ _07229_ vssd1 vssd1 vccd1 vccd1 _07230_ sky130_fd_sc_hd__nand2_1
XANTENNA__13010__A1 net240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout891_X net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout989_X net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18114__B _03691_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11211_ net1201 control.body\[841\] vssd1 vssd1 vccd1 vccd1 _06184_ sky130_fd_sc_hd__xnor2_1
X_20409_ clknet_leaf_31_clk _01296_ net1338 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[45\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_47_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12191_ net1054 ag2.apple_cord\[7\] vssd1 vssd1 vccd1 vccd1 _07163_ sky130_fd_sc_hd__nand2_1
Xoutput10 net10 vssd1 vssd1 vccd1 vccd1 gpio_out[0] sky130_fd_sc_hd__buf_2
XANTENNA__11572__A1 net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput21 net21 vssd1 vssd1 vccd1 vccd1 gpio_out[1] sky130_fd_sc_hd__buf_2
XANTENNA__19124__CLK clknet_leaf_141_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput32 net32 vssd1 vssd1 vccd1 vccd1 gpio_out[7] sky130_fd_sc_hd__buf_2
X_11142_ ag2.body\[409\] net1209 vssd1 vssd1 vccd1 vccd1 _06115_ sky130_fd_sc_hd__xor2_1
XANTENNA__14510__A1 net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15950_ ag2.body\[155\] net199 _01656_ ag2.body\[147\] vssd1 vssd1 vccd1 vccd1 _01181_
+ sky130_fd_sc_hd__a22o_1
X_11073_ ag2.body\[363\] net772 net784 ag2.body\[360\] vssd1 vssd1 vccd1 vccd1 _06046_
+ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__14510__B2 net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10024_ _04967_ _04968_ _04978_ _04986_ _04996_ vssd1 vssd1 vccd1 vccd1 _04997_ sky130_fd_sc_hd__o32a_1
X_14901_ control.body\[1094\] net177 _01540_ net2323 vssd1 vssd1 vccd1 vccd1 _00248_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_95_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15881_ ag2.body\[222\] net192 _01648_ ag2.body\[214\] vssd1 vssd1 vccd1 vccd1 _01120_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11875__A2 net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13274__A net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17620_ _03295_ _03297_ _03298_ vssd1 vssd1 vccd1 vccd1 _03299_ sky130_fd_sc_hd__or3b_2
XFILLER_0_99_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14832_ _08594_ _08597_ _08602_ _08623_ vssd1 vssd1 vccd1 vccd1 _01503_ sky130_fd_sc_hd__o31a_1
X_17551_ _03223_ _03229_ vssd1 vssd1 vccd1 vccd1 _03230_ sky130_fd_sc_hd__or2_2
XFILLER_0_53_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14763_ _08915_ _08916_ _08918_ _08923_ vssd1 vssd1 vccd1 vccd1 _08924_ sky130_fd_sc_hd__or4b_4
XFILLER_0_114_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11975_ img_gen.tracker.frame\[574\] net588 net575 vssd1 vssd1 vccd1 vccd1 _06947_
+ sky130_fd_sc_hd__o21a_1
X_16502_ _02180_ _02057_ _02176_ vssd1 vssd1 vccd1 vccd1 _02181_ sky130_fd_sc_hd__or3b_1
XANTENNA__17212__B1 net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13714_ track.highScore\[3\] _04641_ net356 vssd1 vssd1 vccd1 vccd1 track.nextHighScore\[3\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17482_ ag2.body\[131\] net721 net694 ag2.body\[135\] vssd1 vssd1 vccd1 vccd1 _03161_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_19_1486 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10926_ net769 control.body\[1035\] control.body\[1036\] net761 _05898_ vssd1 vssd1
+ vccd1 vccd1 _05899_ sky130_fd_sc_hd__a221o_1
X_14694_ net978 ag2.body\[323\] vssd1 vssd1 vccd1 vccd1 _08855_ sky130_fd_sc_hd__xor2_1
X_19221_ clknet_leaf_85_clk _00165_ net1483 vssd1 vssd1 vccd1 vccd1 ag2.body\[84\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_116_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16433_ obsg2.obstacleArray\[79\] _02059_ net397 _02111_ vssd1 vssd1 vccd1 vccd1
+ _02112_ sky130_fd_sc_hd__o211a_1
X_13645_ _08003_ _08004_ vssd1 vssd1 vccd1 vccd1 control.divider.next_count\[15\]
+ sky130_fd_sc_hd__nor2_1
X_10857_ net1046 control.body\[695\] vssd1 vssd1 vccd1 vccd1 _05830_ sky130_fd_sc_hd__xor2_1
XANTENNA__13721__B net25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19152_ clknet_leaf_52_clk _00096_ net1367 vssd1 vssd1 vccd1 vccd1 ag2.body\[16\]
+ sky130_fd_sc_hd__dfrtp_4
X_16364_ obsg2.obstacleArray\[14\] obsg2.obstacleArray\[15\] net409 vssd1 vssd1 vccd1
+ vccd1 _02043_ sky130_fd_sc_hd__mux2_1
X_13576_ control.divider.count\[18\] _07949_ vssd1 vssd1 vccd1 vccd1 _07951_ sky130_fd_sc_hd__nand2_1
X_10788_ net1097 control.body\[629\] vssd1 vssd1 vccd1 vccd1 _05761_ sky130_fd_sc_hd__xor2_1
XFILLER_0_67_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18103_ obsg2.obstacleArray\[54\] _03684_ net524 vssd1 vssd1 vccd1 vccd1 _01305_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_82_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10063__A1 _04445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_59_Right_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_270 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11241__B net1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15315_ net2585 net74 _01588_ net2305 vssd1 vssd1 vccd1 vccd1 _00614_ sky130_fd_sc_hd__a22o_1
XFILLER_0_42_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14329__B2 net1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15929__A _05922_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12527_ net387 net306 _07460_ vssd1 vssd1 vccd1 vccd1 _07461_ sky130_fd_sc_hd__or3b_1
X_19083_ clknet_leaf_9_clk img_gen.tracker.next_frame\[521\] net1271 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[521\] sky130_fd_sc_hd__dfrtp_1
X_16295_ obsg2.obstacleArray\[114\] net406 vssd1 vssd1 vccd1 vccd1 _01974_ sky130_fd_sc_hd__or2_1
XANTENNA__10138__A net1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1115 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_966 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18034_ obsg2.obstacleArray\[30\] _03639_ net527 vssd1 vssd1 vccd1 vccd1 _01281_
+ sky130_fd_sc_hd__o21a_1
X_15246_ control.body\[776\] net99 _01579_ net2113 vssd1 vssd1 vccd1 vccd1 _00554_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_112_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12458_ net687 _07276_ _07300_ _07417_ vssd1 vssd1 vccd1 vccd1 net32 sky130_fd_sc_hd__a22o_1
XANTENNA__14552__B ag2.body\[68\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17279__B1 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11409_ _06372_ _06373_ _06375_ _06376_ vssd1 vssd1 vccd1 vccd1 _06382_ sky130_fd_sc_hd__a22o_1
XFILLER_0_111_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12389_ _07253_ _07291_ vssd1 vssd1 vccd1 vccd1 _07354_ sky130_fd_sc_hd__nor2_2
X_15177_ control.body\[843\] net101 _01571_ net2262 vssd1 vssd1 vccd1 vccd1 _00493_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_2_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_1326 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14128_ net843 ag2.body\[368\] ag2.body\[373\] net807 vssd1 vssd1 vccd1 vccd1 _08289_
+ sky130_fd_sc_hd__o22ai_1
X_19985_ clknet_leaf_64_clk _00929_ net1474 vssd1 vssd1 vccd1 vccd1 ag2.body\[415\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_103_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14501__A1 net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14501__B2 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14059_ net832 ag2.body\[33\] ag2.body\[34\] net824 _08217_ vssd1 vssd1 vccd1 vccd1
+ _08220_ sky130_fd_sc_hd__a221o_1
X_18936_ clknet_leaf_139_clk img_gen.tracker.next_frame\[374\] net1288 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[374\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__12640__X _07523_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18040__A _03542_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_68_Right_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16479__B net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09662__A net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1200 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18867_ clknet_leaf_17_clk img_gen.tracker.next_frame\[305\] net1342 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[305\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_118_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17451__B1 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17818_ _03481_ _03484_ vssd1 vssd1 vccd1 vccd1 _03485_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_94_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__20348__RESET_B net1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10601__A net1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18641__CLK clknet_leaf_131_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18798_ clknet_leaf_22_clk img_gen.tracker.next_frame\[236\] net1358 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[236\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_1400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11079__B1 net1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17749_ _02976_ _02983_ _03427_ _02712_ vssd1 vssd1 vccd1 vccd1 _03428_ sky130_fd_sc_hd__o211a_1
XANTENNA__12815__A1 net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10320__B net1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkload87_A clknet_leaf_105_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14568__A1 _03965_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19419_ clknet_leaf_108_clk _00363_ net1434 vssd1 vssd1 vccd1 vccd1 control.body\[969\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14568__B2 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_77_Right_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout148_A net154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16309__A2 net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1163 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13240__A1 net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09103_ ag2.body\[359\] vssd1 vssd1 vccd1 vccd1 _04128_ sky130_fd_sc_hd__inv_2
XFILLER_0_94_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16434__S net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10048__A _04551_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_966 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout315_A net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19147__CLK clknet_leaf_51_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09034_ ag2.body\[183\] vssd1 vssd1 vccd1 vccd1 _04059_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout1057_A net1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11578__S net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold320 img_gen.tracker.frame\[525\] vssd1 vssd1 vccd1 vccd1 net1882 sky130_fd_sc_hd__dlygate4sd3_1
Xhold331 img_gen.tracker.frame\[414\] vssd1 vssd1 vccd1 vccd1 net1893 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold342 img_gen.tracker.frame\[472\] vssd1 vssd1 vccd1 vccd1 net1904 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1224_A net1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold353 img_gen.tracker.frame\[412\] vssd1 vssd1 vccd1 vccd1 net1915 sky130_fd_sc_hd__dlygate4sd3_1
Xhold364 img_gen.tracker.frame\[479\] vssd1 vssd1 vccd1 vccd1 net1926 sky130_fd_sc_hd__dlygate4sd3_1
Xhold375 img_gen.tracker.frame\[19\] vssd1 vssd1 vccd1 vccd1 net1937 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout800 net805 vssd1 vssd1 vccd1 vccd1 net800 sky130_fd_sc_hd__buf_4
XFILLER_0_1_880 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold386 img_gen.tracker.frame\[242\] vssd1 vssd1 vccd1 vccd1 net1948 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout684_A _04393_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_86_Right_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout811 net813 vssd1 vssd1 vccd1 vccd1 net811 sky130_fd_sc_hd__clkbuf_4
Xhold397 img_gen.tracker.frame\[371\] vssd1 vssd1 vccd1 vccd1 net1959 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__17690__B1 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20125_ clknet_leaf_81_clk _01069_ net1485 vssd1 vssd1 vccd1 vccd1 ag2.body\[267\]
+ sky130_fd_sc_hd__dfrtp_4
Xfanout822 net823 vssd1 vssd1 vccd1 vccd1 net822 sky130_fd_sc_hd__buf_2
X_09936_ ag2.body\[26\] net1175 vssd1 vssd1 vccd1 vccd1 _04909_ sky130_fd_sc_hd__and2b_1
XANTENNA_fanout1012_X net1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout833 net835 vssd1 vssd1 vccd1 vccd1 net833 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_0_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout844 net846 vssd1 vssd1 vccd1 vccd1 net844 sky130_fd_sc_hd__clkbuf_4
Xfanout855 net856 vssd1 vssd1 vccd1 vccd1 net855 sky130_fd_sc_hd__clkbuf_4
Xfanout866 net867 vssd1 vssd1 vccd1 vccd1 net866 sky130_fd_sc_hd__clkbuf_4
X_20056_ clknet_leaf_72_clk _01000_ net1504 vssd1 vssd1 vccd1 vccd1 ag2.body\[342\]
+ sky130_fd_sc_hd__dfrtp_4
Xfanout877 net878 vssd1 vssd1 vccd1 vccd1 net877 sky130_fd_sc_hd__buf_4
XANTENNA_fanout851_A net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09867_ ag2.body\[158\] net1092 vssd1 vssd1 vccd1 vccd1 _04840_ sky130_fd_sc_hd__xor2_1
XANTENNA_fanout472_X net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11857__A2 net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout888 net889 vssd1 vssd1 vccd1 vccd1 net888 sky130_fd_sc_hd__buf_4
Xhold1020 control.body\[1102\] vssd1 vssd1 vccd1 vccd1 net2582 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout949_A net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1031 control.body\[802\] vssd1 vssd1 vccd1 vccd1 net2593 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout899 control.body_update.curr_length\[6\] vssd1 vssd1 vccd1 vccd1 net899 sky130_fd_sc_hd__clkbuf_4
Xhold1042 control.body\[916\] vssd1 vssd1 vccd1 vccd1 net2604 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13094__A net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1053 control.body\[1083\] vssd1 vssd1 vccd1 vccd1 net2615 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_73_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1064 control.body\[725\] vssd1 vssd1 vccd1 vccd1 net2626 sky130_fd_sc_hd__dlygate4sd3_1
X_09798_ _04767_ _04768_ _04769_ _04770_ vssd1 vssd1 vccd1 vccd1 _04771_ sky130_fd_sc_hd__or4_1
XFILLER_0_9_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_1388 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1075 control.body\[888\] vssd1 vssd1 vccd1 vccd1 net2637 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1086 control.body\[935\] vssd1 vssd1 vccd1 vccd1 net2648 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1097 control.body\[672\] vssd1 vssd1 vccd1 vccd1 net2659 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_115_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout737_X net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16609__S net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10230__B net1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11760_ img_gen.tracker.frame\[287\] net581 net542 img_gen.tracker.frame\[284\] _06731_
+ vssd1 vssd1 vccd1 vccd1 _06732_ sky130_fd_sc_hd__o221a_1
XFILLER_0_51_1506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11045__C _05936_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_95_Right_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10711_ _05676_ _05677_ _05678_ _05683_ vssd1 vssd1 vccd1 vccd1 _05684_ sky130_fd_sc_hd__or4_1
XFILLER_0_67_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14559__A1 net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14559__B2 net1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11691_ img_gen.tracker.frame\[98\] net618 net585 img_gen.tracker.frame\[107\] vssd1
+ vssd1 vccd1 vccd1 _06663_ sky130_fd_sc_hd__o22a_1
XFILLER_0_138_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12438__A net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_639 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14912__A_N _05375_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10642_ _05611_ _05612_ _05613_ _05614_ vssd1 vssd1 vccd1 vccd1 _05615_ sky130_fd_sc_hd__or4_1
X_13430_ net388 _07460_ _07813_ vssd1 vssd1 vccd1 vccd1 _07884_ sky130_fd_sc_hd__and3_1
XANTENNA__12034__A2 net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11061__B net1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13361_ net274 _07856_ _07857_ net1671 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[461\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__15749__A _05255_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10573_ ag2.body\[188\] net1138 vssd1 vssd1 vccd1 vccd1 _05546_ sky130_fd_sc_hd__xor2_1
XANTENNA__14653__A net1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16344__S net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15100_ control.body\[918\] net145 _01563_ net2194 vssd1 vssd1 vccd1 vccd1 _00424_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_107_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12312_ _07228_ _07202_ _07210_ vssd1 vssd1 vccd1 vccd1 _07279_ sky130_fd_sc_hd__or3b_1
XFILLER_0_49_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16080_ net346 _01758_ _01755_ _01742_ vssd1 vssd1 vccd1 vccd1 _01759_ sky130_fd_sc_hd__o211a_1
XFILLER_0_90_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13292_ net280 _07829_ _07830_ net1736 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[419\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_122_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16720__A2 net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17493__A2_N net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1024 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12243_ _07193_ _07212_ img_gen.updater.commands.count\[14\] img_gen.updater.commands.count\[15\]
+ img_gen.updater.commands.count\[13\] vssd1 vssd1 vccd1 vccd1 _07213_ sky130_fd_sc_hd__o2111a_1
X_15031_ _04445_ _04607_ _01556_ vssd1 vssd1 vccd1 vccd1 _01557_ sky130_fd_sc_hd__a21boi_4
XANTENNA__13269__A net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17964__A net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_2_Left_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12173__A net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11545__A1 net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_39_Left_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12174_ net385 _07119_ _06823_ vssd1 vssd1 vccd1 vccd1 _07146_ sky130_fd_sc_hd__o21ba_2
X_20593__1525 vssd1 vssd1 vccd1 vccd1 _20593__1525/HI net1525 sky130_fd_sc_hd__conb_1
XANTENNA__18473__A2 net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1360 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11125_ net1149 control.body\[867\] vssd1 vssd1 vccd1 vccd1 _06098_ sky130_fd_sc_hd__and2b_1
XFILLER_0_101_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19770_ clknet_leaf_18_clk _00714_ net1323 vssd1 vssd1 vccd1 vccd1 ag2.body\[616\]
+ sky130_fd_sc_hd__dfrtp_2
X_16982_ _02653_ _02654_ _02655_ _02657_ vssd1 vssd1 vccd1 vccd1 _02661_ sky130_fd_sc_hd__and4_1
XFILLER_0_120_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18721_ clknet_leaf_142_clk img_gen.tracker.next_frame\[159\] net1253 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[159\] sky130_fd_sc_hd__dfrtp_1
X_11056_ ag2.body\[437\] net1103 vssd1 vssd1 vccd1 vccd1 _06029_ sky130_fd_sc_hd__xnor2_1
X_15933_ ag2.body\[171\] net136 _01655_ ag2.body\[163\] vssd1 vssd1 vccd1 vccd1 _01165_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_95_1411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17433__B1 net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10007_ net898 net901 vssd1 vssd1 vccd1 vccd1 _04980_ sky130_fd_sc_hd__and2b_2
X_18652_ clknet_leaf_131_clk img_gen.tracker.next_frame\[90\] net1317 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[90\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__11517__A net1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10421__A net1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15864_ ag2.body\[239\] net175 _01646_ ag2.body\[231\] vssd1 vssd1 vccd1 vccd1 _01105_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_91_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10520__A2 net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17603_ ag2.body\[421\] net949 vssd1 vssd1 vccd1 vccd1 _03282_ sky130_fd_sc_hd__xor2_1
XFILLER_0_118_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14815_ net1018 ag2.body\[382\] vssd1 vssd1 vccd1 vccd1 _01486_ sky130_fd_sc_hd__or2_1
XANTENNA__11236__B net1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18583_ clknet_leaf_4_clk img_gen.tracker.next_frame\[21\] net1278 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[21\] sky130_fd_sc_hd__dfrtp_1
X_15795_ ag2.body\[288\] net207 _01640_ ag2.body\[280\] vssd1 vssd1 vccd1 vccd1 _01042_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_118_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_48_Left_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10808__B1 _05765_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17534_ _03207_ _03208_ _03209_ _03210_ _03212_ vssd1 vssd1 vccd1 vccd1 _03213_ sky130_fd_sc_hd__a221o_1
X_14746_ net1038 ag2.body\[108\] vssd1 vssd1 vccd1 vccd1 _08907_ sky130_fd_sc_hd__xor2_1
XFILLER_0_86_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11958_ net466 _06928_ _06929_ _06902_ _06903_ vssd1 vssd1 vccd1 vccd1 _06930_ sky130_fd_sc_hd__o32a_1
XTAP_TAPCELL_ROW_120_3990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10909_ _05878_ _05879_ _05880_ _05881_ vssd1 vssd1 vccd1 vccd1 _05882_ sky130_fd_sc_hd__or4_1
X_17465_ ag2.body\[535\] net932 vssd1 vssd1 vccd1 vccd1 _03144_ sky130_fd_sc_hd__xor2_1
XFILLER_0_58_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14677_ net1028 ag2.body\[389\] vssd1 vssd1 vccd1 vccd1 _08838_ sky130_fd_sc_hd__or2_1
XANTENNA__12348__A net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11889_ img_gen.tracker.frame\[37\] net623 net552 img_gen.tracker.frame\[43\] _06860_
+ vssd1 vssd1 vccd1 vccd1 _06861_ sky130_fd_sc_hd__o221a_1
X_19204_ clknet_leaf_88_clk _00148_ net1459 vssd1 vssd1 vccd1 vccd1 ag2.body\[67\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_55_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16416_ obsg2.obstacleArray\[112\] obsg2.obstacleArray\[113\] net455 vssd1 vssd1
+ vccd1 vccd1 _02095_ sky130_fd_sc_hd__mux2_1
X_13628_ _07992_ _07993_ vssd1 vssd1 vccd1 vccd1 control.divider.next_count\[9\] sky130_fd_sc_hd__nor2_1
XFILLER_0_104_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17396_ ag2.body\[504\] net739 net700 ag2.body\[510\] _03074_ vssd1 vssd1 vccd1 vccd1
+ _03075_ sky130_fd_sc_hd__a221o_1
XANTENNA__12025__A2 net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19135_ clknet_leaf_132_clk img_gen.tracker.next_frame\[573\] net1297 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[573\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__09977__A1 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16347_ _02024_ _02025_ net417 vssd1 vssd1 vccd1 vccd1 _02026_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09977__B2 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16254__S net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13559_ ssdec1.in\[2\] _07938_ vssd1 vssd1 vccd1 vccd1 _07940_ sky130_fd_sc_hd__nand2_1
XFILLER_0_55_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14563__A net1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_max_cap368_X net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19066_ clknet_leaf_29_clk img_gen.tracker.next_frame\[504\] net1335 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[504\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16278_ obsg2.obstacleArray\[19\] net414 _01956_ net417 vssd1 vssd1 vccd1 vccd1 _01957_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_120_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18017_ _03540_ _03581_ vssd1 vssd1 vccd1 vccd1 _03627_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_57_Left_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15229_ net2447 net96 _01577_ control.body\[785\] vssd1 vssd1 vccd1 vccd1 _00539_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_114_3794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12083__A net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_110_3669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10315__B net1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout107 net114 vssd1 vssd1 vccd1 vccd1 net107 sky130_fd_sc_hd__buf_2
Xfanout118 net119 vssd1 vssd1 vccd1 vccd1 net118 sky130_fd_sc_hd__buf_2
Xfanout129 net132 vssd1 vssd1 vccd1 vccd1 net129 sky130_fd_sc_hd__buf_2
X_19968_ clknet_leaf_62_clk _00912_ net1469 vssd1 vssd1 vccd1 vccd1 ag2.body\[430\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_10_499 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1620 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09721_ _04669_ _04679_ _04693_ vssd1 vssd1 vccd1 vccd1 _04694_ sky130_fd_sc_hd__o21a_1
X_18919_ clknet_leaf_145_clk img_gen.tracker.next_frame\[357\] net1253 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[357\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__11839__A2 net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16002__B net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19899_ clknet_leaf_86_clk _00843_ net1464 vssd1 vssd1 vccd1 vccd1 ag2.body\[489\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_78_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17424__B1 net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_1506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09652_ net1220 control.body\[744\] vssd1 vssd1 vccd1 vccd1 _04625_ sky130_fd_sc_hd__xor2_1
XANTENNA__16778__A2 net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16937__B net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09583_ _04238_ _04471_ vssd1 vssd1 vccd1 vccd1 _04556_ sky130_fd_sc_hd__or2_2
XFILLER_0_96_219 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10050__B _04962_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16429__S net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09466__A2_N net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17727__A1 net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16953__A ag2.body\[290\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1174_A net1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12016__A2 net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16950__A2 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16164__S net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18152__A1 net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1341_A net1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout318_X net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1439_A net1442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16163__B1 net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16702__A2 net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14192__B ag2.body\[165\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_947 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09017_ ag2.body\[148\] vssd1 vssd1 vccd1 vccd1 _04042_ sky130_fd_sc_hd__inv_2
XFILLER_0_115_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14713__A1 net993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13089__A net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14713__B2 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10506__A net1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1227_X net1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold150 obsg2.obsNeeded\[1\] vssd1 vssd1 vccd1 vccd1 net1712 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold161 img_gen.tracker.frame\[113\] vssd1 vssd1 vccd1 vccd1 net1723 sky130_fd_sc_hd__dlygate4sd3_1
Xhold172 img_gen.tracker.frame\[118\] vssd1 vssd1 vccd1 vccd1 net1734 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10225__B net1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout687_X net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold183 img_gen.tracker.frame\[405\] vssd1 vssd1 vccd1 vccd1 net1745 sky130_fd_sc_hd__dlygate4sd3_1
Xhold194 img_gen.tracker.frame\[400\] vssd1 vssd1 vccd1 vccd1 net1756 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12721__A net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout630 _06473_ vssd1 vssd1 vccd1 vccd1 net630 sky130_fd_sc_hd__clkbuf_4
X_20108_ clknet_leaf_79_clk _01052_ net1487 vssd1 vssd1 vccd1 vccd1 ag2.body\[282\]
+ sky130_fd_sc_hd__dfrtp_4
Xfanout641 _04419_ vssd1 vssd1 vccd1 vccd1 net641 sky130_fd_sc_hd__buf_4
X_09919_ _04103_ net1236 net1212 _04104_ vssd1 vssd1 vccd1 vccd1 _04892_ sky130_fd_sc_hd__a22o_1
Xfanout652 net653 vssd1 vssd1 vccd1 vccd1 net652 sky130_fd_sc_hd__clkbuf_2
Xfanout663 _04394_ vssd1 vssd1 vccd1 vccd1 net663 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout854_X net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout674 _04393_ vssd1 vssd1 vccd1 vccd1 net674 sky130_fd_sc_hd__clkbuf_4
Xfanout685 net686 vssd1 vssd1 vccd1 vccd1 net685 sky130_fd_sc_hd__clkbuf_4
XANTENNA__17415__B1 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20039_ clknet_leaf_66_clk _00983_ net1476 vssd1 vssd1 vccd1 vccd1 ag2.body\[357\]
+ sky130_fd_sc_hd__dfrtp_4
Xfanout696 _04268_ vssd1 vssd1 vccd1 vccd1 net696 sky130_fd_sc_hd__clkbuf_4
XANTENNA_clkbuf_3_1_0_clk_X clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12930_ net679 _07662_ vssd1 vssd1 vccd1 vccd1 _07663_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_124_4090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16769__A2 net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16847__B net961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11056__B net1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12861_ net240 _07631_ _07632_ net1766 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[186\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__16339__S net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14600_ net829 ag2.body\[306\] _04102_ net1012 _08754_ vssd1 vssd1 vccd1 vccd1 _08761_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_90_1330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11812_ img_gen.tracker.frame\[464\] net540 _06783_ net558 vssd1 vssd1 vccd1 vccd1
+ _06784_ sky130_fd_sc_hd__o211a_1
XFILLER_0_55_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15580_ ag2.body\[480\] net130 _01617_ ag2.body\[472\] vssd1 vssd1 vccd1 vccd1 _00850_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__13452__A1 net235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12792_ net667 _07599_ vssd1 vssd1 vccd1 vccd1 _07600_ sky130_fd_sc_hd__nor2_1
XFILLER_0_96_786 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11463__B1 net1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14531_ net983 ag2.body\[250\] vssd1 vssd1 vccd1 vccd1 _08692_ sky130_fd_sc_hd__or2_1
XFILLER_0_132_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17959__A net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11743_ img_gen.tracker.frame\[5\] net606 net590 img_gen.tracker.frame\[11\] _06714_
+ vssd1 vssd1 vccd1 vccd1 _06715_ sky130_fd_sc_hd__o221a_1
XFILLER_0_95_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17250_ net723 ag2.body\[546\] _04200_ net874 vssd1 vssd1 vccd1 vccd1 _02929_ sky130_fd_sc_hd__a2bb2o_1
X_14462_ _08615_ _08617_ _08620_ _08622_ vssd1 vssd1 vccd1 vccd1 _08623_ sky130_fd_sc_hd__or4_2
XANTENNA__13204__A1 net242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12007__A2 net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_4495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11674_ _06641_ _06644_ vssd1 vssd1 vccd1 vccd1 _06646_ sky130_fd_sc_hd__xnor2_1
XANTENNA__16941__A2 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16201_ obsg2.obstacleArray\[42\] obsg2.obstacleArray\[43\] net422 vssd1 vssd1 vccd1
+ vccd1 _01880_ sky130_fd_sc_hd__mux2_1
X_13413_ net257 _07876_ _07877_ net1699 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[493\]
+ sky130_fd_sc_hd__a22o_1
X_17181_ ag2.body\[461\] net948 vssd1 vssd1 vccd1 vccd1 _02860_ sky130_fd_sc_hd__xor2_1
XFILLER_0_92_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10625_ _03992_ net1177 net1102 _03993_ _05592_ vssd1 vssd1 vccd1 vccd1 _05598_ sky130_fd_sc_hd__a221o_1
XFILLER_0_10_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14393_ net1032 ag2.body\[125\] vssd1 vssd1 vccd1 vccd1 _08554_ sky130_fd_sc_hd__xnor2_1
X_16132_ _01743_ _01806_ _01810_ _01728_ vssd1 vssd1 vccd1 vccd1 _01811_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_12_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16154__B1 net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13344_ net228 _07850_ _07851_ net1894 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[450\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_49_1254 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10556_ _04553_ _05509_ _05526_ _05528_ vssd1 vssd1 vccd1 vccd1 _05529_ sky130_fd_sc_hd__o22a_1
XFILLER_0_126_1411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16063_ _01727_ _01741_ vssd1 vssd1 vccd1 vccd1 _01742_ sky130_fd_sc_hd__and2_2
XFILLER_0_11_208 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13275_ net234 _07823_ _07824_ net1701 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[408\]
+ sky130_fd_sc_hd__a22o_1
X_10487_ ag2.body\[585\] net1196 vssd1 vssd1 vccd1 vccd1 _05460_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_51_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_254 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15014_ control.body\[986\] net168 _01553_ control.body\[978\] vssd1 vssd1 vccd1
+ vccd1 _00348_ sky130_fd_sc_hd__a22o_1
X_12226_ img_gen.updater.commands.cmd_num\[1\] img_gen.updater.commands.cmd_num\[0\]
+ vssd1 vssd1 vccd1 vccd1 _07196_ sky130_fd_sc_hd__nand2_1
XANTENNA__16457__A1 net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12157_ img_gen.tracker.frame\[459\] net597 net578 img_gen.tracker.frame\[465\] vssd1
+ vssd1 vccd1 vccd1 _07129_ sky130_fd_sc_hd__o22a_1
X_19822_ clknet_leaf_125_clk _00766_ net1411 vssd1 vssd1 vccd1 vccd1 ag2.body\[572\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_62_1487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09924__B _04640_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11108_ net1207 control.body\[1097\] vssd1 vssd1 vccd1 vccd1 _06081_ sky130_fd_sc_hd__nand2b_1
X_16965_ ag2.body\[414\] net940 vssd1 vssd1 vccd1 vccd1 _02644_ sky130_fd_sc_hd__xor2_1
X_19753_ clknet_leaf_130_clk net2445 net1317 vssd1 vssd1 vccd1 vccd1 control.body\[647\]
+ sky130_fd_sc_hd__dfrtp_1
X_12088_ img_gen.tracker.frame\[303\] net612 net595 img_gen.tracker.frame\[309\] _07059_
+ vssd1 vssd1 vccd1 vccd1 _07060_ sky130_fd_sc_hd__a221o_1
X_15916_ ag2.body\[189\] net131 _01652_ ag2.body\[181\] vssd1 vssd1 vccd1 vccd1 _01151_
+ sky130_fd_sc_hd__a22o_1
X_11039_ net1231 control.body\[1040\] vssd1 vssd1 vccd1 vccd1 _06012_ sky130_fd_sc_hd__nand2b_1
X_18704_ clknet_leaf_10_clk img_gen.tracker.next_frame\[142\] net1274 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[142\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__10151__A ag2.body\[57\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19684_ clknet_leaf_117_clk _00628_ net1384 vssd1 vssd1 vccd1 vccd1 control.body\[706\]
+ sky130_fd_sc_hd__dfrtp_1
X_16896_ ag2.body\[211\] net719 net706 ag2.body\[213\] vssd1 vssd1 vccd1 vccd1 _02575_
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_56_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18635_ clknet_leaf_131_clk img_gen.tracker.next_frame\[73\] net1295 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[73\] sky130_fd_sc_hd__dfrtp_1
X_15847_ _04688_ net59 vssd1 vssd1 vccd1 vccd1 _01645_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_103_3451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_103_3462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18566_ clknet_leaf_14_clk img_gen.tracker.next_frame\[4\] net1313 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[4\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_103_3473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15778_ ag2.body\[305\] net210 _01638_ ag2.body\[297\] vssd1 vssd1 vccd1 vccd1 _01027_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_91_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13443__A1 net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13181__B net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17517_ _03188_ _03191_ _03194_ _03195_ vssd1 vssd1 vccd1 vccd1 _03196_ sky130_fd_sc_hd__or4_1
X_14729_ net821 ag2.body\[115\] _04027_ net1012 vssd1 vssd1 vccd1 vccd1 _08890_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__11454__B1 _06413_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18497_ net1515 net1509 vssd1 vssd1 vccd1 vccd1 _00028_ sky130_fd_sc_hd__or2_1
XANTENNA__19805__CLK clknet_leaf_124_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1578 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17448_ _04136_ net960 net691 ag2.body\[383\] _03122_ vssd1 vssd1 vccd1 vccd1 _03127_
+ sky130_fd_sc_hd__a221o_1
XANTENNA__16393__B1 net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_458 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17379_ ag2.body\[491\] net853 vssd1 vssd1 vccd1 vccd1 _03058_ sky130_fd_sc_hd__xor2_1
XANTENNA__12806__A net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_508 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_3856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_65_Left_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_116_3867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19118_ clknet_leaf_131_clk img_gen.tracker.next_frame\[556\] net1295 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[556\] sky130_fd_sc_hd__dfrtp_1
X_20390_ clknet_leaf_40_clk _01277_ net1374 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[26\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__15499__A2 net113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19049_ clknet_leaf_10_clk img_gen.tracker.next_frame\[487\] net1275 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[487\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17754__D _03432_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16448__A1 net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18212__B net40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17891__X _03531_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10613__X _05586_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12541__A net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_2484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_1005 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_2495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_74_Left_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09704_ _04663_ _04664_ _04667_ _04668_ vssd1 vssd1 vccd1 vccd1 _04677_ sky130_fd_sc_hd__a22o_1
XFILLER_0_39_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19335__CLK clknet_leaf_103_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16667__B net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_88_2992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11693__B1 net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_4_clk_A clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09635_ net1206 _04251_ control.body\[1019\] net771 _04607_ vssd1 vssd1 vccd1 vccd1
+ _04608_ sky130_fd_sc_hd__a221o_1
XANTENNA__16159__S net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10996__A ag2.body\[341\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14468__A net1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1291_A net1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout268_X net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout647_A net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1389_A net1404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13372__A net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_2878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13434__A1 net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09566_ net908 _04446_ net641 vssd1 vssd1 vccd1 vccd1 _04539_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_84_2889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14187__B ag2.body\[166\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13091__B net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_65_2299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09497_ net909 net913 vssd1 vssd1 vccd1 vccd1 _04470_ sky130_fd_sc_hd__or2_4
XANTENNA_fanout814_A net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20592__1524 vssd1 vssd1 vccd1 vccd1 _20592__1524/HI net1524 sky130_fd_sc_hd__conb_1
XANTENNA_fanout1177_X net1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11540__S0 net1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09849__X _04822_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17498__B net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_83_Left_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout602_X net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12716__A net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10410_ net1112 control.body\[1077\] vssd1 vssd1 vccd1 vccd1 _05383_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_22_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16136__B1 net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11390_ _06359_ _06360_ _06361_ _06362_ vssd1 vssd1 vccd1 vccd1 _06363_ sky130_fd_sc_hd__a22o_1
X_20588_ net1520 vssd1 vssd1 vccd1 vccd1 gpio_oeb[0] sky130_fd_sc_hd__buf_2
XANTENNA__09810__B1 _04782_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16687__A1 net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17718__S net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10341_ ag2.body\[522\] net775 net1059 _04192_ _05313_ vssd1 vssd1 vccd1 vccd1 _05314_
+ sky130_fd_sc_hd__a221o_1
XANTENNA__17884__B1 _03523_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13060_ net680 _07723_ vssd1 vssd1 vccd1 vccd1 _07724_ sky130_fd_sc_hd__nor2_1
XFILLER_0_131_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10272_ ag2.body\[137\] net1211 vssd1 vssd1 vccd1 vccd1 _05245_ sky130_fd_sc_hd__xor2_1
XANTENNA__11484__A_N _06122_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout971_X net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16439__A1 net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12011_ _06964_ _06970_ _06976_ _06982_ net471 net440 vssd1 vssd1 vccd1 vccd1 _06983_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__13547__A net226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09744__B net1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1403 net1404 vssd1 vssd1 vccd1 vccd1 net1403 sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_92_Left_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1414 net1415 vssd1 vssd1 vccd1 vccd1 net1414 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_126_4152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1425 net1430 vssd1 vssd1 vccd1 vccd1 net1425 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_54_1970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1436 net1442 vssd1 vssd1 vccd1 vccd1 net1436 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_126_4163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1447 net1448 vssd1 vssd1 vccd1 vccd1 net1447 sky130_fd_sc_hd__clkbuf_2
Xfanout460 _01710_ vssd1 vssd1 vccd1 vccd1 net460 sky130_fd_sc_hd__clkbuf_8
Xfanout1458 net1465 vssd1 vssd1 vccd1 vccd1 net1458 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_35_1380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1469 net1470 vssd1 vssd1 vccd1 vccd1 net1469 sky130_fd_sc_hd__clkbuf_4
Xfanout471 net472 vssd1 vssd1 vccd1 vccd1 net471 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_35_1391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16750_ obsg2.obstacleArray\[60\] net491 net482 obsg2.obstacleArray\[61\] vssd1 vssd1
+ vccd1 vccd1 _02429_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_122_4038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout482 net483 vssd1 vssd1 vccd1 vccd1 net482 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_50_1856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout493 _01736_ vssd1 vssd1 vccd1 vccd1 net493 sky130_fd_sc_hd__buf_4
X_13962_ ag2.body\[102\] net189 _08156_ ag2.body\[94\] vssd1 vssd1 vccd1 vccd1 _00183_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_6_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_4049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15701_ ag2.body\[382\] net140 _01628_ ag2.body\[374\] vssd1 vssd1 vccd1 vccd1 _00960_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_96_1583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12913_ net679 _07654_ vssd1 vssd1 vccd1 vccd1 _07655_ sky130_fd_sc_hd__nor2_1
X_16681_ _02227_ _02345_ _02349_ _02359_ _02211_ vssd1 vssd1 vccd1 vccd1 _02360_ sky130_fd_sc_hd__a311o_1
XANTENNA__11684__B1 net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14378__A net1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16069__S net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13893_ ag2.body\[40\] net118 _08149_ ag2.body\[32\] vssd1 vssd1 vccd1 vccd1 _00121_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__19828__CLK clknet_leaf_124_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11354__X _06327_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16072__C1 _01743_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18420_ _03857_ _03909_ net434 vssd1 vssd1 vccd1 vccd1 _03910_ sky130_fd_sc_hd__a21oi_1
X_15632_ _06028_ net64 vssd1 vssd1 vccd1 vccd1 _01622_ sky130_fd_sc_hd__and2_2
XFILLER_0_9_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12844_ net1767 _07623_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[178\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_70_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18351_ _04645_ _08033_ vssd1 vssd1 vccd1 vccd1 _03847_ sky130_fd_sc_hd__or2_1
XFILLER_0_55_1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15563_ ag2.body\[498\] net185 _01614_ ag2.body\[490\] vssd1 vssd1 vccd1 vccd1 _00836_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_48_1774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_263 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1182 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12775_ net2034 net647 _07590_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[142\]
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_48_1785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17167__A2 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17302_ _02973_ _02974_ _02977_ _02978_ _02980_ vssd1 vssd1 vccd1 vccd1 _02981_ sky130_fd_sc_hd__a221o_1
XFILLER_0_84_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_48_1796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14514_ net985 ag2.body\[314\] vssd1 vssd1 vccd1 vccd1 _08675_ sky130_fd_sc_hd__xor2_1
XFILLER_0_127_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18282_ net319 _03583_ obsg2.obstacleArray\[138\] vssd1 vssd1 vccd1 vccd1 _03780_
+ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_29_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11726_ img_gen.tracker.frame\[194\] net624 vssd1 vssd1 vccd1 vccd1 _06698_ sky130_fd_sc_hd__or2_1
X_15494_ ag2.body\[565\] net110 _01606_ ag2.body\[557\] vssd1 vssd1 vccd1 vccd1 _00775_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_51_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17233_ _04156_ net883 net703 ag2.body\[445\] vssd1 vssd1 vccd1 vccd1 _02912_ sky130_fd_sc_hd__a22o_1
XANTENNA__16470__S0 net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14445_ net1038 ag2.body\[228\] vssd1 vssd1 vccd1 vccd1 _08606_ sky130_fd_sc_hd__xor2_1
X_11657_ net1119 net1094 vssd1 vssd1 vccd1 vccd1 _06630_ sky130_fd_sc_hd__nand2_2
XANTENNA__12626__A net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10608_ net1110 control.body\[989\] vssd1 vssd1 vccd1 vccd1 _05581_ sky130_fd_sc_hd__xor2_1
X_17164_ ag2.body\[592\] net879 vssd1 vssd1 vccd1 vccd1 _02843_ sky130_fd_sc_hd__or2_1
X_14376_ net834 ag2.body\[417\] ag2.body\[423\] net793 _08532_ vssd1 vssd1 vccd1 vccd1
+ _08537_ sky130_fd_sc_hd__a221o_1
XFILLER_0_29_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11588_ _06506_ _06557_ _06559_ vssd1 vssd1 vccd1 vccd1 _06561_ sky130_fd_sc_hd__and3_1
XFILLER_0_40_815 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16115_ _01742_ _01789_ _01793_ _01729_ vssd1 vssd1 vccd1 vccd1 _01794_ sky130_fd_sc_hd__a31o_1
XANTENNA__16678__A1 net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_94_3185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_3720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_3196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold908 control.body\[713\] vssd1 vssd1 vccd1 vccd1 net2470 sky130_fd_sc_hd__dlygate4sd3_1
X_13327_ _06823_ _07502_ vssd1 vssd1 vccd1 vccd1 _07844_ sky130_fd_sc_hd__nor2_1
X_17095_ ag2.body\[296\] net886 vssd1 vssd1 vccd1 vccd1 _02774_ sky130_fd_sc_hd__nand2_1
Xhold919 control.body\[909\] vssd1 vssd1 vccd1 vccd1 net2481 sky130_fd_sc_hd__dlygate4sd3_1
X_10539_ ag2.body\[226\] net1182 vssd1 vssd1 vccd1 vccd1 _05512_ sky130_fd_sc_hd__xor2_1
XFILLER_0_10_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16046_ net956 _01717_ vssd1 vssd1 vccd1 vccd1 _01725_ sky130_fd_sc_hd__and2_2
X_13258_ net310 _07449_ vssd1 vssd1 vccd1 vccd1 _07817_ sky130_fd_sc_hd__nor2_1
XFILLER_0_62_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18032__B net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17627__B1 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12209_ score_detect.sig_out\[0\] _04271_ _04948_ vssd1 vssd1 vccd1 vccd1 _07181_
+ sky130_fd_sc_hd__o21ai_4
X_13189_ net289 _07783_ _07784_ net1801 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[362\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__17722__S0 net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19805_ clknet_leaf_124_clk _00749_ net1405 vssd1 vssd1 vccd1 vccd1 ag2.body\[587\]
+ sky130_fd_sc_hd__dfrtp_4
X_17997_ obsg2.obstacleArray\[20\] _03612_ net533 vssd1 vssd1 vccd1 vccd1 _01271_
+ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_109_3660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15653__A2 net139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16948_ ag2.body\[385\] net872 vssd1 vssd1 vccd1 vccd1 _02627_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_105_3513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19736_ clknet_leaf_132_clk _00680_ net1305 vssd1 vssd1 vccd1 vccd1 control.body\[662\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_105_3524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20335__CLK clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12011__S1 net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_3535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10478__A1 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16879_ ag2.body\[21\] net946 vssd1 vssd1 vccd1 vccd1 _02558_ sky130_fd_sc_hd__xor2_1
X_19667_ clknet_leaf_119_clk _00611_ net1390 vssd1 vssd1 vccd1 vccd1 control.body\[721\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14288__A net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_1201 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09420_ ag2.goodColl net530 _04398_ vssd1 vssd1 vccd1 vccd1 _04399_ sky130_fd_sc_hd__and3_1
XFILLER_0_56_1055 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18618_ clknet_leaf_145_clk img_gen.tracker.next_frame\[56\] net1241 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[56\] sky130_fd_sc_hd__dfrtp_1
X_19598_ clknet_leaf_118_clk _00542_ net1393 vssd1 vssd1 vccd1 vccd1 control.body\[796\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_133_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__20485__CLK clknet_leaf_37_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09351_ net270 _04352_ _04353_ vssd1 vssd1 vccd1 vccd1 _01421_ sky130_fd_sc_hd__and3_1
X_18549_ clknet_leaf_131_clk _00075_ net1297 vssd1 vssd1 vccd1 vccd1 ag2.y\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_133_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18355__B2 net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_959 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_118_3907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_118_3918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09282_ sound_gen.posDetector1.N\[1\] sound_gen.posDetector1.N\[0\] sound_gen.osc1.keepCounting
+ vssd1 vssd1 vccd1 vccd1 _04305_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_118_3929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_2141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_2152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_2163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20511_ clknet_leaf_113_clk track.nextHighScore\[1\] net1403 vssd1 vssd1 vccd1 vccd1
+ track.highScore\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16008__A net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout228_A net233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20442_ clknet_leaf_25_clk _01329_ net1345 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[78\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_16_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1102 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_2660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20373_ clknet_leaf_23_clk _01260_ net1362 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[9\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_77_2671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15847__A _04688_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16442__S net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_2682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload70 clknet_leaf_46_clk vssd1 vssd1 vccd1 vccd1 clkload70/Y sky130_fd_sc_hd__inv_8
XTAP_TAPCELL_ROW_73_2535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1137_A net1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_2081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload81 clknet_leaf_92_clk vssd1 vssd1 vccd1 vccd1 clkload81/Y sky130_fd_sc_hd__inv_6
XTAP_TAPCELL_ROW_58_2092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload92 clknet_leaf_110_clk vssd1 vssd1 vccd1 vccd1 clkload92/Y sky130_fd_sc_hd__bufinv_16
XFILLER_0_11_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_1347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout597_A net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11439__X _06412_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13367__A net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17618__B1 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09564__B _04239_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17713__S0 net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08997_ ag2.body\[95\] vssd1 vssd1 vccd1 vccd1 _04022_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout764_A net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18725__CLK clknet_leaf_142_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout385_X net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15644__A2 net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_3_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09859__B1 _04831_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout931_A obsg2.randCord\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14198__A net1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout552_X net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09618_ net1170 control.body\[802\] vssd1 vssd1 vccd1 vccd1 _04591_ sky130_fd_sc_hd__xor2_1
XANTENNA__13407__A1 net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout43_A net44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1128 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10890_ net1146 control.body\[651\] vssd1 vssd1 vccd1 vccd1 _05863_ sky130_fd_sc_hd__nand2_1
XANTENNA__18875__CLK clknet_leaf_13_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09549_ _04445_ net637 _04520_ vssd1 vssd1 vccd1 vccd1 _04522_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout1461_X net1461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1498 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout817_X net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11902__X _06874_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_134_4410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12560_ net612 _06638_ net436 net576 vssd1 vssd1 vccd1 vccd1 _07479_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_134_4421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18117__B _03693_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11511_ _06480_ _06481_ vssd1 vssd1 vccd1 vccd1 _06484_ sky130_fd_sc_hd__xnor2_1
XANTENNA__17021__B net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09739__B net1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12491_ _07431_ _07439_ vssd1 vssd1 vccd1 vccd1 _07440_ sky130_fd_sc_hd__nor2_1
XFILLER_0_47_992 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14230_ _08389_ _08390_ vssd1 vssd1 vccd1 vccd1 _08391_ sky130_fd_sc_hd__or2_1
XANTENNA__16109__B1 net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11442_ net1204 control.body\[953\] vssd1 vssd1 vccd1 vccd1 _06415_ sky130_fd_sc_hd__xor2_1
XFILLER_0_46_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11373_ ag2.body\[476\] net1128 vssd1 vssd1 vccd1 vccd1 _06346_ sky130_fd_sc_hd__xor2_1
XFILLER_0_81_1104 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14161_ net832 ag2.body\[617\] ag2.body\[616\] net840 vssd1 vssd1 vccd1 vccd1 _08322_
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_85_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17321__A2 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14661__A net1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10944__A2 net1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10324_ ag2.body\[615\] net1047 vssd1 vssd1 vccd1 vccd1 _05297_ sky130_fd_sc_hd__xor2_1
X_13112_ net2127 net652 _07748_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[321\]
+ sky130_fd_sc_hd__and3_1
XANTENNA__19500__CLK clknet_leaf_115_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14092_ net1002 ag2.body\[280\] vssd1 vssd1 vccd1 vccd1 _08253_ sky130_fd_sc_hd__xor2_1
XFILLER_0_24_1500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_128_4214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_4225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_1571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_128_4236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17920_ net345 _03553_ vssd1 vssd1 vccd1 vccd1 _03554_ sky130_fd_sc_hd__nor2_2
XANTENNA__17972__A net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10255_ net1075 control.body\[790\] vssd1 vssd1 vccd1 vccd1 _05228_ sky130_fd_sc_hd__xor2_1
X_13043_ net342 _07546_ vssd1 vssd1 vccd1 vccd1 _07716_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_37_1442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10157__B1 _04232_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12181__A net1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1200 ag2.y\[1\] vssd1 vssd1 vccd1 vccd1 net1200 sky130_fd_sc_hd__buf_2
Xfanout1211 net1212 vssd1 vssd1 vccd1 vccd1 net1211 sky130_fd_sc_hd__clkbuf_8
X_17851_ img_gen.updater.commands.rR1.rainbowRNG\[14\] _03506_ vssd1 vssd1 vccd1 vccd1
+ _03507_ sky130_fd_sc_hd__nand2_1
XFILLER_0_24_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09562__A2 _04518_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17691__B net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10186_ ag2.body\[420\] net1139 vssd1 vssd1 vccd1 vccd1 _05159_ sky130_fd_sc_hd__xor2_1
XFILLER_0_79_1022 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1222 net1224 vssd1 vssd1 vccd1 vccd1 net1222 sky130_fd_sc_hd__clkbuf_4
Xfanout1233 net1238 vssd1 vssd1 vccd1 vccd1 net1233 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_33_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1244 net1250 vssd1 vssd1 vccd1 vccd1 net1244 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10413__B _05375_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16802_ _02086_ _02107_ _02170_ _02480_ vssd1 vssd1 vccd1 vccd1 _02481_ sky130_fd_sc_hd__or4_1
Xfanout1255 net1257 vssd1 vssd1 vccd1 vccd1 net1255 sky130_fd_sc_hd__clkbuf_4
X_17782_ net842 net990 net825 net974 net969 vssd1 vssd1 vccd1 vccd1 _03460_ sky130_fd_sc_hd__a41o_1
XFILLER_0_98_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1266 net1267 vssd1 vssd1 vccd1 vccd1 net1266 sky130_fd_sc_hd__clkbuf_2
X_14994_ control.body\[1000\] net152 _01551_ net2451 vssd1 vssd1 vccd1 vccd1 _00330_
+ sky130_fd_sc_hd__a22o_1
Xfanout1277 net1280 vssd1 vssd1 vccd1 vccd1 net1277 sky130_fd_sc_hd__clkbuf_4
Xfanout1288 net1291 vssd1 vssd1 vccd1 vccd1 net1288 sky130_fd_sc_hd__clkbuf_4
Xfanout290 net294 vssd1 vssd1 vccd1 vccd1 net290 sky130_fd_sc_hd__clkbuf_4
Xfanout1299 net1310 vssd1 vssd1 vccd1 vccd1 net1299 sky130_fd_sc_hd__clkbuf_2
XANTENNA__18034__B1 net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16733_ obsg2.obstacleArray\[103\] net500 net481 obsg2.obstacleArray\[101\] vssd1
+ vssd1 vccd1 vccd1 _02412_ sky130_fd_sc_hd__a22o_1
X_19521_ clknet_leaf_121_clk net2530 net1402 vssd1 vssd1 vccd1 vccd1 control.body\[879\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13283__Y _07827_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13945_ ag2.body\[87\] net197 _08154_ ag2.body\[79\] vssd1 vssd1 vccd1 vccd1 _00168_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__10254__A_N net1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17388__A2 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkload6_A clknet_4_12__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19452_ clknet_leaf_109_clk _00396_ net1420 vssd1 vssd1 vccd1 vccd1 control.body\[938\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_134_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16664_ obsg2.obstacleArray\[22\] net448 vssd1 vssd1 vccd1 vccd1 _02343_ sky130_fd_sc_hd__or2_1
XANTENNA__16596__B1 net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13876_ ag2.body\[25\] net121 _08147_ ag2.body\[17\] vssd1 vssd1 vccd1 vccd1 _00106_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_88_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_1162 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15615_ ag2.body\[448\] net123 _01613_ ag2.body\[440\] vssd1 vssd1 vccd1 vccd1 _00882_
+ sky130_fd_sc_hd__a22o_1
X_18403_ _04493_ _04639_ _03831_ _03892_ vssd1 vssd1 vccd1 vccd1 _03893_ sky130_fd_sc_hd__o211a_1
XANTENNA__11244__B net1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12827_ net288 _07613_ _07614_ net1873 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[170\]
+ sky130_fd_sc_hd__a22o_1
X_19383_ clknet_leaf_93_clk _00327_ net1436 vssd1 vssd1 vccd1 vccd1 control.body\[1013\]
+ sky130_fd_sc_hd__dfrtp_1
X_16595_ obsg2.obstacleArray\[78\] net443 vssd1 vssd1 vccd1 vccd1 _02274_ sky130_fd_sc_hd__or2_1
XANTENNA__14071__A1 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14071__B2 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18334_ _03822_ _03829_ vssd1 vssd1 vccd1 vccd1 _03830_ sky130_fd_sc_hd__nand2_1
XFILLER_0_70_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15546_ ag2.body\[516\] net184 _01580_ ag2.body\[508\] vssd1 vssd1 vccd1 vccd1 _00822_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12082__B1 net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12758_ net237 _07582_ _07583_ net1743 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[132\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_45_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_96_3236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18265_ obsg2.obstacleArray\[129\] _03771_ net530 vssd1 vssd1 vccd1 vccd1 _01380_
+ sky130_fd_sc_hd__o21a_1
X_11709_ _06678_ _06680_ net565 vssd1 vssd1 vccd1 vccd1 _06681_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_96_3247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15477_ ag2.body\[582\] net111 _01604_ net1584 vssd1 vssd1 vccd1 vccd1 _00760_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_96_3258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19200__Q ag2.body\[63\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12689_ net238 _07549_ _07550_ net2036 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[96\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_115_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17216_ _02885_ _02886_ _02887_ _02888_ vssd1 vssd1 vccd1 vccd1 _02895_ sky130_fd_sc_hd__a22o_1
XFILLER_0_53_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14428_ net988 _04203_ _04204_ net971 _08588_ vssd1 vssd1 vccd1 vccd1 _08589_ sky130_fd_sc_hd__a221o_1
X_18196_ _03640_ _03703_ obsg2.obstacleArray\[95\] vssd1 vssd1 vccd1 vccd1 _03737_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_112_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11188__A2 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17147_ ag2.body\[613\] net946 vssd1 vssd1 vccd1 vccd1 _02826_ sky130_fd_sc_hd__or2_1
X_14359_ _08510_ _08511_ _08513_ _08514_ vssd1 vssd1 vccd1 vccd1 _08520_ sky130_fd_sc_hd__a22o_1
XANTENNA__16262__S net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold705 control.body\[791\] vssd1 vssd1 vccd1 vccd1 net2267 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__18043__A net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold716 control.body\[1026\] vssd1 vssd1 vccd1 vccd1 net2278 sky130_fd_sc_hd__dlygate4sd3_1
Xhold727 control.body\[634\] vssd1 vssd1 vccd1 vccd1 net2289 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10935__A2 _05890_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19180__CLK clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_1623 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold738 control.body\[941\] vssd1 vssd1 vccd1 vccd1 net2300 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09665__A _04425_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17078_ ag2.body\[193\] net731 net849 _04061_ _02756_ vssd1 vssd1 vccd1 vccd1 _02757_
+ sky130_fd_sc_hd__a221o_1
Xhold749 control.body\[865\] vssd1 vssd1 vccd1 vccd1 net2311 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_126_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16029_ net958 net538 vssd1 vssd1 vccd1 vccd1 _01708_ sky130_fd_sc_hd__and2_2
XFILLER_0_99_1409 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12091__A net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10604__A net1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20591__1523 vssd1 vssd1 vccd1 vccd1 _20591__1523/HI net1523 sky130_fd_sc_hd__conb_1
XFILLER_0_42_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10323__B net1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16284__C1 _01911_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18898__CLK clknet_leaf_144_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19719_ clknet_leaf_134_clk net2522 net1303 vssd1 vssd1 vccd1 vccd1 control.body\[677\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_81_2804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_2350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_1020 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_2203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16945__B net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09403_ net1603 _04342_ _04385_ vssd1 vssd1 vccd1 vccd1 _01401_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_48_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_62_2214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11154__B net1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_2225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14746__A net1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18328__A1 net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1087_A net1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09334_ _04335_ _04340_ vssd1 vssd1 vccd1 vccd1 _01429_ sky130_fd_sc_hd__nor2_1
XANTENNA__10993__B net1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09265_ _04288_ vssd1 vssd1 vccd1 vccd1 sound_gen.osc1.timer_nxt\[14\] sky130_fd_sc_hd__inv_2
XFILLER_0_5_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11820__B1 net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout512_A net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_2722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout133_X net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_2733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1254_A net1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_79_2744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09196_ ag2.body\[615\] vssd1 vssd1 vccd1 vccd1 _04221_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_75_2608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_2619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11179__A2 _06135_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20425_ clknet_leaf_37_clk _01312_ net1353 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[61\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_133_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout300_X net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_2018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1042_X net1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16172__S net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_56_2029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17303__A2 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20500__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20356_ clknet_leaf_18_clk _01247_ net1323 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleCount\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA_fanout881_A net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout979_A net980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20287_ clknet_leaf_35_clk control.divider.next_count\[8\] net1348 vssd1 vssd1 vccd1
+ vccd1 control.divider.count\[8\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_120_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10040_ net1107 control.body\[901\] vssd1 vssd1 vccd1 vccd1 _05013_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_8_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold10 obsmode.sOBSMODE.pb_1 vssd1 vssd1 vccd1 vccd1 net1572 sky130_fd_sc_hd__dlygate4sd3_1
Xhold21 img_gen.control.button5.Q\[1\] vssd1 vssd1 vccd1 vccd1 net1583 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout767_X net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16275__C1 net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold32 img_gen.tracker.frame\[423\] vssd1 vssd1 vccd1 vccd1 net1594 sky130_fd_sc_hd__dlygate4sd3_1
Xhold43 img_gen.tracker.frame\[403\] vssd1 vssd1 vccd1 vccd1 net1605 sky130_fd_sc_hd__dlygate4sd3_1
Xhold54 img_gen.tracker.frame\[193\] vssd1 vssd1 vccd1 vccd1 net1616 sky130_fd_sc_hd__dlygate4sd3_1
Xhold65 img_gen.tracker.frame\[265\] vssd1 vssd1 vccd1 vccd1 net1627 sky130_fd_sc_hd__dlygate4sd3_1
Xhold76 img_gen.tracker.frame\[194\] vssd1 vssd1 vccd1 vccd1 net1638 sky130_fd_sc_hd__dlygate4sd3_1
Xhold87 control.divider.fsm.current_mode\[1\] vssd1 vssd1 vccd1 vccd1 net1649 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11639__B1 _06610_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17016__B net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout934_X net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold98 img_gen.tracker.frame\[176\] vssd1 vssd1 vccd1 vccd1 net1660 sky130_fd_sc_hd__dlygate4sd3_1
X_11991_ img_gen.tracker.frame\[388\] net601 net584 img_gen.tracker.frame\[394\] _06962_
+ vssd1 vssd1 vccd1 vccd1 _06963_ sky130_fd_sc_hd__o221a_1
XANTENNA__11103__A2 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_1613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13730_ _04390_ _07218_ _07251_ _07259_ vssd1 vssd1 vccd1 vccd1 _00053_ sky130_fd_sc_hd__a22o_1
X_10942_ ag2.body\[298\] net1187 vssd1 vssd1 vccd1 vccd1 _05915_ sky130_fd_sc_hd__xor2_1
XANTENNA_fanout46_X net46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16855__B net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11064__B net1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13661_ net825 _08013_ vssd1 vssd1 vccd1 vccd1 _08015_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_45_1700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16347__S net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10873_ ag2.body\[529\] net1203 vssd1 vssd1 vccd1 vccd1 _05846_ sky130_fd_sc_hd__or2_1
X_15400_ control.body\[641\] net80 _01581_ net2416 vssd1 vssd1 vccd1 vccd1 _00691_
+ sky130_fd_sc_hd__a22o_1
X_12612_ net277 _07506_ _07507_ net1620 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[62\]
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_26_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16380_ _01900_ _02058_ vssd1 vssd1 vccd1 vccd1 _02059_ sky130_fd_sc_hd__and2_4
XANTENNA__11999__B net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13592_ control.divider.count\[10\] _07954_ _07965_ _07966_ vssd1 vssd1 vccd1 vccd1
+ _07967_ sky130_fd_sc_hd__o22a_1
XFILLER_0_17_1392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15331_ control.body\[707\] net73 _01587_ net2400 vssd1 vssd1 vccd1 vccd1 _00629_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__17967__A net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10614__B2 _05586_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12543_ net2013 net653 _07469_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[31\]
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_22_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18050_ net43 _03649_ vssd1 vssd1 vccd1 vccd1 _03650_ sky130_fd_sc_hd__nor2_1
XANTENNA__12607__C net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15262_ _04416_ net58 vssd1 vssd1 vccd1 vccd1 _01580_ sky130_fd_sc_hd__nor2_2
X_12474_ _07426_ _07427_ vssd1 vssd1 vccd1 vccd1 _07429_ sky130_fd_sc_hd__nand2b_1
XANTENNA__16750__B1 net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_3100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17001_ ag2.body\[136\] net741 net708 ag2.body\[141\] _02679_ vssd1 vssd1 vccd1 vccd1
+ _02680_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_91_3111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18134__Y _03705_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_91_clk_A clknet_4_11__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14213_ net982 ag2.body\[410\] vssd1 vssd1 vccd1 vccd1 _08374_ sky130_fd_sc_hd__xor2_1
XFILLER_0_65_1622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11425_ _06371_ _06384_ _06390_ _06397_ vssd1 vssd1 vccd1 vccd1 _06398_ sky130_fd_sc_hd__o22a_1
XFILLER_0_62_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15193_ control.body\[825\] net94 _01573_ net2494 vssd1 vssd1 vccd1 vccd1 _00507_
+ sky130_fd_sc_hd__a22o_1
XANTENNA_7 _03442_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_20_Left_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_1515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_1526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14144_ _08293_ _08294_ _08303_ _08304_ vssd1 vssd1 vccd1 vccd1 _08305_ sky130_fd_sc_hd__a211o_1
XFILLER_0_10_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13278__Y _07825_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11356_ net1201 control.body\[809\] vssd1 vssd1 vccd1 vccd1 _06329_ sky130_fd_sc_hd__or2_1
XANTENNA__12119__A1 net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10307_ net1072 control.body\[702\] vssd1 vssd1 vccd1 vccd1 _05280_ sky130_fd_sc_hd__or2_1
XANTENNA__18013__D net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14075_ _08230_ _08233_ _08234_ _08235_ vssd1 vssd1 vccd1 vccd1 _08236_ sky130_fd_sc_hd__or4b_1
X_18952_ clknet_leaf_5_clk img_gen.tracker.next_frame\[390\] net1276 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[390\] sky130_fd_sc_hd__dfrtp_1
X_11287_ net1232 control.body\[1104\] vssd1 vssd1 vccd1 vccd1 _06260_ sky130_fd_sc_hd__xor2_1
X_17903_ net432 _02054_ vssd1 vssd1 vccd1 vccd1 _03538_ sky130_fd_sc_hd__and2_1
X_13026_ net385 _07535_ _07638_ vssd1 vssd1 vccd1 vccd1 _07708_ sky130_fd_sc_hd__and3_1
X_10238_ ag2.body\[325\] net1116 vssd1 vssd1 vccd1 vccd1 _05211_ sky130_fd_sc_hd__xor2_4
XTAP_TAPCELL_ROW_89_3040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11239__B net1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_3051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18883_ clknet_leaf_12_clk img_gen.tracker.next_frame\[321\] net1283 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[321\] sky130_fd_sc_hd__dfrtp_1
Xfanout1030 net1031 vssd1 vssd1 vccd1 vccd1 net1030 sky130_fd_sc_hd__buf_4
XANTENNA__16266__C1 net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15608__A2 net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1041 net1042 vssd1 vssd1 vccd1 vccd1 net1041 sky130_fd_sc_hd__buf_2
XFILLER_0_101_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09932__B net1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17834_ net1034 ag2.apple_cord\[4\] net224 vssd1 vssd1 vccd1 vccd1 _03494_ sky130_fd_sc_hd__mux2_1
Xfanout1052 net1053 vssd1 vssd1 vccd1 vccd1 net1052 sky130_fd_sc_hd__buf_4
X_10169_ _05137_ _05139_ _05140_ _05141_ vssd1 vssd1 vccd1 vccd1 _05142_ sky130_fd_sc_hd__or4_1
XFILLER_0_83_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1063 net1069 vssd1 vssd1 vccd1 vccd1 net1063 sky130_fd_sc_hd__buf_2
XFILLER_0_94_1328 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1074 net1082 vssd1 vssd1 vccd1 vccd1 net1074 sky130_fd_sc_hd__buf_4
Xfanout1085 net1093 vssd1 vssd1 vccd1 vccd1 net1085 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_59_1459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1096 net1098 vssd1 vssd1 vccd1 vccd1 net1096 sky130_fd_sc_hd__clkbuf_4
X_14977_ control.body\[1016\] net158 _01550_ control.body\[1008\] vssd1 vssd1 vccd1
+ vccd1 _00314_ sky130_fd_sc_hd__a22o_1
X_17765_ _02807_ _02810_ _02815_ _03218_ vssd1 vssd1 vccd1 vccd1 _03444_ sky130_fd_sc_hd__o31a_2
XFILLER_0_107_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19504_ clknet_leaf_113_clk _00448_ net1401 vssd1 vssd1 vccd1 vccd1 control.body\[894\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11255__A net1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16716_ obsg2.obstacleArray\[123\] net501 net487 obsg2.obstacleArray\[122\] vssd1
+ vssd1 vccd1 vccd1 _02395_ sky130_fd_sc_hd__a22o_1
X_13928_ _04863_ net61 vssd1 vssd1 vccd1 vccd1 _08153_ sky130_fd_sc_hd__nor2_2
XFILLER_0_88_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17696_ _04044_ net877 net713 ag2.body\[156\] _03374_ vssd1 vssd1 vccd1 vccd1 _03375_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_117_1048 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1052 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16647_ obsg2.obstacleArray\[2\] obsg2.obstacleArray\[3\] net446 vssd1 vssd1 vccd1
+ vccd1 _02326_ sky130_fd_sc_hd__mux2_1
X_19435_ clknet_leaf_108_clk net2520 net1421 vssd1 vssd1 vccd1 vccd1 control.body\[953\]
+ sky130_fd_sc_hd__dfrtp_1
X_13859_ ag2.body\[22\] net116 _08134_ ag2.body\[14\] vssd1 vssd1 vccd1 vccd1 _00102_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_18_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_44_clk_A clknet_4_7__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_3309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18038__A _03543_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15241__B1 _01578_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13470__A _07592_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12055__B1 net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16578_ obsg2.obstacleArray\[114\] net443 vssd1 vssd1 vccd1 vccd1 _02257_ sky130_fd_sc_hd__or2_1
XANTENNA__19546__CLK clknet_leaf_115_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19366_ clknet_leaf_102_clk _00310_ net1438 vssd1 vssd1 vccd1 vccd1 control.body\[1028\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__19231__RESET_B net1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15792__B2 ag2.body\[294\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18317_ _03786_ _03790_ _08053_ vssd1 vssd1 vccd1 vccd1 _03813_ sky130_fd_sc_hd__o21ai_1
X_15529_ ag2.body\[532\] net158 _01610_ ag2.body\[524\] vssd1 vssd1 vccd1 vccd1 _00806_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11802__B1 net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19297_ clknet_leaf_99_clk net2200 net1447 vssd1 vssd1 vccd1 vccd1 control.body\[1103\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__17533__A2 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09050_ ag2.body\[240\] vssd1 vssd1 vccd1 vccd1 _04075_ sky130_fd_sc_hd__inv_2
X_18248_ _03689_ net35 vssd1 vssd1 vccd1 vccd1 _03763_ sky130_fd_sc_hd__nor2_1
XANTENNA__20523__CLK clknet_leaf_93_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_59_clk_A clknet_4_13__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16741__B1 net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10318__B net1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18179_ obsg2.obstacleArray\[86\] _03728_ net532 vssd1 vssd1 vccd1 vccd1 _01337_
+ sky130_fd_sc_hd__o21a_1
XANTENNA_clkbuf_leaf_102_clk_A clknet_4_10__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold502 img_gen.tracker.frame\[48\] vssd1 vssd1 vccd1 vccd1 net2064 sky130_fd_sc_hd__dlygate4sd3_1
X_20210_ clknet_leaf_60_clk _01154_ net1466 vssd1 vssd1 vccd1 vccd1 ag2.body\[176\]
+ sky130_fd_sc_hd__dfrtp_4
Xhold513 img_gen.tracker.frame\[249\] vssd1 vssd1 vccd1 vccd1 net2075 sky130_fd_sc_hd__dlygate4sd3_1
Xhold524 img_gen.tracker.frame\[568\] vssd1 vssd1 vccd1 vccd1 net2086 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold535 img_gen.tracker.frame\[54\] vssd1 vssd1 vccd1 vccd1 net2097 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold546 img_gen.tracker.frame\[570\] vssd1 vssd1 vccd1 vccd1 net2108 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__16005__B net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold557 img_gen.tracker.frame\[243\] vssd1 vssd1 vccd1 vccd1 net2119 sky130_fd_sc_hd__dlygate4sd3_1
Xhold568 img_gen.updater.commands.rR1.rainbowRNG\[15\] vssd1 vssd1 vccd1 vccd1 net2130
+ sky130_fd_sc_hd__dlygate4sd3_1
X_20141_ clknet_leaf_97_clk _01085_ net1449 vssd1 vssd1 vccd1 vccd1 ag2.body\[251\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_64_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09952_ control.body\[740\] net1119 vssd1 vssd1 vccd1 vccd1 _04925_ sky130_fd_sc_hd__nand2b_1
Xhold579 control.body\[1047\] vssd1 vssd1 vccd1 vccd1 net2141 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09682__X _04655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20072_ clknet_leaf_73_clk _01016_ net1500 vssd1 vssd1 vccd1 vccd1 ag2.body\[326\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA_clkbuf_leaf_117_clk_A clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11869__B1 net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09883_ ag2.body\[160\] net784 net1209 _04050_ _04850_ vssd1 vssd1 vccd1 vccd1 _04856_
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_42_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16257__C1 net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18220__B net40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout295_A _07335_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_2401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1002_A net1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_2412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14283__A1 net1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout462_A net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14283__B2 net1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15480__B1 _01605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17757__C1 net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16675__B net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout250_X net250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14476__A net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout348_X net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout727_A net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1469_A net1470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12046__B1 net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16980__B1 net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12597__A1 net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09317_ _04323_ _04332_ sound_gen.osc1.count\[3\] net272 vssd1 vssd1 vccd1 vccd1
+ _01438_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA_fanout515_X net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14763__X _08924_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17524__A2 net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_1644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09857__X _04830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09248_ img_gen.updater.commands.cmd_num\[0\] vssd1 vssd1 vccd1 vccd1 _04273_ sky130_fd_sc_hd__inv_2
XFILLER_0_105_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16732__B1 net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10228__B net1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09179_ ag2.body\[555\] vssd1 vssd1 vccd1 vccd1 _04204_ sky130_fd_sc_hd__inv_2
X_11210_ net1051 control.body\[847\] vssd1 vssd1 vccd1 vccd1 _06183_ sky130_fd_sc_hd__xnor2_1
X_20408_ clknet_leaf_31_clk _01295_ net1338 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[44\]
+ sky130_fd_sc_hd__dfrtp_2
X_12190_ net1222 ag2.apple_cord\[0\] vssd1 vssd1 vccd1 vccd1 _07162_ sky130_fd_sc_hd__or2_1
XFILLER_0_82_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13539__B net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout884_X net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09935__A_N net1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput11 net11 vssd1 vssd1 vccd1 vccd1 gpio_out[10] sky130_fd_sc_hd__buf_2
XFILLER_0_124_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput22 net22 vssd1 vssd1 vccd1 vccd1 gpio_out[20] sky130_fd_sc_hd__buf_2
X_11141_ ag2.body\[408\] net1234 vssd1 vssd1 vccd1 vccd1 _06114_ sky130_fd_sc_hd__xor2_1
Xoutput33 net33 vssd1 vssd1 vccd1 vccd1 gpio_out[8] sky130_fd_sc_hd__buf_2
X_20339_ clknet_leaf_20_clk _01230_ net1364 vssd1 vssd1 vccd1 vccd1 ag2.apple_cord\[7\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_120_1406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17953__C _03579_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13849__B2 net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11059__B net1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11072_ ag2.body\[367\] net747 net772 ag2.body\[363\] vssd1 vssd1 vccd1 vccd1 _06045_
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_21_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10023_ _04991_ _04993_ _04995_ vssd1 vssd1 vccd1 vccd1 _04996_ sky130_fd_sc_hd__or3_4
XANTENNA__11774__S net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14900_ control.body\[1093\] net177 _01540_ net2253 vssd1 vssd1 vccd1 vccd1 _00247_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__09752__B net1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15880_ ag2.body\[221\] net192 _01648_ ag2.body\[213\] vssd1 vssd1 vccd1 vccd1 _01119_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_95_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14831_ _08327_ _08333_ _01500_ _01501_ _08268_ vssd1 vssd1 vccd1 vccd1 _01502_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_118_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14274__A1 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_1335 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14274__B2 net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17550_ _03224_ _03225_ _03226_ _03228_ vssd1 vssd1 vccd1 vccd1 _03229_ sky130_fd_sc_hd__a211o_1
XFILLER_0_54_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14762_ net840 ag2.body\[40\] _08922_ vssd1 vssd1 vccd1 vccd1 _08923_ sky130_fd_sc_hd__o21a_1
XFILLER_0_99_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11974_ img_gen.tracker.frame\[571\] net550 vssd1 vssd1 vccd1 vccd1 _06946_ sky130_fd_sc_hd__or2_1
XANTENNA__09820__A1_N net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16501_ net367 _02177_ _02179_ vssd1 vssd1 vccd1 vccd1 _02180_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_98_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16585__B net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_486 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13713_ net326 vssd1 vssd1 vccd1 vccd1 _08051_ sky130_fd_sc_hd__inv_2
X_17481_ ag2.body\[128\] net887 vssd1 vssd1 vccd1 vccd1 _03160_ sky130_fd_sc_hd__or2_1
X_10925_ net1231 control.body\[1032\] vssd1 vssd1 vccd1 vccd1 _05898_ sky130_fd_sc_hd__xor2_1
X_14693_ net993 _04110_ _04112_ net1012 _08853_ vssd1 vssd1 vccd1 vccd1 _08854_ sky130_fd_sc_hd__a221o_1
XANTENNA__16077__S net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14026__A1 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14026__B2 net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1498 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19220_ clknet_leaf_75_clk _00164_ net1494 vssd1 vssd1 vccd1 vccd1 ag2.body\[83\]
+ sky130_fd_sc_hd__dfrtp_4
X_16432_ obsg2.obstacleArray\[78\] net453 vssd1 vssd1 vccd1 vccd1 _02111_ sky130_fd_sc_hd__or2_1
X_13644_ control.divider.count\[15\] _08002_ vssd1 vssd1 vccd1 vccd1 _08004_ sky130_fd_sc_hd__and2_1
XANTENNA__20546__CLK clknet_leaf_105_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12037__B1 net557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10856_ net1218 control.body\[688\] vssd1 vssd1 vccd1 vccd1 _05829_ sky130_fd_sc_hd__xor2_1
XFILLER_0_85_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19151_ clknet_leaf_51_clk _00095_ net1367 vssd1 vssd1 vccd1 vccd1 ag2.body\[15\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__18593__CLK clknet_leaf_13_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20590__1522 vssd1 vssd1 vccd1 vccd1 _20590__1522/HI net1522 sky130_fd_sc_hd__conb_1
X_16363_ net420 _02039_ _02041_ net370 vssd1 vssd1 vccd1 vccd1 _02042_ sky130_fd_sc_hd__a211o_1
XFILLER_0_32_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13575_ control.divider.fsm.current_mode\[2\] _03961_ vssd1 vssd1 vccd1 vccd1 _07950_
+ sky130_fd_sc_hd__nor2_1
XANTENNA__10419__A net1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10787_ net1219 control.body\[624\] vssd1 vssd1 vccd1 vccd1 _05760_ sky130_fd_sc_hd__xor2_1
X_18102_ net44 _03683_ vssd1 vssd1 vccd1 vccd1 _03684_ sky130_fd_sc_hd__nor2_1
XANTENNA__11796__C1 net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17515__A2 net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15314_ control.body\[723\] net74 _01588_ control.body\[715\] vssd1 vssd1 vccd1 vccd1
+ _00613_ sky130_fd_sc_hd__a22o_1
XFILLER_0_82_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11260__A1 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10063__A2 _04519_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12526_ net629 net437 net473 net561 vssd1 vssd1 vccd1 vccd1 _07460_ sky130_fd_sc_hd__and4_2
XANTENNA__09767__X _04740_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19082_ clknet_leaf_29_clk img_gen.tracker.next_frame\[520\] net1334 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[520\] sky130_fd_sc_hd__dfrtp_1
X_16294_ _01971_ _01972_ net419 vssd1 vssd1 vccd1 vccd1 _01973_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15929__B net57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18033_ net351 net38 _03638_ vssd1 vssd1 vccd1 vccd1 _03639_ sky130_fd_sc_hd__and3_1
XFILLER_0_124_444 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15245_ _06138_ net53 vssd1 vssd1 vccd1 vccd1 _01579_ sky130_fd_sc_hd__nor2_2
X_12457_ img_gen.updater.commands.rR1.rainbowRNG\[15\] _07319_ _07320_ _07409_ _07416_
+ vssd1 vssd1 vccd1 vccd1 _07417_ sky130_fd_sc_hd__a221o_1
XFILLER_0_78_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12634__A net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11408_ ag2.body\[572\] net1132 vssd1 vssd1 vccd1 vccd1 _06381_ sky130_fd_sc_hd__xor2_1
X_15176_ net2610 net102 _01571_ control.body\[834\] vssd1 vssd1 vccd1 vccd1 _00492_
+ sky130_fd_sc_hd__a22o_1
X_12388_ _07299_ _07351_ net1122 vssd1 vssd1 vccd1 vccd1 _07353_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16487__C1 net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12760__A1 net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14127_ _08285_ _08286_ _08287_ _08284_ vssd1 vssd1 vccd1 vccd1 _08288_ sky130_fd_sc_hd__a211o_1
XFILLER_0_61_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_1030 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11339_ _06306_ _06308_ _06310_ _06311_ vssd1 vssd1 vccd1 vccd1 _06312_ sky130_fd_sc_hd__or4_2
X_19984_ clknet_leaf_64_clk _00928_ net1474 vssd1 vssd1 vccd1 vccd1 ag2.body\[414\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__11581__C_N _06497_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10154__A ag2.body\[59\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13168__C _07508_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09508__A2 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19099__CLK clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18935_ clknet_leaf_139_clk img_gen.tracker.next_frame\[373\] net1288 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[373\] sky130_fd_sc_hd__dfrtp_1
X_14058_ net996 ag2.body\[32\] vssd1 vssd1 vccd1 vccd1 _08219_ sky130_fd_sc_hd__xor2_1
XANTENNA__18040__B net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13009_ net668 _07699_ vssd1 vssd1 vccd1 vccd1 _07700_ sky130_fd_sc_hd__nor2_1
XANTENNA__09662__B net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1212 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18866_ clknet_leaf_12_clk img_gen.tracker.next_frame\[304\] net1285 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[304\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_118_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17817_ _03482_ _03483_ vssd1 vssd1 vccd1 vccd1 _03484_ sky130_fd_sc_hd__nor2_1
XANTENNA__10160__Y _05133_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14848__X _01519_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18797_ clknet_leaf_12_clk img_gen.tracker.next_frame\[235\] net1285 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[235\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__15462__B1 _01603_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17748_ _02626_ _02629_ _02631_ _03098_ vssd1 vssd1 vccd1 vccd1 _03427_ sky130_fd_sc_hd__o31a_1
XANTENNA__17739__C1 _03415_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14017__A1 net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14017__B2 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17679_ ag2.body\[474\] net725 net929 _04172_ vssd1 vssd1 vccd1 vccd1 _03358_ sky130_fd_sc_hd__a22o_1
XFILLER_0_33_1418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16411__C1 net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19418_ clknet_leaf_111_clk _00362_ net1427 vssd1 vssd1 vccd1 vccd1 control.body\[968\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_130_1023 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_704 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12579__A1 net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11432__B net1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19349_ clknet_leaf_101_clk _00293_ net1444 vssd1 vssd1 vccd1 vccd1 control.body\[1043\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_116_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17506__A2 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09102_ ag2.body\[355\] vssd1 vssd1 vccd1 vccd1 _04127_ sky130_fd_sc_hd__inv_2
XFILLER_0_2_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16714__B1 net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09033_ ag2.body\[182\] vssd1 vssd1 vccd1 vccd1 _04058_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout210_A net218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12544__A net225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout308_A net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11003__A1 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18467__B1 net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold310 img_gen.tracker.frame\[548\] vssd1 vssd1 vccd1 vccd1 net1872 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11003__B2 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold321 img_gen.tracker.frame\[266\] vssd1 vssd1 vccd1 vccd1 net1883 sky130_fd_sc_hd__dlygate4sd3_1
Xhold332 img_gen.tracker.frame\[450\] vssd1 vssd1 vccd1 vccd1 net1894 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold343 img_gen.tracker.frame\[322\] vssd1 vssd1 vccd1 vccd1 net1905 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold354 img_gen.tracker.frame\[167\] vssd1 vssd1 vccd1 vccd1 net1916 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10064__A net1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold365 img_gen.tracker.frame\[432\] vssd1 vssd1 vccd1 vccd1 net1927 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold376 img_gen.tracker.frame\[245\] vssd1 vssd1 vccd1 vccd1 net1938 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__16885__A2_N net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1217_A net1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold387 img_gen.tracker.frame\[318\] vssd1 vssd1 vccd1 vccd1 net1949 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout801 net805 vssd1 vssd1 vccd1 vccd1 net801 sky130_fd_sc_hd__clkbuf_2
XANTENNA__18219__B1 net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20124_ clknet_leaf_79_clk _01068_ net1486 vssd1 vssd1 vccd1 vccd1 ag2.body\[266\]
+ sky130_fd_sc_hd__dfrtp_4
Xhold398 img_gen.tracker.frame\[513\] vssd1 vssd1 vccd1 vccd1 net1960 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09853__A net1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout812 net813 vssd1 vssd1 vccd1 vccd1 net812 sky130_fd_sc_hd__buf_4
X_09935_ net1198 ag2.body\[25\] vssd1 vssd1 vccd1 vccd1 _04908_ sky130_fd_sc_hd__and2b_1
Xfanout823 _03968_ vssd1 vssd1 vccd1 vccd1 net823 sky130_fd_sc_hd__buf_2
Xfanout834 net835 vssd1 vssd1 vccd1 vccd1 net834 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout677_A net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout845 net846 vssd1 vssd1 vccd1 vccd1 net845 sky130_fd_sc_hd__buf_4
XANTENNA_fanout298_X net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout856 net857 vssd1 vssd1 vccd1 vccd1 net856 sky130_fd_sc_hd__buf_4
X_20055_ clknet_leaf_73_clk _00999_ net1502 vssd1 vssd1 vccd1 vccd1 ag2.body\[341\]
+ sky130_fd_sc_hd__dfrtp_4
Xfanout867 obsg2.randCord\[2\] vssd1 vssd1 vccd1 vccd1 net867 sky130_fd_sc_hd__clkbuf_8
X_09866_ _04835_ _04836_ _04837_ _04838_ vssd1 vssd1 vccd1 vccd1 _04839_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout1005_X net1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout878 obsg2.randCord\[1\] vssd1 vssd1 vccd1 vccd1 net878 sky130_fd_sc_hd__clkbuf_4
Xhold1010 control.body\[662\] vssd1 vssd1 vccd1 vccd1 net2572 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1021 control.body\[642\] vssd1 vssd1 vccd1 vccd1 net2583 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout889 obsg2.randCord\[0\] vssd1 vssd1 vccd1 vccd1 net889 sky130_fd_sc_hd__buf_6
XFILLER_0_77_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1032 control.body\[777\] vssd1 vssd1 vccd1 vccd1 net2594 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13094__B _07460_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1043 control.body\[1069\] vssd1 vssd1 vccd1 vccd1 net2605 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14256__A1 net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout844_A net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09797_ net1060 control.body\[967\] vssd1 vssd1 vccd1 vccd1 _04770_ sky130_fd_sc_hd__xor2_1
Xhold1054 control.body\[703\] vssd1 vssd1 vccd1 vccd1 net2616 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14256__B2 net1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1065 control.body\[792\] vssd1 vssd1 vccd1 vccd1 net2627 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout465_X net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15453__B1 _01602_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1076 control.body\[633\] vssd1 vssd1 vccd1 vccd1 net2638 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1087 control.body\[1050\] vssd1 vssd1 vccd1 vccd1 net2649 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14812__A1_N net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1098 control.body\[901\] vssd1 vssd1 vccd1 vccd1 net2660 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__16973__X _02652_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout632_X net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1374_X net1374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14008__B2 net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15205__B1 _01574_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11045__D _06017_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10710_ _05679_ _05680_ _05681_ _05682_ vssd1 vssd1 vccd1 vccd1 _05683_ sky130_fd_sc_hd__or4_1
XANTENNA__12019__B1 net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11690_ img_gen.tracker.frame\[101\] net602 vssd1 vssd1 vccd1 vccd1 _06662_ sky130_fd_sc_hd__or2_1
XANTENNA__11342__B net1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10641_ net1168 control.body\[666\] vssd1 vssd1 vccd1 vccd1 _05614_ sky130_fd_sc_hd__xor2_1
XANTENNA__14493__X _08654_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_843 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_271 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13360_ net249 _07856_ _07857_ net1962 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[460\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__15749__B net60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10572_ ag2.body\[189\] net1104 vssd1 vssd1 vccd1 vccd1 _05545_ sky130_fd_sc_hd__xor2_1
XFILLER_0_36_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11793__A2 net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12311_ _07221_ _07272_ _07218_ vssd1 vssd1 vccd1 vccd1 _07278_ sky130_fd_sc_hd__nor3b_1
XFILLER_0_23_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12990__A1 net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09747__B net1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13291_ net255 _07829_ _07830_ net1720 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[418\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_106_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15030_ _04772_ net66 vssd1 vssd1 vccd1 vccd1 _01556_ sky130_fd_sc_hd__and2_2
XFILLER_0_106_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12242_ img_gen.updater.commands.count\[8\] img_gen.updater.commands.count\[7\] _07211_
+ img_gen.updater.commands.count\[9\] img_gen.updater.commands.count\[11\] vssd1 vssd1
+ vccd1 vccd1 _07212_ sky130_fd_sc_hd__o311a_1
XFILLER_0_107_1036 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16469__C1 _02076_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12742__A1 net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16360__S net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12173_ net387 _07144_ vssd1 vssd1 vccd1 vccd1 _07145_ sky130_fd_sc_hd__or2_1
XFILLER_0_48_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17130__B1 net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16484__A2 _02059_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11124_ _06093_ _06094_ _06095_ _06096_ _06092_ vssd1 vssd1 vccd1 vccd1 _06097_ sky130_fd_sc_hd__a221o_1
X_16981_ ag2.body\[429\] net703 net696 ag2.body\[430\] _02656_ vssd1 vssd1 vccd1 vccd1
+ _02660_ sky130_fd_sc_hd__o221a_1
XFILLER_0_60_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19923__RESET_B net1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17980__A net39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18720_ clknet_leaf_142_clk img_gen.tracker.next_frame\[158\] net1258 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[158\] sky130_fd_sc_hd__dfrtp_1
X_15932_ ag2.body\[170\] net126 _01655_ ag2.body\[162\] vssd1 vssd1 vccd1 vccd1 _01164_
+ sky130_fd_sc_hd__a22o_1
X_11055_ _04427_ _04758_ net642 vssd1 vssd1 vccd1 vccd1 _06028_ sky130_fd_sc_hd__a21o_2
XANTENNA__19391__CLK clknet_leaf_102_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10006_ net911 net906 net918 net914 vssd1 vssd1 vccd1 vccd1 _04979_ sky130_fd_sc_hd__or4_2
XFILLER_0_137_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18651_ clknet_leaf_130_clk img_gen.tracker.next_frame\[89\] net1317 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[89\] sky130_fd_sc_hd__dfrtp_1
X_15863_ ag2.body\[238\] net174 _01646_ ag2.body\[230\] vssd1 vssd1 vccd1 vccd1 _01104_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_21_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14247__B2 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15444__B1 _01601_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17602_ ag2.body\[416\] net889 vssd1 vssd1 vccd1 vccd1 _03281_ sky130_fd_sc_hd__xor2_1
XFILLER_0_118_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14814_ net1018 ag2.body\[382\] vssd1 vssd1 vccd1 vccd1 _01485_ sky130_fd_sc_hd__nand2_1
XFILLER_0_99_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15794_ _04983_ net49 vssd1 vssd1 vccd1 vccd1 _01640_ sky130_fd_sc_hd__and2b_2
X_18582_ clknet_leaf_14_clk img_gen.tracker.next_frame\[20\] net1280 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[20\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10808__A1 _05670_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14745_ net985 ag2.body\[106\] vssd1 vssd1 vccd1 vccd1 _08906_ sky130_fd_sc_hd__xor2_1
X_17533_ ag2.body\[274\] net726 net933 _04095_ _03211_ vssd1 vssd1 vccd1 vccd1 _03212_
+ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_103_Left_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11957_ net469 _06917_ _06920_ _06926_ net437 vssd1 vssd1 vccd1 vccd1 _06929_ sky130_fd_sc_hd__o311a_1
XFILLER_0_131_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_120_3980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11533__A net1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_3991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10908_ net1045 control.body\[679\] vssd1 vssd1 vccd1 vccd1 _05881_ sky130_fd_sc_hd__xor2_1
X_17464_ ag2.body\[533\] net952 vssd1 vssd1 vccd1 vccd1 _03143_ sky130_fd_sc_hd__xor2_1
XFILLER_0_131_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15747__A1 ag2.body\[342\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14676_ net1028 ag2.body\[389\] vssd1 vssd1 vccd1 vccd1 _08837_ sky130_fd_sc_hd__nand2_1
XANTENNA__20410__RESET_B net1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_309 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11888_ img_gen.tracker.frame\[40\] net607 net591 img_gen.tracker.frame\[46\] vssd1
+ vssd1 vccd1 vccd1 _06860_ sky130_fd_sc_hd__o22a_1
XFILLER_0_131_1354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_101_3390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16415_ net401 _02093_ _02092_ net366 vssd1 vssd1 vccd1 vccd1 _02094_ sky130_fd_sc_hd__a211o_1
X_19203_ clknet_leaf_86_clk _00147_ net1460 vssd1 vssd1 vccd1 vccd1 ag2.body\[66\]
+ sky130_fd_sc_hd__dfrtp_4
X_13627_ control.divider.count\[9\] _07990_ net220 vssd1 vssd1 vccd1 vccd1 _07993_
+ sky130_fd_sc_hd__o21ai_1
X_17395_ _04184_ net886 net712 ag2.body\[508\] vssd1 vssd1 vccd1 vccd1 _03074_ sky130_fd_sc_hd__a22o_1
X_10839_ _05787_ _05797_ _05798_ _05811_ vssd1 vssd1 vccd1 vccd1 _05812_ sky130_fd_sc_hd__o22a_1
XANTENNA__10149__A ag2.body\[58\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11769__C1 net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_8__f_clk clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_8__leaf_clk sky130_fd_sc_hd__clkbuf_16
XANTENNA__09497__X _04470_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16346_ obsg2.obstacleArray\[90\] obsg2.obstacleArray\[91\] net411 vssd1 vssd1 vccd1
+ vccd1 _02025_ sky130_fd_sc_hd__mux2_1
XANTENNA__10036__A2 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19134_ clknet_leaf_140_clk img_gen.tracker.next_frame\[572\] net1296 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[572\] sky130_fd_sc_hd__dfrtp_1
X_13558_ _07935_ _07937_ _07939_ vssd1 vssd1 vccd1 vccd1 net17 sky130_fd_sc_hd__or3_1
XANTENNA__15659__B net57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_132_Right_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11784__A2 net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_904 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15011__Y _01553_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12509_ net1898 net649 _07450_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[16\]
+ sky130_fd_sc_hd__and3_1
X_19065_ clknet_leaf_10_clk img_gen.tracker.next_frame\[503\] net1274 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[503\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16277_ obsg2.obstacleArray\[18\] net412 vssd1 vssd1 vccd1 vccd1 _01956_ sky130_fd_sc_hd__or2_1
XFILLER_0_89_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13489_ net2002 net644 _07906_ _07907_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[539\]
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_112_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18016_ obsg2.obstacleArray\[25\] _03626_ net532 vssd1 vssd1 vccd1 vccd1 _01276_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_129_1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15228_ net2627 net98 _01577_ net2191 vssd1 vssd1 vccd1 vccd1 _00538_ sky130_fd_sc_hd__a22o_1
XFILLER_0_120_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_114_3795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_112_Left_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15159_ control.body\[859\] net98 _01569_ control.body\[851\] vssd1 vssd1 vccd1 vccd1
+ _00477_ sky130_fd_sc_hd__a22o_1
XANTENNA__16270__S net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16475__A2 _02059_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09673__A net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout108 net110 vssd1 vssd1 vccd1 vccd1 net108 sky130_fd_sc_hd__buf_2
XFILLER_0_120_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19967_ clknet_leaf_62_clk _00911_ net1470 vssd1 vssd1 vccd1 vccd1 ag2.body\[429\]
+ sky130_fd_sc_hd__dfrtp_4
Xfanout119 net120 vssd1 vssd1 vccd1 vccd1 net119 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__15683__B1 _01627_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09720_ _04685_ _04688_ _04690_ _04692_ vssd1 vssd1 vccd1 vccd1 _04693_ sky130_fd_sc_hd__or4b_2
X_18918_ clknet_leaf_142_clk img_gen.tracker.next_frame\[356\] net1258 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[356\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19898_ clknet_leaf_57_clk _00842_ net1464 vssd1 vssd1 vccd1 vccd1 ag2.body\[488\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_78_1632 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11427__B net1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09651_ net1048 control.body\[751\] vssd1 vssd1 vccd1 vccd1 _04624_ sky130_fd_sc_hd__xor2_1
XFILLER_0_78_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18849_ clknet_leaf_4_clk img_gen.tracker.next_frame\[287\] net1259 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[287\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_1042 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14238__A1 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14238__B2 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09582_ net891 net897 net901 net921 vssd1 vssd1 vccd1 vccd1 _04555_ sky130_fd_sc_hd__nand4b_2
XPHY_EDGE_ROW_121_Left_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17114__B net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout160_A net161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12539__A net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11443__A net1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout258_A net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19114__CLK clknet_leaf_141_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20151__RESET_B net1452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15738__B2 ag2.body\[342\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16953__B net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout425_A _01735_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17768__C _02768_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14754__A net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1167_A net1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09848__A net1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15569__B net61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1360 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18152__A2 _03579_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14183__A1_N net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11775__A2 net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17568__A2_N net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09567__B _04539_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1334_A net1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09016_ ag2.body\[147\] vssd1 vssd1 vccd1 vccd1 _04041_ sky130_fd_sc_hd__inv_2
XFILLER_0_104_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11527__A2 net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout794_A net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12724__A1 net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold140 img_gen.tracker.frame\[188\] vssd1 vssd1 vccd1 vccd1 net1702 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_108_1389 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16180__S net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold151 img_gen.tracker.frame\[125\] vssd1 vssd1 vccd1 vccd1 net1713 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1501_A net1502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold162 img_gen.tracker.frame\[512\] vssd1 vssd1 vccd1 vccd1 net1724 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1122_X net1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10735__B1 net1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold173 img_gen.tracker.frame\[59\] vssd1 vssd1 vccd1 vccd1 net1735 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_125_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09583__A _04238_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold184 img_gen.tracker.frame\[2\] vssd1 vssd1 vccd1 vccd1 net1746 sky130_fd_sc_hd__dlygate4sd3_1
Xhold195 img_gen.tracker.frame\[544\] vssd1 vssd1 vccd1 vccd1 net1757 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout961_A net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout582_X net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout620 net626 vssd1 vssd1 vccd1 vccd1 net620 sky130_fd_sc_hd__buf_2
XANTENNA__12721__B _07564_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout631 _06462_ vssd1 vssd1 vccd1 vccd1 net631 sky130_fd_sc_hd__buf_4
XFILLER_0_121_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09918_ _04105_ net1186 net1140 _04106_ _04890_ vssd1 vssd1 vccd1 vccd1 _04891_ sky130_fd_sc_hd__a221o_1
X_20107_ clknet_leaf_79_clk _01051_ net1487 vssd1 vssd1 vccd1 vccd1 ag2.body\[281\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_22_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout642 _04417_ vssd1 vssd1 vccd1 vccd1 net642 sky130_fd_sc_hd__buf_4
Xfanout653 net654 vssd1 vssd1 vccd1 vccd1 net653 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout664 net674 vssd1 vssd1 vccd1 vccd1 net664 sky130_fd_sc_hd__clkbuf_4
Xfanout675 net676 vssd1 vssd1 vccd1 vccd1 net675 sky130_fd_sc_hd__clkbuf_4
X_20038_ clknet_leaf_68_clk _00982_ net1494 vssd1 vssd1 vccd1 vccd1 ag2.body\[356\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_57_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout686 _04393_ vssd1 vssd1 vccd1 vccd1 net686 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_137_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout697 net698 vssd1 vssd1 vccd1 vccd1 net697 sky130_fd_sc_hd__buf_2
X_09849_ _04445_ _04607_ _04819_ _04820_ _04821_ vssd1 vssd1 vccd1 vccd1 _04822_ sky130_fd_sc_hd__a221o_1
XANTENNA__10241__B net1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout847_X net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_4091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12860_ net675 _07631_ vssd1 vssd1 vccd1 vccd1 _07632_ sky130_fd_sc_hd__nor2_1
XFILLER_0_119_1463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11811_ img_gen.tracker.frame\[458\] net614 net578 img_gen.tracker.frame\[467\] _06782_
+ vssd1 vssd1 vccd1 vccd1 _06783_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_1_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17179__B1 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12791_ net316 _07598_ vssd1 vssd1 vccd1 vccd1 _07599_ sky130_fd_sc_hd__nor2_1
XFILLER_0_138_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14530_ net983 ag2.body\[250\] vssd1 vssd1 vccd1 vccd1 _08691_ sky130_fd_sc_hd__nand2_1
X_11742_ img_gen.tracker.frame\[8\] net551 vssd1 vssd1 vccd1 vccd1 _06714_ sky130_fd_sc_hd__or2_1
XFILLER_0_7_1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16863__B net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14461_ net981 _04154_ ag2.body\[439\] net792 _08621_ vssd1 vssd1 vccd1 vccd1 _08622_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_95_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11673_ _06641_ _06644_ vssd1 vssd1 vccd1 vccd1 _06645_ sky130_fd_sc_hd__xor2_1
XFILLER_0_138_377 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14664__A net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_137_4496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16200_ obsg2.obstacleArray\[40\] obsg2.obstacleArray\[41\] net422 vssd1 vssd1 vccd1
+ vccd1 _01879_ sky130_fd_sc_hd__mux2_1
XANTENNA__10018__A2 net1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13412_ net234 _07876_ _07877_ net1651 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[492\]
+ sky130_fd_sc_hd__a22o_1
X_17180_ ag2.body\[460\] net960 vssd1 vssd1 vccd1 vccd1 _02859_ sky130_fd_sc_hd__xor2_1
XANTENNA__09758__A ag2.body\[214\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10624_ ag2.body\[48\] net1223 vssd1 vssd1 vccd1 vccd1 _05597_ sky130_fd_sc_hd__or2_1
X_14392_ net846 ag2.body\[120\] ag2.body\[126\] net803 vssd1 vssd1 vccd1 vccd1 _08553_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_119_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15479__B net54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16131_ net373 _01809_ _01808_ net346 vssd1 vssd1 vccd1 vccd1 _01810_ sky130_fd_sc_hd__a211o_1
XANTENNA__11766__A2 net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17975__A net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13343_ net664 _07850_ vssd1 vssd1 vccd1 vccd1 _07851_ sky130_fd_sc_hd__nor2_1
XFILLER_0_49_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09477__B net1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_1599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10555_ _05512_ _05524_ _05527_ _05517_ vssd1 vssd1 vccd1 vccd1 _05528_ sky130_fd_sc_hd__or4b_1
XANTENNA__12184__A net1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16062_ net497 _01726_ vssd1 vssd1 vccd1 vccd1 _01741_ sky130_fd_sc_hd__or2_1
XFILLER_0_84_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13274_ net670 _07823_ vssd1 vssd1 vccd1 vccd1 _07824_ sky130_fd_sc_hd__nor2_1
X_10486_ _04214_ net1173 net1048 _04217_ _05454_ vssd1 vssd1 vccd1 vccd1 _05459_ sky130_fd_sc_hd__o221a_1
XFILLER_0_59_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15013_ control.body\[985\] net166 _01553_ control.body\[977\] vssd1 vssd1 vccd1
+ vccd1 _00347_ sky130_fd_sc_hd__a22o_1
XFILLER_0_126_1467 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12225_ img_gen.updater.commands.count\[14\] img_gen.updater.commands.count\[15\]
+ _07194_ img_gen.updater.commands.count\[16\] vssd1 vssd1 vccd1 vccd1 _07195_ sky130_fd_sc_hd__o31a_1
XFILLER_0_121_266 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17103__B1 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12912__A net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19821_ clknet_leaf_124_clk _00765_ net1408 vssd1 vssd1 vccd1 vccd1 ag2.body\[571\]
+ sky130_fd_sc_hd__dfrtp_4
X_12156_ img_gen.tracker.frame\[468\] net614 net597 img_gen.tracker.frame\[471\] _07126_
+ vssd1 vssd1 vccd1 vccd1 _07128_ sky130_fd_sc_hd__o221a_1
XFILLER_0_75_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11107_ net779 control.body\[1097\] _06078_ _06079_ vssd1 vssd1 vccd1 vccd1 _06080_
+ sky130_fd_sc_hd__o22a_1
X_19752_ clknet_leaf_130_clk _00696_ net1317 vssd1 vssd1 vccd1 vccd1 control.body\[646\]
+ sky130_fd_sc_hd__dfrtp_1
X_16964_ ag2.body\[413\] net949 vssd1 vssd1 vccd1 vccd1 _02643_ sky130_fd_sc_hd__xor2_1
X_12087_ img_gen.tracker.frame\[300\] net630 net557 img_gen.tracker.frame\[306\] vssd1
+ vssd1 vccd1 vccd1 _07059_ sky130_fd_sc_hd__a22o_1
XFILLER_0_21_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18703_ clknet_leaf_10_clk img_gen.tracker.next_frame\[141\] net1274 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[141\] sky130_fd_sc_hd__dfrtp_1
X_15915_ ag2.body\[188\] net131 _01652_ ag2.body\[180\] vssd1 vssd1 vccd1 vccd1 _01150_
+ sky130_fd_sc_hd__a22o_1
X_11038_ net750 control.body\[1046\] _06008_ _06009_ _06010_ vssd1 vssd1 vccd1 vccd1
+ _06011_ sky130_fd_sc_hd__o2111a_1
XANTENNA__11247__B net1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1242 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19683_ clknet_leaf_117_clk _00627_ net1384 vssd1 vssd1 vccd1 vccd1 control.body\[705\]
+ sky130_fd_sc_hd__dfrtp_1
X_16895_ ag2.body\[215\] net932 vssd1 vssd1 vccd1 vccd1 _02574_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10151__B net1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09940__B net1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18634_ clknet_leaf_131_clk img_gen.tracker.next_frame\[72\] net1295 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[72\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_91_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15846_ ag2.body\[255\] net176 _01644_ ag2.body\[247\] vssd1 vssd1 vccd1 vccd1 _01089_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_99_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_103_3452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_3463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18565_ clknet_leaf_15_clk img_gen.tracker.next_frame\[3\] net1313 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[3\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_103_3474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15777_ ag2.body\[304\] net208 _01638_ ag2.body\[296\] vssd1 vssd1 vccd1 vccd1 _01026_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__19203__Q ag2.body\[66\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12989_ _07690_ net254 _07688_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[256\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_115_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17516_ ag2.body\[586\] net722 net928 _04217_ _03189_ vssd1 vssd1 vccd1 vccd1 _03195_
+ sky130_fd_sc_hd__a221o_1
X_14728_ _08885_ _08886_ _08887_ _08888_ vssd1 vssd1 vccd1 vccd1 _08889_ sky130_fd_sc_hd__or4_1
XFILLER_0_87_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11454__B2 _06426_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18496_ net1517 net1511 vssd1 vssd1 vccd1 vccd1 _00027_ sky130_fd_sc_hd__or2_1
XANTENNA__19287__CLK clknet_leaf_98_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16393__A1 net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17447_ ag2.body\[379\] net852 vssd1 vssd1 vccd1 vccd1 _03126_ sky130_fd_sc_hd__xor2_1
XFILLER_0_46_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14659_ net991 ag2.body\[521\] vssd1 vssd1 vccd1 vccd1 _08820_ sky130_fd_sc_hd__xnor2_1
XANTENNA__14574__A net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18046__A net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17590__B1 net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11206__A1 _06160_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17378_ _03020_ _03048_ _03054_ _03056_ _03039_ vssd1 vssd1 vccd1 vccd1 _03057_ sky130_fd_sc_hd__o2111a_1
XTAP_TAPCELL_ROW_116_3846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20264__CLK clknet_leaf_43_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_116_3857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12806__B net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11757__A2 net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12954__A1 net246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19117_ clknet_leaf_131_clk img_gen.tracker.next_frame\[555\] net1296 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[555\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_116_3868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16329_ net415 _02007_ _02006_ net369 vssd1 vssd1 vccd1 vccd1 _02008_ sky130_fd_sc_hd__a211o_1
XANTENNA__12094__A net1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16696__A2 net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19048_ clknet_leaf_10_clk img_gen.tracker.next_frame\[486\] net1275 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[486\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__17893__A1 _03531_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19845__RESET_B net1414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09674__Y _04647_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12822__A net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10717__B1 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_4__f_clk_A clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16013__B _01691_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_2474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_2485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_2496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15120__A2 net107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16948__B net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09703_ ag2.body\[66\] net1184 vssd1 vssd1 vccd1 vccd1 _04676_ sky130_fd_sc_hd__xor2_1
XANTENNA__13131__A1 net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11157__B net1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13682__A2 net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09634_ net892 net922 vssd1 vssd1 vccd1 vccd1 _04607_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_88_2993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10996__B net1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13372__B _07535_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09565_ net923 _04445_ _04519_ vssd1 vssd1 vccd1 vccd1 _04538_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_84_2879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout542_A net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09638__B2 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11173__A net1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09496_ _04463_ _04468_ _04430_ _04458_ vssd1 vssd1 vccd1 vccd1 _04469_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__16908__B1 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11540__S1 net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11996__A2 net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout428_X net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17581__B1 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout807_A net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1072_X net1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1451_A net1452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11460__X _06433_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13198__A1 net240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18654__CLK clknet_leaf_131_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_1268 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xwire317 _06459_ vssd1 vssd1 vccd1 vccd1 net317 sky130_fd_sc_hd__buf_2
XANTENNA__12945__A1 net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_132_4360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16136__A1 net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20587_ clknet_leaf_105_clk ag2.goodColl _00051_ vssd1 vssd1 vccd1 vccd1 sound_gen.posDetector1.N\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09810__A1 _04418_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10340_ ag2.body\[525\] net1108 vssd1 vssd1 vccd1 vccd1 _05313_ sky130_fd_sc_hd__xor2_1
XFILLER_0_61_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout797_X net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10236__B net1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10271_ ag2.body\[142\] net1088 vssd1 vssd1 vccd1 vccd1 _05244_ sky130_fd_sc_hd__xor2_1
XANTENNA_fanout1504_X net1504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12732__A net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09574__B1 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12010_ _06977_ _06979_ _06981_ net558 vssd1 vssd1 vccd1 vccd1 _06982_ sky130_fd_sc_hd__a22o_1
XANTENNA__17019__B net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout964_X net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15647__B1 _01623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1404 net1453 vssd1 vssd1 vccd1 vccd1 net1404 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11920__A2 net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1415 net1453 vssd1 vssd1 vccd1 vccd1 net1415 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_54_1960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10252__A net1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1426 net1430 vssd1 vssd1 vccd1 vccd1 net1426 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_54_1971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1437 net1442 vssd1 vssd1 vccd1 vccd1 net1437 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_54_1982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout450 net451 vssd1 vssd1 vccd1 vccd1 net450 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_22_1461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1448 net1452 vssd1 vssd1 vccd1 vccd1 net1448 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_126_4175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout461 _01710_ vssd1 vssd1 vccd1 vccd1 net461 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_50_1835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1459 net1461 vssd1 vssd1 vccd1 vccd1 net1459 sky130_fd_sc_hd__clkbuf_4
XANTENNA__16858__B net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout472 _06647_ vssd1 vssd1 vccd1 vccd1 net472 sky130_fd_sc_hd__clkbuf_4
X_13961_ ag2.body\[101\] net189 _08156_ ag2.body\[93\] vssd1 vssd1 vccd1 vccd1 _00182_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_35_1392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_4039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout483 _02373_ vssd1 vssd1 vccd1 vccd1 net483 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_6_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_1502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout494 _01736_ vssd1 vssd1 vccd1 vccd1 net494 sky130_fd_sc_hd__clkbuf_2
XANTENNA__14659__A net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_1573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_31_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17035__A ag2.body\[122\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15700_ ag2.body\[381\] net140 _01628_ ag2.body\[373\] vssd1 vssd1 vccd1 vccd1 _00959_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_31_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12912_ net386 _07460_ _07638_ vssd1 vssd1 vccd1 vccd1 _07654_ sky130_fd_sc_hd__and3_1
X_16680_ net360 _02352_ _02358_ _02228_ vssd1 vssd1 vccd1 vccd1 _02359_ sky130_fd_sc_hd__o211a_1
XFILLER_0_96_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_518 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13892_ _05813_ net52 vssd1 vssd1 vccd1 vccd1 _08149_ sky130_fd_sc_hd__nor2_2
X_15631_ ag2.body\[447\] net125 _01621_ ag2.body\[439\] vssd1 vssd1 vccd1 vccd1 _00897_
+ sky130_fd_sc_hd__a22o_1
X_12843_ net1680 _07623_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[177\]
+ sky130_fd_sc_hd__and2_1
XANTENNA__12179__A net1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_551 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15562_ ag2.body\[497\] net185 _01614_ ag2.body\[489\] vssd1 vssd1 vccd1 vccd1 _00835_
+ sky130_fd_sc_hd__a22o_1
X_18350_ _03842_ _03844_ _03821_ vssd1 vssd1 vccd1 vccd1 _03846_ sky130_fd_sc_hd__a21o_1
XANTENNA__10239__A2 _04493_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17689__B net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_1157 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_4_15__f_clk_A clknet_3_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12774_ net2003 net647 _07590_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[141\]
+ sky130_fd_sc_hd__and3_1
XFILLER_0_69_787 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_275 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17301_ ag2.body\[344\] net739 net953 _04123_ _02979_ vssd1 vssd1 vccd1 vccd1 _02980_
+ sky130_fd_sc_hd__a221o_1
X_14513_ net821 ag2.body\[315\] _04108_ net1012 vssd1 vssd1 vccd1 vccd1 _08674_ sky130_fd_sc_hd__a22o_1
XFILLER_0_90_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11987__A2 net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11725_ img_gen.tracker.frame\[203\] net591 net566 vssd1 vssd1 vccd1 vccd1 _06697_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_68_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16085__S net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18281_ net529 _03779_ vssd1 vssd1 vccd1 vccd1 _01388_ sky130_fd_sc_hd__and2_1
X_15493_ ag2.body\[564\] net109 _01606_ ag2.body\[556\] vssd1 vssd1 vccd1 vccd1 _00774_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_29_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13189__A1 net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17232_ ag2.body\[445\] net703 net690 ag2.body\[447\] vssd1 vssd1 vccd1 vccd1 _02911_
+ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__14386__B1 ag2.body\[303\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14444_ net1030 ag2.body\[229\] vssd1 vssd1 vccd1 vccd1 _08605_ sky130_fd_sc_hd__or2_1
XANTENNA__16470__S1 net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11656_ net1094 net1045 vssd1 vssd1 vccd1 vccd1 _06629_ sky130_fd_sc_hd__nand2_1
XANTENNA__12626__B _06639_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout90 net91 vssd1 vssd1 vccd1 vccd1 net90 sky130_fd_sc_hd__buf_2
XFILLER_0_65_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10607_ _05576_ _05577_ _05578_ _05579_ vssd1 vssd1 vccd1 vccd1 _05580_ sky130_fd_sc_hd__a22o_1
XFILLER_0_52_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17163_ ag2.body\[592\] net879 vssd1 vssd1 vccd1 vccd1 _02842_ sky130_fd_sc_hd__nand2_1
X_14375_ net973 ag2.body\[419\] vssd1 vssd1 vccd1 vccd1 _08536_ sky130_fd_sc_hd__nand2_1
XFILLER_0_135_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16127__A1 net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15002__B net58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10427__A net1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11587_ net773 net588 vssd1 vssd1 vccd1 vccd1 _06560_ sky130_fd_sc_hd__nand2_1
XFILLER_0_52_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16114_ net347 _01792_ vssd1 vssd1 vccd1 vccd1 _01793_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_94_3175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_3186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13326_ net275 _07842_ _07843_ net2031 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[440\]
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_111_3710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17094_ _02771_ _02772_ _02770_ vssd1 vssd1 vccd1 vccd1 _02773_ sky130_fd_sc_hd__or3b_1
Xhold909 control.body\[966\] vssd1 vssd1 vccd1 vccd1 net2471 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_827 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10538_ ag2.body\[229\] net1111 vssd1 vssd1 vccd1 vccd1 _05511_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_111_3721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_3197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14689__A1 net1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14689__B2 net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16045_ net352 _01720_ vssd1 vssd1 vccd1 vccd1 _01724_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_10_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13257_ net280 _07815_ _07816_ net1992 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[398\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_86_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12642__A net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10469_ _05438_ _05439_ _05440_ _05441_ vssd1 vssd1 vccd1 vccd1 _05442_ sky130_fd_sc_hd__a22o_1
XANTENNA__16114__A net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19256__RESET_B net1484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18032__C net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12208_ score_detect.sig_out\[0\] _04271_ _04948_ vssd1 vssd1 vccd1 vccd1 _07180_
+ sky130_fd_sc_hd__o21a_1
XANTENNA__12164__A2 net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13188_ net263 _07783_ _07784_ net1993 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[361\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11372__B1 net1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_1304 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1247 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17722__S1 net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11911__A2 net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11258__A net1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19804_ clknet_leaf_125_clk _00748_ net1410 vssd1 vssd1 vccd1 vccd1 ag2.body\[586\]
+ sky130_fd_sc_hd__dfrtp_4
X_12139_ net562 _07107_ _07108_ _07110_ vssd1 vssd1 vccd1 vccd1 _07111_ sky130_fd_sc_hd__a22o_1
X_17996_ net46 _03611_ vssd1 vssd1 vccd1 vccd1 _03612_ sky130_fd_sc_hd__nor2_1
XFILLER_0_100_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_109_3650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16850__A2 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_3661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19735_ clknet_leaf_132_clk _00679_ net1304 vssd1 vssd1 vccd1 vccd1 control.body\[661\]
+ sky130_fd_sc_hd__dfrtp_1
X_16947_ _04140_ net852 net940 _04141_ _02625_ vssd1 vssd1 vccd1 vccd1 _02626_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_105_3514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_3525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_3536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18052__A1 net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10478__A2 _04695_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19666_ clknet_leaf_134_clk _00610_ net1390 vssd1 vssd1 vccd1 vccd1 control.body\[720\]
+ sky130_fd_sc_hd__dfrtp_1
X_16878_ ag2.body\[16\] net880 vssd1 vssd1 vccd1 vccd1 _02557_ sky130_fd_sc_hd__xor2_1
XFILLER_0_126_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18617_ clknet_leaf_145_clk img_gen.tracker.next_frame\[55\] net1241 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[55\] sky130_fd_sc_hd__dfrtp_1
X_15829_ ag2.body\[271\] net201 _01643_ ag2.body\[263\] vssd1 vssd1 vccd1 vccd1 _01073_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_56_1067 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1213 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19597_ clknet_leaf_118_clk _00541_ net1390 vssd1 vssd1 vccd1 vccd1 control.body\[795\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15810__B1 _01641_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09350_ sound_gen.osc1.stayCount\[22\] _04351_ vssd1 vssd1 vccd1 vccd1 _04353_ sky130_fd_sc_hd__or2_1
X_18548_ clknet_leaf_132_clk _00074_ net1304 vssd1 vssd1 vccd1 vccd1 ag2.y\[0\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__17599__B net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19922__CLK clknet_leaf_51_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_118_3908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11978__A2 net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_118_3919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09281_ sound_gen.posDetector1.N\[1\] sound_gen.posDetector1.N\[0\] sound_gen.osc1.keepCounting
+ vssd1 vssd1 vccd1 vccd1 _04304_ sky130_fd_sc_hd__nor3_1
XFILLER_0_117_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18479_ net1512 net1507 vssd1 vssd1 vccd1 vccd1 _00010_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_60_2142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12817__A net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11280__X _06253_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_2153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20510_ clknet_leaf_112_clk track.nextHighScore\[0\] net1403 vssd1 vssd1 vccd1 vccd1
+ track.highScore\[0\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_60_2164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkload62_A clknet_leaf_51_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16008__B net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12927__A1 net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20441_ clknet_leaf_25_clk _01328_ net1343 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[77\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_127_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16723__S net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout123_A net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_2661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_77_2672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20372_ clknet_leaf_26_clk _01259_ net1343 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[8\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__15847__B net59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10056__B net1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_2683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload60 clknet_leaf_24_clk vssd1 vssd1 vccd1 vccd1 clkload60/Y sky130_fd_sc_hd__inv_16
XFILLER_0_113_575 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload71 clknet_leaf_47_clk vssd1 vssd1 vccd1 vccd1 clkload71/Y sky130_fd_sc_hd__inv_8
XTAP_TAPCELL_ROW_73_2536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_2082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload82 clknet_leaf_122_clk vssd1 vssd1 vccd1 vccd1 clkload82/Y sky130_fd_sc_hd__clkinv_8
XTAP_TAPCELL_ROW_58_2093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1032_A ag2.randCord\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_2558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload93 clknet_leaf_111_clk vssd1 vssd1 vccd1 vccd1 clkload93/Y sky130_fd_sc_hd__inv_12
XFILLER_0_45_1472 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1359 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13367__B net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15629__B1 _01621_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout492_A _01736_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16959__A ag2.body\[288\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17713__S1 net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11168__A net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10072__A net1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08996_ ag2.body\[94\] vssd1 vssd1 vccd1 vccd1 _04021_ sky130_fd_sc_hd__inv_2
XANTENNA__20513__RESET_B net1403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout280_X net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14479__A net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14852__A1 _08485_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout378_X net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout757_A _04232_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1499_A net1504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13383__A net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09617_ net778 control.body\[801\] control.body\[804\] net758 vssd1 vssd1 vccd1 vccd1
+ _04590_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__16694__A net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout545_X net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1287_X net1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09548_ net897 net904 _04446_ net636 vssd1 vssd1 vccd1 vccd1 _04521_ sky130_fd_sc_hd__a31o_1
XFILLER_0_6_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout36_A _03706_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11969__A2 net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_134_4400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_1416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_134_4411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09479_ ag2.body\[465\] net782 net768 ag2.body\[467\] vssd1 vssd1 vccd1 vccd1 _04452_
+ sky130_fd_sc_hd__o22a_1
XANTENNA_fanout712_X net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_144_clk clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_144_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_134_4422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12727__A net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11190__X _06163_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11510_ _06481_ _06480_ vssd1 vssd1 vccd1 vccd1 _06483_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_109_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12490_ net334 _07438_ vssd1 vssd1 vccd1 vccd1 _07439_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_24_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11350__B net1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11441_ net1060 control.body\[959\] vssd1 vssd1 vccd1 vccd1 _06414_ sky130_fd_sc_hd__xor2_1
XFILLER_0_0_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14160_ net996 _04222_ ag2.body\[623\] net790 vssd1 vssd1 vccd1 vccd1 _08321_ sky130_fd_sc_hd__o22a_1
X_11372_ ag2.body\[474\] net774 net1155 _04169_ _06344_ vssd1 vssd1 vccd1 vccd1 _06345_
+ sky130_fd_sc_hd__a221o_1
XANTENNA__08940__A net994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_1127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13111_ net344 _07578_ vssd1 vssd1 vccd1 vccd1 _07748_ sky130_fd_sc_hd__or2_1
XFILLER_0_0_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10323_ ag2.body\[609\] net1195 vssd1 vssd1 vccd1 vccd1 _05296_ sky130_fd_sc_hd__xor2_1
X_14091_ net1031 ag2.body\[285\] vssd1 vssd1 vccd1 vccd1 _08252_ sky130_fd_sc_hd__or2_1
XANTENNA__12462__A net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_4215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_4226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13042_ net279 _07713_ _07714_ net1969 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[284\]
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_128_4237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10254_ net1130 control.body\[788\] vssd1 vssd1 vccd1 vccd1 _05227_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_123_1459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_37_1443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10157__B2 ag2.body\[61\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1201 net1202 vssd1 vssd1 vccd1 vccd1 net1201 sky130_fd_sc_hd__buf_4
Xfanout1212 net1213 vssd1 vssd1 vccd1 vccd1 net1212 sky130_fd_sc_hd__clkbuf_8
XANTENNA__18282__A1 net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17085__A2 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17850_ img_gen.updater.commands.rR1.rainbowRNG\[13\] _03505_ vssd1 vssd1 vccd1 vccd1
+ _03506_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_33_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10185_ ag2.body\[422\] net1081 vssd1 vssd1 vccd1 vccd1 _05158_ sky130_fd_sc_hd__xor2_1
XFILLER_0_121_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1223 net1224 vssd1 vssd1 vccd1 vccd1 net1223 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_24_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_33_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1234 net1238 vssd1 vssd1 vccd1 vccd1 net1234 sky130_fd_sc_hd__buf_4
XANTENNA__16588__B net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16801_ _02475_ _02479_ _02057_ vssd1 vssd1 vccd1 vccd1 _02480_ sky130_fd_sc_hd__o21ai_1
Xfanout1245 net1250 vssd1 vssd1 vccd1 vccd1 net1245 sky130_fd_sc_hd__clkbuf_2
Xfanout1256 net1257 vssd1 vssd1 vccd1 vccd1 net1256 sky130_fd_sc_hd__buf_2
X_17781_ net2189 net516 _04398_ _03457_ _03459_ vssd1 vssd1 vccd1 vccd1 _01209_ sky130_fd_sc_hd__o32a_1
Xfanout1267 net1287 vssd1 vssd1 vccd1 vccd1 net1267 sky130_fd_sc_hd__buf_2
X_14993_ _05937_ net65 vssd1 vssd1 vccd1 vccd1 _01551_ sky130_fd_sc_hd__and2_2
Xfanout1278 net1280 vssd1 vssd1 vccd1 vccd1 net1278 sky130_fd_sc_hd__clkbuf_4
Xfanout280 net282 vssd1 vssd1 vccd1 vccd1 net280 sky130_fd_sc_hd__clkbuf_4
Xfanout291 net294 vssd1 vssd1 vccd1 vccd1 net291 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_79_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1289 net1291 vssd1 vssd1 vccd1 vccd1 net1289 sky130_fd_sc_hd__clkbuf_2
X_19520_ clknet_leaf_121_clk _00464_ net1402 vssd1 vssd1 vccd1 vccd1 control.body\[878\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13293__A _07476_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16732_ obsg2.obstacleArray\[96\] net490 net486 obsg2.obstacleArray\[98\] _02410_
+ vssd1 vssd1 vccd1 vccd1 _02411_ sky130_fd_sc_hd__a221o_1
X_13944_ ag2.body\[86\] net197 _08154_ ag2.body\[78\] vssd1 vssd1 vccd1 vccd1 _00167_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_88_315 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19451_ clknet_leaf_109_clk _00395_ net1416 vssd1 vssd1 vccd1 vccd1 control.body\[937\]
+ sky130_fd_sc_hd__dfrtp_1
X_16663_ obsg2.obstacleArray\[20\] obsg2.obstacleArray\[21\] net447 vssd1 vssd1 vccd1
+ vccd1 _02342_ sky130_fd_sc_hd__mux2_1
X_13875_ ag2.body\[24\] net115 _08147_ ag2.body\[16\] vssd1 vssd1 vccd1 vccd1 _00105_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_134_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18402_ _04644_ _08025_ _03890_ vssd1 vssd1 vccd1 vccd1 _03892_ sky130_fd_sc_hd__o21ai_1
X_15614_ ag2.body\[463\] net123 _01620_ ag2.body\[455\] vssd1 vssd1 vccd1 vccd1 _00881_
+ sky130_fd_sc_hd__a22o_1
X_12826_ net262 _07613_ _07614_ net2063 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[169\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_9_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19382_ clknet_leaf_102_clk _00326_ net1426 vssd1 vssd1 vccd1 vccd1 control.body\[1012\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16594_ _02271_ _02272_ net394 vssd1 vssd1 vccd1 vccd1 _02273_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18333_ net906 net638 _04638_ _04641_ net902 vssd1 vssd1 vccd1 vccd1 _03829_ sky130_fd_sc_hd__a2111o_1
X_12757_ net683 _07582_ vssd1 vssd1 vccd1 vccd1 _07583_ sky130_fd_sc_hd__nor2_1
X_15545_ ag2.body\[515\] net162 _01580_ ag2.body\[507\] vssd1 vssd1 vccd1 vccd1 _00821_
+ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_135_clk clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_135_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_57_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_1290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11708_ img_gen.tracker.frame\[299\] net591 net552 img_gen.tracker.frame\[296\] _06679_
+ vssd1 vssd1 vccd1 vccd1 _06680_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_96_3237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18264_ _03530_ _03547_ _03549_ vssd1 vssd1 vccd1 vccd1 _03771_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_13_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15476_ ag2.body\[581\] net111 _01604_ ag2.body\[573\] vssd1 vssd1 vccd1 vccd1 _00759_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_96_3248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12688_ net673 _07549_ vssd1 vssd1 vccd1 vccd1 _07550_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_96_3259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17215_ ag2.body\[49\] net731 net688 ag2.body\[55\] _02891_ vssd1 vssd1 vccd1 vccd1
+ _02894_ sky130_fd_sc_hd__a221o_1
XFILLER_0_25_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14427_ net1019 ag2.body\[558\] vssd1 vssd1 vccd1 vccd1 _08588_ sky130_fd_sc_hd__xor2_1
XFILLER_0_126_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11639_ _06521_ _06555_ _06610_ _06611_ _06562_ vssd1 vssd1 vccd1 vccd1 _06612_ sky130_fd_sc_hd__o221a_1
X_18195_ obsg2.obstacleArray\[94\] _03736_ net526 vssd1 vssd1 vccd1 vccd1 _01345_
+ sky130_fd_sc_hd__o21a_1
XANTENNA__15571__A2 net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_548 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14358_ net994 _04142_ ag2.body\[403\] net819 vssd1 vssd1 vccd1 vccd1 _08519_ sky130_fd_sc_hd__a22o_1
XFILLER_0_108_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17146_ ag2.body\[613\] net946 vssd1 vssd1 vccd1 vccd1 _02825_ sky130_fd_sc_hd__nand2_1
XFILLER_0_68_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_3_clk_A clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold706 control.body\[659\] vssd1 vssd1 vccd1 vccd1 net2268 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__18043__B _03554_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold717 control.body\[948\] vssd1 vssd1 vccd1 vccd1 net2279 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_873 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13309_ net2066 net648 _07837_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[429\]
+ sky130_fd_sc_hd__and3_1
XANTENNA__10935__A3 _05897_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold728 ag2.body\[221\] vssd1 vssd1 vccd1 vccd1 net2290 sky130_fd_sc_hd__dlygate4sd3_1
X_17077_ ag2.body\[199\] obsg2.randCord\[7\] vssd1 vssd1 vccd1 vccd1 _02756_ sky130_fd_sc_hd__xor2_1
X_14289_ net812 ag2.body\[476\] vssd1 vssd1 vccd1 vccd1 _08450_ sky130_fd_sc_hd__nor2_1
Xhold739 coll.badColl vssd1 vssd1 vccd1 vccd1 net2301 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1635 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__20302__CLK clknet_leaf_37_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16028_ net883 net948 vssd1 vssd1 vccd1 vccd1 _01707_ sky130_fd_sc_hd__xnor2_2
XANTENNA__17882__B _04758_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17979_ _01714_ _03540_ net298 vssd1 vssd1 vccd1 vccd1 _03600_ sky130_fd_sc_hd__and3_1
X_19718_ clknet_leaf_133_clk _00662_ net1308 vssd1 vssd1 vccd1 vccd1 control.body\[676\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_46_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_85_2930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11435__B net1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19649_ clknet_leaf_128_clk _00593_ net1329 vssd1 vssd1 vccd1 vccd1 control.body\[751\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_66_2340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16587__A1 net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_2805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_2351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16718__S net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09402_ sound_gen.osc1.stayCount\[2\] _04342_ net270 vssd1 vssd1 vccd1 vccd1 _04385_
+ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_62_2204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_62_2215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_2226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18328__A2 _04519_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18218__B net40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09333_ net2173 _04334_ vssd1 vssd1 vccd1 vccd1 _04340_ sky130_fd_sc_hd__nor2_1
XFILLER_0_47_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17122__B net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout240_A net242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_126_clk clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_126_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_8_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17536__B1 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11451__A net1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout338_A net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17000__A2 net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09264_ sound_gen.osc1.timer\[2\] _04285_ _04284_ vssd1 vssd1 vccd1 vccd1 _04288_
+ sky130_fd_sc_hd__o21bai_4
XFILLER_0_63_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_79_2723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16961__B net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_2734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_2745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10067__A net1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09195_ ag2.body\[611\] vssd1 vssd1 vccd1 vccd1 _04220_ sky130_fd_sc_hd__inv_2
XFILLER_0_90_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_75_2609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1247_A net1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11179__A3 _06137_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20424_ clknet_leaf_38_clk _01311_ net1355 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[60\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__09856__A _04772_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_56_2019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_1594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13378__A net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20355_ clknet_leaf_140_clk _01246_ net1291 vssd1 vssd1 vccd1 vccd1 img_gen.updater.commands.rR1.rainbowRNG\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09575__B net1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1035_X net1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1414_A net1415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_534 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20286_ clknet_leaf_35_clk control.divider.next_count\[7\] net1348 vssd1 vssd1 vccd1
+ vccd1 control.divider.count\[7\] sky130_fd_sc_hd__dfrtp_2
XANTENNA_fanout495_X net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout874_A net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10514__B net1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_1470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1202_X net1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold11 score_detect.N\[1\] vssd1 vssd1 vccd1 vccd1 net1573 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__18842__CLK clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09591__A net1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold22 ag2.body\[574\] vssd1 vssd1 vccd1 vccd1 net1584 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__16814__A2 net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold33 img_gen.tracker.frame\[104\] vssd1 vssd1 vccd1 vccd1 net1595 sky130_fd_sc_hd__dlygate4sd3_1
X_08979_ ag2.body\[73\] vssd1 vssd1 vccd1 vccd1 _04004_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout662_X net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold44 img_gen.tracker.frame\[117\] vssd1 vssd1 vccd1 vccd1 net1606 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14825__A1 net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold55 img_gen.tracker.frame\[5\] vssd1 vssd1 vccd1 vccd1 net1617 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14825__B2 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold66 control.fsm.temp\[1\] vssd1 vssd1 vccd1 vccd1 net1628 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11639__A1 _06521_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold77 img_gen.tracker.frame\[3\] vssd1 vssd1 vccd1 vccd1 net1639 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14002__A net1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold88 img_gen.tracker.frame\[110\] vssd1 vssd1 vccd1 vccd1 net1650 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10530__A net1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11990_ img_gen.tracker.frame\[385\] net618 net546 img_gen.tracker.frame\[391\] vssd1
+ vssd1 vccd1 vccd1 _06962_ sky130_fd_sc_hd__o22a_1
Xhold99 img_gen.tracker.frame\[325\] vssd1 vssd1 vccd1 vccd1 net1661 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_19_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11345__B net1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10941_ ag2.body\[300\] net1142 vssd1 vssd1 vccd1 vccd1 _05914_ sky130_fd_sc_hd__xor2_1
XANTENNA_fanout927_X net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18992__CLK clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13841__A net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13660_ net825 _08013_ vssd1 vssd1 vccd1 vccd1 _08014_ sky130_fd_sc_hd__nor2_1
XFILLER_0_97_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10872_ ag2.body\[529\] net1203 vssd1 vssd1 vccd1 vccd1 _05845_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_45_1701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout39_X net39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12611_ net252 _07506_ _07507_ net1645 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[61\]
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_26_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13591_ _03961_ control.divider.count\[9\] control.divider.count\[8\] _07953_ vssd1
+ vssd1 vccd1 vccd1 _07966_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_117_clk clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_117_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_26_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15330_ net2350 net74 _01587_ control.body\[698\] vssd1 vssd1 vccd1 vccd1 _00628_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__19348__CLK clknet_leaf_102_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1295 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12542_ net2027 net653 _07469_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[30\]
+ sky130_fd_sc_hd__and3_1
XANTENNA__10614__A2 _05572_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17967__B _03531_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09480__A2 net1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15261_ control.body\[775\] net97 net50 net2162 vssd1 vssd1 vccd1 vccd1 _00569_ sky130_fd_sc_hd__a22o_1
XANTENNA__11080__B net1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12473_ _07426_ _07427_ vssd1 vssd1 vccd1 vccd1 _07428_ sky130_fd_sc_hd__and2b_1
XFILLER_0_123_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14212_ _08369_ _08370_ _08371_ _08372_ vssd1 vssd1 vccd1 vccd1 _08373_ sky130_fd_sc_hd__or4_1
X_17000_ _04036_ net889 net866 _04037_ vssd1 vssd1 vccd1 vccd1 _02679_ sky130_fd_sc_hd__a22o_1
XANTENNA__20325__CLK clknet_4_7__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_3101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_91_3112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11424_ _06181_ _06394_ _06395_ _06396_ vssd1 vssd1 vccd1 vccd1 _06397_ sky130_fd_sc_hd__or4_1
X_15192_ control.body\[824\] net94 _01573_ net2497 vssd1 vssd1 vccd1 vccd1 _00506_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_22_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11575__B1 net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_8 _03442_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19498__CLK clknet_leaf_113_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14143_ net1037 ag2.body\[172\] vssd1 vssd1 vccd1 vccd1 _08304_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_39_1516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13288__A _07472_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11355_ net1075 control.body\[814\] vssd1 vssd1 vccd1 vccd1 _06328_ sky130_fd_sc_hd__xor2_1
XFILLER_0_21_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_39_1527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12192__A net1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10306_ net1193 control.body\[697\] vssd1 vssd1 vccd1 vccd1 _05279_ sky130_fd_sc_hd__xor2_1
X_14074_ net808 ag2.body\[213\] ag2.body\[215\] net794 _08228_ vssd1 vssd1 vccd1 vccd1
+ _08235_ sky130_fd_sc_hd__o221a_1
X_18951_ clknet_leaf_5_clk img_gen.tracker.next_frame\[389\] net1268 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[389\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_120_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11286_ net1159 control.body\[1107\] vssd1 vssd1 vccd1 vccd1 _06259_ sky130_fd_sc_hd__xor2_1
XFILLER_0_67_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13867__A2 _04519_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17058__A2 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17902_ net530 _03537_ vssd1 vssd1 vccd1 vccd1 _01251_ sky130_fd_sc_hd__and2_1
X_13025_ net288 _07705_ _07706_ net1921 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[275\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_123_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10237_ ag2.body\[321\] net1211 vssd1 vssd1 vccd1 vccd1 _05210_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_89_3030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_3041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18882_ clknet_leaf_11_clk img_gen.tracker.next_frame\[320\] net1283 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[320\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_89_3052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1020 net1022 vssd1 vssd1 vccd1 vccd1 net1020 sky130_fd_sc_hd__buf_4
Xfanout1031 ag2.randCord\[5\] vssd1 vssd1 vccd1 vccd1 net1031 sky130_fd_sc_hd__buf_4
Xfanout1042 ag2.randCord\[4\] vssd1 vssd1 vccd1 vccd1 net1042 sky130_fd_sc_hd__buf_8
XANTENNA__16805__A2 net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17833_ net662 _03493_ vssd1 vssd1 vccd1 vccd1 _01226_ sky130_fd_sc_hd__and2_1
Xfanout1053 net1069 vssd1 vssd1 vccd1 vccd1 net1053 sky130_fd_sc_hd__buf_2
X_10168_ ag2.body\[577\] net1196 vssd1 vssd1 vccd1 vccd1 _05141_ sky130_fd_sc_hd__xor2_1
XANTENNA__17207__B net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14816__A1 net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1064 net1068 vssd1 vssd1 vccd1 vccd1 net1064 sky130_fd_sc_hd__buf_4
XANTENNA__18007__A1 net38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1075 net1077 vssd1 vssd1 vccd1 vccd1 net1075 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_89_602 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1086 net1093 vssd1 vssd1 vccd1 vccd1 net1086 sky130_fd_sc_hd__buf_2
X_17764_ _03289_ _03299_ _02742_ _03276_ vssd1 vssd1 vccd1 vccd1 _03443_ sky130_fd_sc_hd__and4b_1
XANTENNA__10440__A net1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1097 net1098 vssd1 vssd1 vccd1 vccd1 net1097 sky130_fd_sc_hd__clkbuf_8
XANTENNA__16018__A0 net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10099_ _05068_ _05069_ _05070_ _05071_ vssd1 vssd1 vccd1 vccd1 _05072_ sky130_fd_sc_hd__or4_1
X_14976_ _04607_ _01549_ vssd1 vssd1 vccd1 vccd1 _01550_ sky130_fd_sc_hd__and2b_2
X_19503_ clknet_leaf_113_clk _00447_ net1396 vssd1 vssd1 vccd1 vccd1 control.body\[893\]
+ sky130_fd_sc_hd__dfrtp_1
X_16715_ obsg2.obstacleArray\[124\] net491 net482 obsg2.obstacleArray\[125\] _02393_
+ vssd1 vssd1 vccd1 vccd1 _02394_ sky130_fd_sc_hd__a221o_1
XANTENNA__16569__A1 net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13927_ ag2.body\[71\] net134 _08152_ ag2.body\[63\] vssd1 vssd1 vccd1 vccd1 _00152_
+ sky130_fd_sc_hd__a22o_1
X_17695_ ag2.body\[159\] net693 net728 ag2.body\[154\] vssd1 vssd1 vccd1 vccd1 _03374_
+ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__14847__A _08280_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17230__A2 net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19434_ clknet_leaf_108_clk _00378_ net1423 vssd1 vssd1 vccd1 vccd1 control.body\[952\]
+ sky130_fd_sc_hd__dfrtp_1
X_16646_ _02322_ _02323_ _02324_ net395 net361 vssd1 vssd1 vccd1 vccd1 _02325_ sky130_fd_sc_hd__a221o_1
X_13858_ ag2.body\[21\] net116 _08134_ ag2.body\[13\] vssd1 vssd1 vccd1 vccd1 _00101_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_88_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_18_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18038__B net42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13470__B net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12809_ net253 _07605_ _07606_ net1817 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[160\]
+ sky130_fd_sc_hd__a22o_1
X_19365_ clknet_leaf_102_clk _00309_ net1438 vssd1 vssd1 vccd1 vccd1 control.body\[1027\]
+ sky130_fd_sc_hd__dfrtp_1
X_16577_ net395 _02255_ _02254_ net359 vssd1 vssd1 vccd1 vccd1 _02256_ sky130_fd_sc_hd__a211o_1
Xclkbuf_leaf_108_clk clknet_4_10__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_108_clk
+ sky130_fd_sc_hd__clkbuf_8
X_13789_ _04390_ _07209_ net320 vssd1 vssd1 vccd1 vccd1 _08096_ sky130_fd_sc_hd__a21o_1
XFILLER_0_2_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18316_ _08137_ _03810_ vssd1 vssd1 vccd1 vccd1 _03812_ sky130_fd_sc_hd__nand2_1
XANTENNA__11802__A1 net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15528_ ag2.body\[531\] net157 _01610_ ag2.body\[523\] vssd1 vssd1 vccd1 vccd1 _00805_
+ sky130_fd_sc_hd__a22o_1
X_19296_ clknet_leaf_98_clk _00240_ net1446 vssd1 vssd1 vccd1 vccd1 control.body\[1102\]
+ sky130_fd_sc_hd__dfrtp_1
X_18247_ obsg2.obstacleArray\[120\] _03762_ net524 vssd1 vssd1 vccd1 vccd1 _01371_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_115_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18715__CLK clknet_leaf_144_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15459_ ag2.body\[598\] net86 _01602_ net2387 vssd1 vssd1 vccd1 vccd1 _00744_ sky130_fd_sc_hd__a22o_1
XANTENNA__15544__A2 net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18054__A net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19271__RESET_B net1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18178_ _03617_ net41 vssd1 vssd1 vccd1 vccd1 _03728_ sky130_fd_sc_hd__nor2_1
XANTENNA__10369__A1 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_270 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19200__RESET_B net1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_367 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10369__B2 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold503 img_gen.tracker.frame\[192\] vssd1 vssd1 vccd1 vccd1 net2065 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17297__A2 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold514 img_gen.tracker.frame\[120\] vssd1 vssd1 vccd1 vccd1 net2076 sky130_fd_sc_hd__dlygate4sd3_1
X_17129_ ag2.body\[514\] net727 net719 ag2.body\[515\] vssd1 vssd1 vccd1 vccd1 _02808_
+ sky130_fd_sc_hd__o22a_1
Xhold525 img_gen.tracker.frame\[537\] vssd1 vssd1 vccd1 vccd1 net2087 sky130_fd_sc_hd__dlygate4sd3_1
Xhold536 img_gen.tracker.frame\[97\] vssd1 vssd1 vccd1 vccd1 net2098 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10615__A net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold547 img_gen.tracker.frame\[285\] vssd1 vssd1 vccd1 vccd1 net2109 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13307__A1 net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09951_ net1170 control.body\[738\] vssd1 vssd1 vccd1 vccd1 _04924_ sky130_fd_sc_hd__nand2b_1
Xhold558 control.body\[1023\] vssd1 vssd1 vccd1 vccd1 net2120 sky130_fd_sc_hd__dlygate4sd3_1
X_20140_ clknet_leaf_96_clk _01084_ net1449 vssd1 vssd1 vccd1 vccd1 ag2.body\[250\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_12_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold569 img_gen.tracker.frame\[567\] vssd1 vssd1 vccd1 vccd1 net2131 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkload25_A clknet_leaf_15_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10334__B net1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09882_ ag2.body\[160\] net784 net763 ag2.body\[164\] _04854_ vssd1 vssd1 vccd1 vccd1
+ _04855_ sky130_fd_sc_hd__a221o_1
X_20071_ clknet_leaf_73_clk _01015_ net1500 vssd1 vssd1 vccd1 vccd1 ag2.body\[325\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__12830__A net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout190_A net191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1042 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_2402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_1549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11446__A net1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout455_A net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18229__A net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13661__A net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1612 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1197_A net1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_1572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10844__A2 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout622_A net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1364_A net1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09316_ sound_gen.osc1.count\[3\] _04321_ _04319_ vssd1 vssd1 vccd1 vccd1 _04332_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_134_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09247_ img_gen.updater.commands.cmd_num\[1\] vssd1 vssd1 vccd1 vccd1 _04272_ sky130_fd_sc_hd__inv_2
XFILLER_0_63_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1152_X net1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout508_X net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09586__A net1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09178_ ag2.body\[553\] vssd1 vssd1 vccd1 vccd1 _04203_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout991_A net995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20498__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20407_ clknet_leaf_31_clk _01294_ net1346 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[43\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_107_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10525__A net1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput12 net12 vssd1 vssd1 vccd1 vccd1 gpio_out[11] sky130_fd_sc_hd__buf_2
X_11140_ ag2.body\[412\] net1139 vssd1 vssd1 vccd1 vccd1 _06113_ sky130_fd_sc_hd__xor2_1
Xoutput23 net23 vssd1 vssd1 vccd1 vccd1 gpio_out[21] sky130_fd_sc_hd__buf_2
X_20338_ clknet_leaf_21_clk _01229_ net1363 vssd1 vssd1 vccd1 vccd1 ag2.apple_cord\[6\]
+ sky130_fd_sc_hd__dfstp_1
Xoutput34 net34 vssd1 vssd1 vccd1 vccd1 gpio_out[9] sky130_fd_sc_hd__buf_2
XANTENNA__19790__CLK clknet_leaf_127_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1520 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout877_X net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17953__D net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11071_ ag2.body\[361\] net1209 vssd1 vssd1 vccd1 vccd1 _06044_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_25_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20269_ clknet_leaf_36_clk net1568 net1347 vssd1 vssd1 vccd1 vccd1 control.detect1.Q\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__16248__B1 _01919_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09922__B1 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10022_ _04988_ _04989_ _04990_ _04994_ vssd1 vssd1 vccd1 vccd1 _04995_ sky130_fd_sc_hd__or4_1
XFILLER_0_60_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11356__A net1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14830_ _08318_ _08319_ _08324_ _08645_ vssd1 vssd1 vccd1 vccd1 _01501_ sky130_fd_sc_hd__o31a_2
XANTENNA__10260__A net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_1460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14761_ net790 ag2.body\[47\] _08920_ _08921_ vssd1 vssd1 vccd1 vccd1 _08922_ sky130_fd_sc_hd__o211a_1
X_11973_ net571 _06942_ _06944_ _06941_ vssd1 vssd1 vccd1 vccd1 _06945_ sky130_fd_sc_hd__a31o_1
XANTENNA__17748__B1 _03098_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16358__S net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10296__B1 net1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16500_ net365 _02178_ _02075_ vssd1 vssd1 vccd1 vccd1 _02179_ sky130_fd_sc_hd__a21o_1
XFILLER_0_54_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10924_ _05894_ _05895_ _05896_ vssd1 vssd1 vccd1 vccd1 _05897_ sky130_fd_sc_hd__and3_2
XANTENNA__17212__A2 net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13712_ track.highScore\[2\] _04638_ net356 vssd1 vssd1 vccd1 vccd1 track.nextHighScore\[2\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17480_ ag2.body\[128\] net887 vssd1 vssd1 vccd1 vccd1 _03159_ sky130_fd_sc_hd__nand2_1
X_14692_ net1003 _04109_ ag2.body\[322\] net830 vssd1 vssd1 vccd1 vccd1 _08853_ sky130_fd_sc_hd__a22o_1
XANTENNA__19170__CLK clknet_leaf_53_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_113_Right_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16431_ _02108_ _02109_ net401 vssd1 vssd1 vccd1 vccd1 _02110_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13643_ control.divider.count\[15\] _08002_ net222 vssd1 vssd1 vccd1 vccd1 _08003_
+ sky130_fd_sc_hd__o21ai_1
XANTENNA__18738__CLK clknet_leaf_141_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10855_ net1167 control.body\[690\] vssd1 vssd1 vccd1 vccd1 _05828_ sky130_fd_sc_hd__xor2_1
XANTENNA__12187__A net1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19150_ clknet_leaf_51_clk _00094_ net1377 vssd1 vssd1 vccd1 vccd1 ag2.body\[14\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_82_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_16_clk_X clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09989__B1 _04937_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13574_ _03960_ control.divider.fsm.current_mode\[0\] vssd1 vssd1 vccd1 vccd1 _07949_
+ sky130_fd_sc_hd__nor2_2
X_16362_ obsg2.obstacleArray\[11\] net414 _02040_ net416 vssd1 vssd1 vccd1 vccd1 _02041_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_82_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10786_ net1195 control.body\[625\] vssd1 vssd1 vccd1 vccd1 _05759_ sky130_fd_sc_hd__or2_1
XFILLER_0_27_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18101_ net300 _03616_ vssd1 vssd1 vccd1 vccd1 _03683_ sky130_fd_sc_hd__nand2_1
XFILLER_0_93_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15313_ control.body\[722\] net77 _01588_ net2552 vssd1 vssd1 vccd1 vccd1 _00612_
+ sky130_fd_sc_hd__a22o_1
X_12525_ net227 _07458_ _07459_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[23\]
+ sky130_fd_sc_hd__o21bai_1
X_16293_ obsg2.obstacleArray\[116\] obsg2.obstacleArray\[117\] net408 vssd1 vssd1
+ vccd1 vccd1 _01972_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10063__A3 _04600_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19081_ clknet_leaf_29_clk img_gen.tracker.next_frame\[519\] net1334 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[519\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__16093__S net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18032_ net539 net432 net462 net489 vssd1 vssd1 vccd1 vccd1 _03638_ sky130_fd_sc_hd__and4_1
XFILLER_0_129_1443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12456_ _07318_ _07333_ _07411_ _07415_ vssd1 vssd1 vccd1 vccd1 _07416_ sky130_fd_sc_hd__a211o_1
X_15244_ control.body\[791\] net97 _01578_ net2372 vssd1 vssd1 vccd1 vccd1 _00553_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_48_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_456 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12634__B _07519_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11407_ ag2.body\[568\] net1228 vssd1 vssd1 vccd1 vccd1 _06380_ sky130_fd_sc_hd__xor2_1
X_15175_ net2653 net103 _01571_ net2363 vssd1 vssd1 vccd1 vccd1 _00491_ sky130_fd_sc_hd__a22o_1
XFILLER_0_23_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17279__A2 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10435__A net1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12387_ _07351_ vssd1 vssd1 vccd1 vccd1 _07352_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14126_ net990 _04131_ _04132_ net981 _08283_ vssd1 vssd1 vccd1 vccd1 _08287_ sky130_fd_sc_hd__a221o_1
XFILLER_0_120_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11338_ _06301_ _06302_ _06305_ _06307_ vssd1 vssd1 vccd1 vccd1 _06311_ sky130_fd_sc_hd__or4_1
X_19983_ clknet_leaf_64_clk _00927_ net1475 vssd1 vssd1 vccd1 vccd1 ag2.body\[413\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_103_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10154__B net1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18934_ clknet_leaf_139_clk img_gen.tracker.next_frame\[372\] net1288 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[372\] sky130_fd_sc_hd__dfrtp_1
X_14057_ net1015 ag2.body\[38\] vssd1 vssd1 vccd1 vccd1 _08218_ sky130_fd_sc_hd__xor2_1
X_11269_ ag2.body\[127\] net1067 vssd1 vssd1 vccd1 vccd1 _06242_ sky130_fd_sc_hd__nand2_1
XFILLER_0_103_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12650__A net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13008_ net342 _07523_ vssd1 vssd1 vccd1 vccd1 _07699_ sky130_fd_sc_hd__nor2_1
X_18865_ clknet_leaf_26_clk img_gen.tracker.next_frame\[303\] net1285 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[303\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__17987__B1 net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11720__B1 net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17816_ net924 _08124_ vssd1 vssd1 vccd1 vccd1 _03483_ sky130_fd_sc_hd__and2_1
XANTENNA__17451__A2 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18796_ clknet_leaf_17_clk img_gen.tracker.next_frame\[234\] net1319 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[234\] sky130_fd_sc_hd__dfrtp_1
X_17747_ _03420_ _03421_ _03423_ _03425_ vssd1 vssd1 vccd1 vccd1 _03426_ sky130_fd_sc_hd__and4_2
XANTENNA__11079__A2 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14959_ net2284 net172 _01547_ control.body\[1025\] vssd1 vssd1 vccd1 vccd1 _00299_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__18049__A net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13481__A net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17203__A2 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17678_ ag2.body\[472\] net737 net716 ag2.body\[475\] vssd1 vssd1 vccd1 vccd1 _03357_
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_76_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19417_ clknet_leaf_105_clk _00361_ net1432 vssd1 vssd1 vccd1 vccd1 control.body\[983\]
+ sky130_fd_sc_hd__dfrtp_1
X_16629_ net359 _02303_ _02307_ net358 vssd1 vssd1 vccd1 vccd1 _02308_ sky130_fd_sc_hd__o211a_1
XANTENNA__14864__X _01535_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16792__A net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19348_ clknet_leaf_102_clk _00292_ net1429 vssd1 vssd1 vccd1 vccd1 control.body\[1042\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09958__X _04931_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14973__B1 net51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09101_ ag2.body\[354\] vssd1 vssd1 vccd1 vccd1 _04126_ sky130_fd_sc_hd__inv_2
XANTENNA__11787__B1 net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19279_ clknet_leaf_97_clk _00223_ net1450 vssd1 vssd1 vccd1 vccd1 control.body\[1117\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11882__S0 net1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09032_ ag2.body\[181\] vssd1 vssd1 vccd1 vccd1 _04057_ sky130_fd_sc_hd__inv_2
XANTENNA__13528__A1 net226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold300 img_gen.tracker.frame\[347\] vssd1 vssd1 vccd1 vccd1 net1862 sky130_fd_sc_hd__dlygate4sd3_1
Xhold311 img_gen.tracker.frame\[170\] vssd1 vssd1 vccd1 vccd1 net1873 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout203_A net204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold322 img_gen.tracker.frame\[366\] vssd1 vssd1 vccd1 vccd1 net1884 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold333 img_gen.tracker.frame\[445\] vssd1 vssd1 vccd1 vccd1 net1895 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold344 img_gen.tracker.frame\[381\] vssd1 vssd1 vccd1 vccd1 net1906 sky130_fd_sc_hd__dlygate4sd3_1
Xhold355 img_gen.tracker.frame\[161\] vssd1 vssd1 vccd1 vccd1 net1917 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold366 img_gen.tracker.frame\[204\] vssd1 vssd1 vccd1 vccd1 net1928 sky130_fd_sc_hd__dlygate4sd3_1
Xhold377 img_gen.tracker.frame\[571\] vssd1 vssd1 vccd1 vccd1 net1939 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout802 net805 vssd1 vssd1 vccd1 vccd1 net802 sky130_fd_sc_hd__buf_4
XFILLER_0_106_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20123_ clknet_leaf_81_clk _01067_ net1486 vssd1 vssd1 vccd1 vccd1 ag2.body\[265\]
+ sky130_fd_sc_hd__dfrtp_4
Xhold388 img_gen.tracker.frame\[338\] vssd1 vssd1 vccd1 vccd1 net1950 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__17690__A2 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09934_ ag2.body\[27\] net1153 vssd1 vssd1 vccd1 vccd1 _04907_ sky130_fd_sc_hd__and2b_1
Xhold399 img_gen.tracker.frame\[368\] vssd1 vssd1 vccd1 vccd1 net1961 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_370 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout813 _03969_ vssd1 vssd1 vccd1 vccd1 net813 sky130_fd_sc_hd__clkbuf_4
XANTENNA__16032__A net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1112_A ag2.x\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12560__A net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout824 net831 vssd1 vssd1 vccd1 vccd1 net824 sky130_fd_sc_hd__buf_4
Xfanout835 net836 vssd1 vssd1 vccd1 vccd1 net835 sky130_fd_sc_hd__clkbuf_4
Xfanout846 net847 vssd1 vssd1 vccd1 vccd1 net846 sky130_fd_sc_hd__buf_4
Xfanout857 obsg2.randCord\[3\] vssd1 vssd1 vccd1 vccd1 net857 sky130_fd_sc_hd__clkbuf_8
X_09865_ ag2.body\[159\] net1065 vssd1 vssd1 vccd1 vccd1 _04838_ sky130_fd_sc_hd__or2_1
X_20054_ clknet_leaf_72_clk _00998_ net1503 vssd1 vssd1 vccd1 vccd1 ag2.body\[340\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_102_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input8_A gpio_in[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1000 control.body\[756\] vssd1 vssd1 vccd1 vccd1 net2562 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout868 net869 vssd1 vssd1 vccd1 vccd1 net868 sky130_fd_sc_hd__buf_4
XFILLER_0_77_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout572_A net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11711__B1 net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1011 control.body\[1086\] vssd1 vssd1 vccd1 vccd1 net2573 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout879 net881 vssd1 vssd1 vccd1 vccd1 net879 sky130_fd_sc_hd__buf_4
Xhold1022 control.body\[995\] vssd1 vssd1 vccd1 vccd1 net2584 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11176__A net1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10080__A net1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1033 control.body\[659\] vssd1 vssd1 vccd1 vccd1 net2595 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__19193__CLK clknet_leaf_53_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09796_ net1205 control.body\[961\] vssd1 vssd1 vccd1 vccd1 _04769_ sky130_fd_sc_hd__xor2_1
Xhold1044 control.body\[679\] vssd1 vssd1 vccd1 vccd1 net2606 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13094__C _07638_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1055 control.body\[1036\] vssd1 vssd1 vccd1 vccd1 net2617 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1066 control.body\[690\] vssd1 vssd1 vccd1 vccd1 net2628 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_1600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1077 control.body\[704\] vssd1 vssd1 vccd1 vccd1 net2639 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout360_X net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1088 control.body\[932\] vssd1 vssd1 vccd1 vccd1 net2650 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14487__A net993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16178__S net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1481_A net1482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1099 control.body\[928\] vssd1 vssd1 vccd1 vccd1 net2661 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout458_X net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout837_A net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout625_X net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19193__RESET_B net1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10640_ net1118 control.body\[668\] vssd1 vssd1 vccd1 vccd1 _05613_ sky130_fd_sc_hd__xor2_1
XANTENNA__14964__B1 _01547_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11778__B1 net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17310__B net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16166__C1 _01743_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10571_ net891 _04423_ _05238_ _05543_ vssd1 vssd1 vccd1 vccd1 _05544_ sky130_fd_sc_hd__o31a_2
XFILLER_0_64_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_283 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12310_ _07275_ _07276_ vssd1 vssd1 vccd1 vccd1 _07277_ sky130_fd_sc_hd__or2_1
X_13290_ net234 _07829_ _07830_ net1798 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[417\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_1_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout994_X net994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_787 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12241_ img_gen.updater.commands.count\[2\] _07190_ img_gen.updater.commands.count\[6\]
+ img_gen.updater.commands.count\[5\] vssd1 vssd1 vccd1 vccd1 _07211_ sky130_fd_sc_hd__o211a_1
XANTENNA__18458__A1 _05075_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10255__A net1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12172_ _07125_ _07131_ _07137_ _07143_ net472 net437 vssd1 vssd1 vccd1 vccd1 _07144_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_130_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11950__B1 net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11123_ net1202 control.body\[865\] vssd1 vssd1 vccd1 vccd1 _06096_ sky130_fd_sc_hd__nand2_1
XANTENNA_clkbuf_leaf_43_clk_A clknet_4_7__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09763__B net1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16980_ _04152_ net950 net941 _04153_ _02658_ vssd1 vssd1 vccd1 vccd1 _02659_ sky130_fd_sc_hd__o221a_1
X_11054_ _06020_ _06025_ _06026_ _04429_ vssd1 vssd1 vccd1 vccd1 _06027_ sky130_fd_sc_hd__and4bb_1
X_15931_ ag2.body\[169\] net136 _01655_ ag2.body\[161\] vssd1 vssd1 vccd1 vccd1 _01163_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__10505__A1 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10702__B net1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10505__B2 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11702__B1 _06671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10005_ _04974_ _04975_ _04976_ _04977_ _04973_ vssd1 vssd1 vccd1 vccd1 _04978_ sky130_fd_sc_hd__a221o_1
XANTENNA__17433__A2 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18650_ clknet_leaf_130_clk img_gen.tracker.next_frame\[88\] net1317 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[88\] sky130_fd_sc_hd__dfrtp_1
X_15862_ ag2.body\[237\] net175 _01646_ ag2.body\[229\] vssd1 vssd1 vccd1 vccd1 _01103_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_64_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__20513__CLK clknet_leaf_113_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17601_ ag2.body\[417\] net733 net725 ag2.body\[418\] _03279_ vssd1 vssd1 vccd1 vccd1
+ _03280_ sky130_fd_sc_hd__a221o_1
XANTENNA__16641__B1 net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_58_clk_A clknet_4_13__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14813_ net1000 ag2.body\[376\] vssd1 vssd1 vccd1 vccd1 _01484_ sky130_fd_sc_hd__xor2_1
XFILLER_0_73_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18581_ clknet_leaf_14_clk img_gen.tracker.next_frame\[19\] net1278 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[19\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_98_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15793_ ag2.body\[303\] net208 _01639_ ag2.body\[295\] vssd1 vssd1 vccd1 vccd1 _01041_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__18560__CLK clknet_leaf_132_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_101_clk_A clknet_4_11__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17532_ ag2.body\[276\] net965 vssd1 vssd1 vccd1 vccd1 _03211_ sky130_fd_sc_hd__xor2_1
X_14744_ net1033 ag2.body\[109\] vssd1 vssd1 vccd1 vccd1 _08905_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_19_1252 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11956_ net472 _06914_ _06927_ _06909_ net438 vssd1 vssd1 vccd1 vccd1 _06928_ sky130_fd_sc_hd__o221a_1
XFILLER_0_118_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12629__B net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_120_3970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_3981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10907_ net1192 control.body\[673\] vssd1 vssd1 vccd1 vccd1 _05880_ sky130_fd_sc_hd__xor2_1
XANTENNA__11533__B net1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17463_ ag2.body\[532\] net964 vssd1 vssd1 vccd1 vccd1 _03142_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_120_3992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14675_ _08834_ _08835_ _08832_ _08833_ vssd1 vssd1 vccd1 vccd1 _08836_ sky130_fd_sc_hd__a211o_1
X_11887_ img_gen.tracker.frame\[31\] net551 _06858_ net565 vssd1 vssd1 vccd1 vccd1
+ _06859_ sky130_fd_sc_hd__o211a_1
XFILLER_0_129_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_101_3391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_1206 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19202_ clknet_leaf_88_clk _00146_ net1459 vssd1 vssd1 vccd1 vccd1 ag2.body\[65\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_129_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16414_ obsg2.obstacleArray\[100\] obsg2.obstacleArray\[101\] net452 vssd1 vssd1
+ vccd1 vccd1 _02093_ sky130_fd_sc_hd__mux2_1
X_13626_ control.divider.count\[9\] _07990_ vssd1 vssd1 vccd1 vccd1 _07992_ sky130_fd_sc_hd__and2_1
X_10838_ _05803_ _05804_ _05805_ _05810_ vssd1 vssd1 vccd1 vccd1 _05811_ sky130_fd_sc_hd__or4_2
XFILLER_0_39_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14955__B1 _01546_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17394_ ag2.body\[508\] net712 net942 _04186_ vssd1 vssd1 vccd1 vccd1 _03073_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__10149__B net1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09582__A_N net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_116_clk_A clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19133_ clknet_leaf_140_clk img_gen.tracker.next_frame\[571\] net1296 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[571\] sky130_fd_sc_hd__dfrtp_1
X_16345_ obsg2.obstacleArray\[88\] obsg2.obstacleArray\[89\] net411 vssd1 vssd1 vccd1
+ vccd1 _02024_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13557_ ssdec1.in\[2\] ssdec1.in\[3\] _07938_ vssd1 vssd1 vccd1 vccd1 _07939_ sky130_fd_sc_hd__and3b_1
X_10769_ ag2.body\[218\] net1184 vssd1 vssd1 vccd1 vccd1 _05742_ sky130_fd_sc_hd__xor2_1
XFILLER_0_67_1504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12508_ net2059 net649 _07450_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[15\]
+ sky130_fd_sc_hd__and3_1
X_19064_ clknet_leaf_9_clk img_gen.tracker.next_frame\[502\] net1272 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[502\] sky130_fd_sc_hd__dfrtp_1
X_16276_ net372 _01950_ _01954_ _01912_ vssd1 vssd1 vccd1 vccd1 _01955_ sky130_fd_sc_hd__o211a_1
X_13488_ net225 _07906_ vssd1 vssd1 vccd1 vccd1 _07907_ sky130_fd_sc_hd__nor2_1
XFILLER_0_113_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18015_ net45 _03625_ vssd1 vssd1 vccd1 vccd1 _03626_ sky130_fd_sc_hd__nor2_1
X_12439_ net1094 _06631_ _07392_ _07399_ vssd1 vssd1 vccd1 vccd1 _07400_ sky130_fd_sc_hd__a211o_1
X_15227_ _05052_ net53 vssd1 vssd1 vccd1 vccd1 _01577_ sky130_fd_sc_hd__nor2_2
XFILLER_0_112_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14183__B2 net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15380__B1 _01594_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_114_3785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_3796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13930__B2 ag2.body\[65\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15158_ control.body\[858\] net102 _01569_ net2365 vssd1 vssd1 vccd1 vccd1 _00476_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_107_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11548__X _06521_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11941__B1 net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13476__A net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14109_ net997 ag2.body\[568\] vssd1 vssd1 vccd1 vccd1 _08270_ sky130_fd_sc_hd__or2_1
X_19966_ clknet_leaf_62_clk _00910_ net1469 vssd1 vssd1 vccd1 vccd1 ag2.body\[428\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_107_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15089_ control.body\[924\] net147 _01562_ net2388 vssd1 vssd1 vccd1 vccd1 _00414_
+ sky130_fd_sc_hd__a22o_1
Xfanout109 net110 vssd1 vssd1 vccd1 vccd1 net109 sky130_fd_sc_hd__buf_2
XANTENNA__20370__Q obsg2.obstacleArray\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18917_ clknet_leaf_142_clk img_gen.tracker.next_frame\[355\] net1253 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[355\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_43_1592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11267__Y _06240_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17890__B _03457_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19897_ clknet_leaf_85_clk _00841_ net1462 vssd1 vssd1 vccd1 vccd1 ag2.body\[503\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__16787__A net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14859__X _01530_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18903__CLK clknet_leaf_144_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09650_ net1073 control.body\[750\] vssd1 vssd1 vccd1 vccd1 _04623_ sky130_fd_sc_hd__nand2_1
XANTENNA__17424__A2 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20193__CLK clknet_leaf_88_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18848_ clknet_leaf_4_clk img_gen.tracker.next_frame\[286\] net1277 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[286\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_78_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09581_ net890 net896 vssd1 vssd1 vccd1 vccd1 _04554_ sky130_fd_sc_hd__and2b_2
X_18779_ clknet_leaf_17_clk img_gen.tracker.next_frame\[217\] net1285 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[217\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_77_402 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10050__D _05022_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14100__A net1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17889__Y _03529_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15199__B1 _01573_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout153_A net154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09688__X _04661_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18226__B net40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17768__D _03140_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19409__CLK clknet_leaf_103_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16148__C1 net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout418_A net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_30_clk clknet_4_4__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_30_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout1062_A net1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18152__A3 net37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16163__A2 net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16794__S0 net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09015_ ag2.body\[143\] vssd1 vssd1 vccd1 vccd1 _04040_ sky130_fd_sc_hd__inv_2
XANTENNA__15371__B1 _01593_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_297 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16461__S net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14770__A net1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18242__A _03683_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19559__CLK clknet_leaf_115_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13921__A1 ag2.body\[65\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold130 img_gen.tracker.frame\[248\] vssd1 vssd1 vccd1 vccd1 net1692 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13921__B2 ag2.body\[57\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold141 img_gen.tracker.frame\[433\] vssd1 vssd1 vccd1 vccd1 net1703 sky130_fd_sc_hd__dlygate4sd3_1
Xhold152 img_gen.tracker.frame\[554\] vssd1 vssd1 vccd1 vccd1 net1714 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12561__Y _07480_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout787_A net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold163 img_gen.tracker.frame\[335\] vssd1 vssd1 vccd1 vccd1 net1725 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold174 img_gen.tracker.frame\[419\] vssd1 vssd1 vccd1 vccd1 net1736 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_125_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09583__B _04471_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10362__X _05335_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold185 img_gen.tracker.frame\[230\] vssd1 vssd1 vccd1 vccd1 net1747 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__16320__C1 net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1115_X net1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold196 img_gen.tracker.frame\[443\] vssd1 vssd1 vccd1 vccd1 net1758 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout610 _06475_ vssd1 vssd1 vccd1 vccd1 net610 sky130_fd_sc_hd__buf_4
Xfanout621 net622 vssd1 vssd1 vccd1 vccd1 net621 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_61_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16871__B1 net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20106_ clknet_leaf_80_clk _01050_ net1487 vssd1 vssd1 vccd1 vccd1 ag2.body\[280\]
+ sky130_fd_sc_hd__dfrtp_4
Xfanout632 _06462_ vssd1 vssd1 vccd1 vccd1 net632 sky130_fd_sc_hd__buf_2
X_09917_ ag2.body\[315\] net772 net776 ag2.body\[314\] vssd1 vssd1 vccd1 vccd1 _04890_
+ sky130_fd_sc_hd__a2bb2o_1
Xfanout643 _04417_ vssd1 vssd1 vccd1 vccd1 net643 sky130_fd_sc_hd__buf_4
XANTENNA__12488__A1 net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout954_A net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout654 _04394_ vssd1 vssd1 vccd1 vccd1 net654 sky130_fd_sc_hd__buf_2
XANTENNA_fanout575_X net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18583__CLK clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout665 net666 vssd1 vssd1 vccd1 vccd1 net665 sky130_fd_sc_hd__dlymetal6s2s_1
Xclkbuf_leaf_97_clk clknet_4_11__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_97_clk
+ sky130_fd_sc_hd__clkbuf_8
Xfanout676 net677 vssd1 vssd1 vccd1 vccd1 net676 sky130_fd_sc_hd__clkbuf_4
X_20037_ clknet_leaf_67_clk _00981_ net1494 vssd1 vssd1 vccd1 vccd1 ag2.body\[355\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__17415__A2 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout687 _04390_ vssd1 vssd1 vccd1 vccd1 net687 sky130_fd_sc_hd__clkbuf_4
X_09848_ net1087 control.body\[974\] vssd1 vssd1 vccd1 vccd1 _04821_ sky130_fd_sc_hd__xor2_1
Xfanout698 _04268_ vssd1 vssd1 vccd1 vccd1 net698 sky130_fd_sc_hd__buf_4
XFILLER_0_38_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout66_A net67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_4092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17305__B net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout742_X net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09779_ _04743_ _04744_ _04747_ _04751_ vssd1 vssd1 vccd1 vccd1 _04752_ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout1484_X net1484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12425__B1_N _06505_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11810_ img_gen.tracker.frame\[461\] net597 vssd1 vssd1 vccd1 vccd1 _06782_ sky130_fd_sc_hd__or2_1
X_12790_ net336 net332 _07497_ vssd1 vssd1 vccd1 vccd1 _07598_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_1_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11741_ img_gen.tracker.frame\[17\] net606 net551 img_gen.tracker.frame\[20\] _06712_
+ vssd1 vssd1 vccd1 vccd1 _06713_ sky130_fd_sc_hd__o221a_1
XFILLER_0_68_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11463__A2 net1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12660__A1 net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16636__S net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15729__A2 net200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_427 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10671__B1 _05634_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14460_ net972 ag2.body\[435\] vssd1 vssd1 vccd1 vccd1 _08621_ sky130_fd_sc_hd__xor2_1
X_11672_ net1094 net1070 _06643_ vssd1 vssd1 vccd1 vccd1 _06644_ sky130_fd_sc_hd__o21a_2
XANTENNA__18128__B1 net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08943__A net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_137_4497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13411_ net671 _07876_ vssd1 vssd1 vccd1 vccd1 _07877_ sky130_fd_sc_hd__nor2_1
X_10623_ ag2.body\[48\] net1223 vssd1 vssd1 vccd1 vccd1 _05596_ sky130_fd_sc_hd__nand2_1
X_14391_ _08544_ _08546_ _08549_ _08551_ vssd1 vssd1 vccd1 vccd1 _08552_ sky130_fd_sc_hd__or4b_1
XANTENNA__09758__B net1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_21_clk clknet_4_6__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_21_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_88_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16130_ obsg2.obstacleArray\[72\] obsg2.obstacleArray\[73\] net425 vssd1 vssd1 vccd1
+ vccd1 _01809_ sky130_fd_sc_hd__mux2_1
X_13342_ _07512_ net304 vssd1 vssd1 vccd1 vccd1 _07850_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_42_1589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10554_ _05510_ _05511_ _05518_ _05519_ vssd1 vssd1 vccd1 vccd1 _05527_ sky130_fd_sc_hd__a22o_1
XANTENNA__17975__B net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16154__A2 net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20066__CLK clknet_leaf_73_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1079 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16061_ _01726_ _01738_ vssd1 vssd1 vccd1 vccd1 _01740_ sky130_fd_sc_hd__or2_1
XANTENNA__15776__A _05798_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15362__B1 _01592_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13273_ net385 _07460_ _07813_ vssd1 vssd1 vccd1 vccd1 _07823_ sky130_fd_sc_hd__and3_1
XFILLER_0_121_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10485_ _04215_ net1150 net754 ag2.body\[589\] _05455_ vssd1 vssd1 vccd1 vccd1 _05458_
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_121_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13912__A1 ag2.body\[57\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12224_ img_gen.updater.commands.count\[12\] img_gen.updater.commands.count\[7\]
+ _07192_ _07193_ img_gen.updater.commands.count\[13\] vssd1 vssd1 vccd1 vccd1 _07194_
+ sky130_fd_sc_hd__o311a_1
X_15012_ control.body\[984\] net166 _01553_ net2556 vssd1 vssd1 vccd1 vccd1 _00346_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_126_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12912__B _07460_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11368__X _06341_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19820_ clknet_leaf_89_clk _00764_ net1411 vssd1 vssd1 vccd1 vccd1 ag2.body\[570\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__09493__B net1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15114__B1 _01554_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_766 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12155_ img_gen.tracker.frame\[477\] net578 net573 vssd1 vssd1 vccd1 vccd1 _07127_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_130_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16311__C1 net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11106_ net1160 control.body\[1099\] vssd1 vssd1 vccd1 vccd1 _06079_ sky130_fd_sc_hd__nor2_1
X_19751_ clknet_leaf_130_clk _00695_ net1317 vssd1 vssd1 vccd1 vccd1 control.body\[645\]
+ sky130_fd_sc_hd__dfrtp_1
X_16963_ _02635_ _02637_ _02641_ _02636_ vssd1 vssd1 vccd1 vccd1 _02642_ sky130_fd_sc_hd__or4b_4
XFILLER_0_75_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12086_ net565 _07057_ _07055_ net474 vssd1 vssd1 vccd1 vccd1 _07058_ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_88_clk clknet_4_12__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_88_clk
+ sky130_fd_sc_hd__clkbuf_8
X_18702_ clknet_leaf_10_clk img_gen.tracker.next_frame\[140\] net1274 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[140\] sky130_fd_sc_hd__dfrtp_1
X_15914_ ag2.body\[187\] net131 _01652_ ag2.body\[179\] vssd1 vssd1 vccd1 vccd1 _01149_
+ sky130_fd_sc_hd__a22o_1
X_11037_ net1111 control.body\[1045\] vssd1 vssd1 vccd1 vccd1 _06010_ sky130_fd_sc_hd__nand2b_1
X_19682_ clknet_leaf_117_clk _00626_ net1384 vssd1 vssd1 vccd1 vccd1 control.body\[704\]
+ sky130_fd_sc_hd__dfrtp_1
X_16894_ ag2.body\[209\] net874 vssd1 vssd1 vccd1 vccd1 _02573_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_95_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18633_ clknet_leaf_0_clk img_gen.tracker.next_frame\[71\] net1242 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[71\] sky130_fd_sc_hd__dfrtp_1
X_15845_ ag2.body\[254\] net181 _01644_ ag2.body\[246\] vssd1 vssd1 vccd1 vccd1 _01088_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_91_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_3453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18564_ clknet_leaf_15_clk img_gen.tracker.next_frame\[2\] net1278 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[2\] sky130_fd_sc_hd__dfrtp_1
X_15776_ _05798_ net60 vssd1 vssd1 vccd1 vccd1 _01638_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_103_3464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12100__B1 net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12988_ img_gen.tracker.frame\[256\] net645 vssd1 vssd1 vccd1 vccd1 _07690_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_103_3475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17515_ _04213_ net868 net858 _04214_ _03190_ vssd1 vssd1 vccd1 vccd1 _03194_ sky130_fd_sc_hd__a221o_1
X_14727_ net1041 ag2.body\[116\] vssd1 vssd1 vccd1 vccd1 _08888_ sky130_fd_sc_hd__xor2_1
XFILLER_0_87_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18495_ net1516 net1510 vssd1 vssd1 vccd1 vccd1 _00026_ sky130_fd_sc_hd__or2_1
X_11939_ img_gen.tracker.frame\[154\] net587 net548 img_gen.tracker.frame\[151\] _06910_
+ vssd1 vssd1 vccd1 vccd1 _06911_ sky130_fd_sc_hd__o221a_1
XANTENNA__12651__A1 net242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11454__A2 _06412_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17446_ ag2.body\[382\] net940 vssd1 vssd1 vccd1 vccd1 _03125_ sky130_fd_sc_hd__xor2_1
XANTENNA__14928__B1 _01543_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14658_ _08813_ _08815_ _08817_ _08818_ vssd1 vssd1 vccd1 vccd1 _08819_ sky130_fd_sc_hd__or4bb_2
XFILLER_0_28_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17590__A1 ag2.body\[59\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18046__B _03558_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13609_ control.divider.count\[1\] control.divider.count\[0\] control.divider.count\[2\]
+ vssd1 vssd1 vccd1 vccd1 _07982_ sky130_fd_sc_hd__a21o_1
XANTENNA__11206__A2 _06163_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17377_ _03049_ _03050_ _03053_ _03055_ _03005_ vssd1 vssd1 vccd1 vccd1 _03056_ sky130_fd_sc_hd__o2111a_1
XANTENNA__09668__B _04640_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14589_ net1004 _04011_ ag2.body\[81\] _03965_ _08744_ vssd1 vssd1 vccd1 vccd1 _08750_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_83_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_12_clk clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_12_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_116_3847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12806__C net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19116_ clknet_leaf_141_clk img_gen.tracker.next_frame\[554\] net1262 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[554\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_116_3858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16328_ obsg2.obstacleArray\[74\] obsg2.obstacleArray\[75\] net406 vssd1 vssd1 vccd1
+ vccd1 _02007_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_116_3869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12094__B net1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_1611 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19047_ clknet_leaf_8_clk img_gen.tracker.next_frame\[485\] net1273 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[485\] sky130_fd_sc_hd__dfrtp_1
X_16259_ net371 _01933_ _01937_ _01912_ vssd1 vssd1 vccd1 vccd1 _01938_ sky130_fd_sc_hd__o211a_1
XANTENNA__16281__S net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12662__X _07536_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12167__B1 net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_768 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_267 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_1210 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19851__CLK clknet_leaf_93_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_71_2475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_2486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19949_ clknet_leaf_45_clk _00893_ net1379 vssd1 vssd1 vccd1 vccd1 ag2.body\[443\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_71_2497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_79_clk clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_79_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_96_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09702_ ag2.body\[70\] net1089 vssd1 vssd1 vccd1 vccd1 _04675_ sky130_fd_sc_hd__xor2_1
XFILLER_0_4_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10910__X _05883_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16605__B1 net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09633_ net917 _04599_ _04601_ _04605_ vssd1 vssd1 vccd1 vccd1 _04606_ sky130_fd_sc_hd__o31a_2
XANTENNA__11693__A2 net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12890__A1 net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17125__B net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_88_2994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10350__C1 _04418_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09564_ net920 _04239_ vssd1 vssd1 vccd1 vccd1 _04537_ sky130_fd_sc_hd__or2_1
XANTENNA__13372__C _07813_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16964__B net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19231__CLK clknet_leaf_75_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09495_ _04464_ _04465_ _04466_ _04467_ vssd1 vssd1 vccd1 vccd1 _04468_ sky130_fd_sc_hd__or4_1
XANTENNA__14765__A net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18237__A net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17030__B1 net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1277_A net1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_1383 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1214 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16028__Y _01707_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17581__B2 ag2.body\[339\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14395__A1 net993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14395__B2 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout702_A _04268_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11828__S0 net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1065_X net1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1444_A net1452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_994 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_4350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_22_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17795__B _03468_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_132_4361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16136__A2 net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20586_ clknet_leaf_105_clk net2301 _00050_ vssd1 vssd1 vccd1 vccd1 sound_gen.posDetector1.N\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_6_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09810__A2 _04723_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18949__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15344__B1 _01590_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1232_X net1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17884__A2 _04445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10270_ ag2.body\[143\] net1065 vssd1 vssd1 vccd1 vccd1 _05243_ sky130_fd_sc_hd__xor2_1
XFILLER_0_14_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout692_X net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11905__B1 net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12732__B _07444_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17097__B1 obsg2.randCord\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14005__A net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1405 net1409 vssd1 vssd1 vccd1 vccd1 net1405 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11348__B net1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1416 net1419 vssd1 vssd1 vccd1 vccd1 net1416 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_54_1961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1427 net1430 vssd1 vssd1 vccd1 vccd1 net1427 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_126_4154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout440 _06645_ vssd1 vssd1 vccd1 vccd1 net440 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_54_1972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout957_X net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_126_4165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1438 net1439 vssd1 vssd1 vccd1 vccd1 net1438 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_54_1983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout451 _02213_ vssd1 vssd1 vccd1 vccd1 net451 sky130_fd_sc_hd__buf_4
Xfanout1449 net1451 vssd1 vssd1 vccd1 vccd1 net1449 sky130_fd_sc_hd__clkbuf_4
Xfanout462 net463 vssd1 vssd1 vccd1 vccd1 net462 sky130_fd_sc_hd__buf_2
XFILLER_0_22_1473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_35_1382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_4029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13960_ ag2.body\[100\] net189 _08156_ ag2.body\[92\] vssd1 vssd1 vccd1 vccd1 _00181_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_35_1393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout473 _06647_ vssd1 vssd1 vccd1 vccd1 net473 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_50_1847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout484 _02373_ vssd1 vssd1 vccd1 vccd1 net484 sky130_fd_sc_hd__buf_4
XANTENNA__08938__A net1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout495 net496 vssd1 vssd1 vccd1 vccd1 net495 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_6_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14870__A2 net182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12911_ net2048 net661 _07315_ _07653_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[215\]
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_57_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17035__B net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13891_ ag2.body\[39\] net115 _08148_ ag2.body\[31\] vssd1 vssd1 vccd1 vccd1 _00120_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11684__A2 net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16072__A1 net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15630_ ag2.body\[446\] net127 _01621_ ag2.body\[438\] vssd1 vssd1 vccd1 vccd1 _00896_
+ sky130_fd_sc_hd__a22o_1
X_12842_ net676 _07622_ vssd1 vssd1 vccd1 vccd1 _07623_ sky130_fd_sc_hd__nor2_1
XANTENNA__11083__B net1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15561_ ag2.body\[496\] net185 _01614_ ag2.body\[488\] vssd1 vssd1 vccd1 vccd1 _00834_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_96_563 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12773_ net338 net333 net312 _07486_ vssd1 vssd1 vccd1 vccd1 _07590_ sky130_fd_sc_hd__or4_1
XFILLER_0_115_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08944__Y _03969_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17300_ ag2.body\[344\] net739 net944 _04124_ vssd1 vssd1 vccd1 vccd1 _02979_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_96_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_1776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14512_ _08670_ _08671_ _08672_ vssd1 vssd1 vccd1 vccd1 _08673_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_48_1787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18280_ net298 _03549_ _03564_ _03579_ obsg2.obstacleArray\[137\] vssd1 vssd1 vccd1
+ vccd1 _03779_ sky130_fd_sc_hd__a41o_1
XTAP_TAPCELL_ROW_48_1798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11724_ img_gen.tracker.frame\[230\] net624 net577 _06695_ vssd1 vssd1 vccd1 vccd1
+ _06696_ sky130_fd_sc_hd__o211a_1
X_15492_ ag2.body\[563\] net109 _01606_ ag2.body\[555\] vssd1 vssd1 vccd1 vccd1 _00773_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_132_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17231_ ag2.body\[441\] net732 net851 _04157_ _02908_ vssd1 vssd1 vccd1 vccd1 _02910_
+ sky130_fd_sc_hd__a221o_1
XANTENNA__14386__A1 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17986__A net46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14386__B2 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11655_ net1118 net1070 vssd1 vssd1 vccd1 vccd1 _06628_ sky130_fd_sc_hd__nand2_1
X_14443_ net1030 ag2.body\[229\] vssd1 vssd1 vccd1 vccd1 _08604_ sky130_fd_sc_hd__nand2_1
XFILLER_0_126_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09488__B net1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout80 net83 vssd1 vssd1 vccd1 vccd1 net80 sky130_fd_sc_hd__buf_2
XFILLER_0_68_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12626__C net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout91 net219 vssd1 vssd1 vccd1 vccd1 net91 sky130_fd_sc_hd__clkbuf_2
X_10606_ net1060 control.body\[991\] vssd1 vssd1 vccd1 vccd1 _05579_ sky130_fd_sc_hd__or2_1
X_17162_ ag2.body\[596\] net959 vssd1 vssd1 vccd1 vccd1 _02841_ sky130_fd_sc_hd__xor2_1
XFILLER_0_64_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14374_ net973 ag2.body\[419\] vssd1 vssd1 vccd1 vccd1 _08535_ sky130_fd_sc_hd__or2_1
XFILLER_0_4_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11586_ _06472_ _06558_ vssd1 vssd1 vccd1 vccd1 _06559_ sky130_fd_sc_hd__or2_1
XFILLER_0_29_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16113_ _01790_ _01791_ net374 vssd1 vssd1 vccd1 vccd1 _01792_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_111_3700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_3176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13325_ net251 _07842_ _07843_ net1846 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[439\]
+ sky130_fd_sc_hd__a22o_1
X_10537_ ag2.body\[229\] net1111 vssd1 vssd1 vccd1 vccd1 _05510_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_111_3711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_3187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17093_ ag2.body\[297\] net875 vssd1 vssd1 vccd1 vccd1 _02772_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_94_3198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_3722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16044_ _01721_ _01722_ vssd1 vssd1 vccd1 vccd1 _01723_ sky130_fd_sc_hd__nor2_1
X_10468_ net1059 control.body\[1015\] vssd1 vssd1 vccd1 vccd1 _05441_ sky130_fd_sc_hd__or2_1
X_13256_ net257 _07815_ _07816_ net1665 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[397\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_126_1276 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12207_ img_gen.control.detect4.Q\[1\] img_gen.control.detect4.Q\[0\] vssd1 vssd1
+ vccd1 vccd1 _07179_ sky130_fd_sc_hd__nand2b_1
XANTENNA__18032__D net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17627__A2 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13187_ net241 _07783_ _07784_ net1777 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[360\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__10443__A net1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10399_ net1086 control.body\[1062\] vssd1 vssd1 vccd1 vccd1 _05372_ sky130_fd_sc_hd__xor2_1
XANTENNA__19104__CLK clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19803_ clknet_leaf_124_clk _00747_ net1405 vssd1 vssd1 vccd1 vccd1 ag2.body\[585\]
+ sky130_fd_sc_hd__dfrtp_2
X_12138_ img_gen.tracker.frame\[501\] net583 net547 img_gen.tracker.frame\[498\] _07109_
+ vssd1 vssd1 vccd1 vccd1 _07110_ sky130_fd_sc_hd__o221a_1
XFILLER_0_97_1316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17995_ net352 _03610_ vssd1 vssd1 vccd1 vccd1 _03611_ sky130_fd_sc_hd__or2_1
XANTENNA__10162__B net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_109_3640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_3651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16946_ ag2.body\[386\] net862 vssd1 vssd1 vccd1 vccd1 _02625_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_109_3662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12069_ img_gen.tracker.frame\[108\] net629 net611 img_gen.tracker.frame\[111\] _07040_
+ vssd1 vssd1 vccd1 vccd1 _07041_ sky130_fd_sc_hd__a221o_1
X_19734_ clknet_leaf_129_clk _00678_ net1325 vssd1 vssd1 vccd1 vccd1 control.body\[660\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10730__X _05703_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_1_clk clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_1_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_105_3515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14861__A2 _08521_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19225__RESET_B net1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_3526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_3537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18052__A2 _03566_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19665_ clknet_leaf_119_clk _00609_ net1391 vssd1 vssd1 vccd1 vccd1 control.body\[735\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__19254__CLK clknet_leaf_75_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16599__C1 net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16877_ _02550_ _02551_ _02553_ _02555_ vssd1 vssd1 vccd1 vccd1 _02556_ sky130_fd_sc_hd__or4_1
XANTENNA__12872__A1 net245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11274__A ag2.body\[122\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18616_ clknet_leaf_144_clk img_gen.tracker.next_frame\[54\] net1242 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[54\] sky130_fd_sc_hd__dfrtp_1
X_15828_ ag2.body\[270\] net205 _01643_ ag2.body\[262\] vssd1 vssd1 vccd1 vccd1 _01072_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_126_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19596_ clknet_leaf_118_clk _00540_ net1392 vssd1 vssd1 vccd1 vccd1 control.body\[794\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_133_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_1079 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__20231__CLK clknet_leaf_66_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18547_ clknet_leaf_137_clk _00073_ net1299 vssd1 vssd1 vccd1 vccd1 img_gen.updater.commands.count\[16\]
+ sky130_fd_sc_hd__dfrtp_2
X_15759_ ag2.body\[320\] net215 _01636_ ag2.body\[312\] vssd1 vssd1 vccd1 vccd1 _01010_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12624__A1 net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14585__A net1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_120 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18057__A net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17012__B1 net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09280_ sound_gen.osc1.stayCount\[23\] _04287_ _04301_ _04302_ vssd1 vssd1 vccd1
+ vccd1 _04303_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_118_3909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18478_ net1512 net1506 vssd1 vssd1 vccd1 vccd1 _00009_ sky130_fd_sc_hd__or2_1
XFILLER_0_30_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_64_2290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16366__A2 net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_2143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_2154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17429_ ag2.body\[116\] net714 net708 ag2.body\[117\] vssd1 vssd1 vccd1 vccd1 _03108_
+ sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_60_2165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20440_ clknet_leaf_26_clk _01327_ net1343 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[76\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_71_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10337__B net1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14129__A1 net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1029 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20371_ clknet_leaf_23_clk _01258_ net1360 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[7\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_77_2662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_2673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload50 clknet_leaf_32_clk vssd1 vssd1 vccd1 vccd1 clkload50/Y sky130_fd_sc_hd__inv_16
XTAP_TAPCELL_ROW_77_2684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload61 clknet_leaf_50_clk vssd1 vssd1 vccd1 vccd1 clkload61/Y sky130_fd_sc_hd__inv_12
XTAP_TAPCELL_ROW_73_2537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload72 clknet_leaf_113_clk vssd1 vssd1 vccd1 vccd1 clkload72/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_3_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_58_2083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_1331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_73_2548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload83 clknet_leaf_124_clk vssd1 vssd1 vccd1 vccd1 clkload83/X sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_58_2094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload94 clknet_leaf_112_clk vssd1 vssd1 vccd1 vccd1 clkload94/Y sky130_fd_sc_hd__clkinv_2
XFILLER_0_62_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11449__A net1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17618__A2 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13367__C _07532_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1025_A net1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18520__A net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16959__B net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08995_ ag2.body\[93\] vssd1 vssd1 vccd1 vccd1 _04020_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout485_A _02373_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14837__C1 _08904_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13664__A net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09861__B net1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14301__B2 net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09859__A2 _04238_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12863__A1 net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10800__B net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1394_A net1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09616_ net1099 control.body\[805\] vssd1 vssd1 vccd1 vccd1 _04589_ sky130_fd_sc_hd__xor2_1
XFILLER_0_116_1423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14065__B1 _08225_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15801__A1 ag2.body\[294\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16694__B net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09547_ net896 _04519_ net636 vssd1 vssd1 vccd1 vccd1 _04520_ sky130_fd_sc_hd__a21oi_4
XANTENNA_fanout440_X net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16186__S net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14495__A net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12567__X _07483_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout538_X net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1182_X net1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17003__B1 net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09589__A net1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_4570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_4401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09478_ ag2.body\[468\] net1128 vssd1 vssd1 vccd1 vccd1 _04451_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_134_4412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_4423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12727__B _07567_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14368__A1 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_1518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_1640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14368__B2 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_123 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout705_X net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18530__RESET_B net1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload0 clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clkload0/X sky130_fd_sc_hd__clkbuf_8
X_11440_ _04424_ _04550_ _04772_ vssd1 vssd1 vccd1 vccd1 _06413_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_62_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20638_ net1555 vssd1 vssd1 vccd1 vccd1 gpio_out[33] sky130_fd_sc_hd__buf_2
XANTENNA__15597__Y _01619_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16109__A2 net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10247__B net1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10929__A1 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11051__B1 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11371_ ag2.body\[479\] net1057 vssd1 vssd1 vccd1 vccd1 _06344_ sky130_fd_sc_hd__xor2_1
XFILLER_0_11_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20569_ clknet_leaf_107_clk net1590 _00033_ vssd1 vssd1 vccd1 vccd1 sound_gen.dac1.dacCount\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_10322_ ag2.body\[608\] net1219 vssd1 vssd1 vccd1 vccd1 _05295_ sky130_fd_sc_hd__xor2_1
X_13110_ net284 _07745_ _07746_ net1972 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[320\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_104_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14090_ net1031 ag2.body\[285\] vssd1 vssd1 vccd1 vccd1 _08251_ sky130_fd_sc_hd__nand2_1
XFILLER_0_46_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1139 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_128_4216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13041_ _07715_ net254 _07713_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[283\]
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_128_4227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10253_ control.body\[788\] net1130 vssd1 vssd1 vccd1 vccd1 _05226_ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_128_4238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10157__A2 net1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16817__B1 net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16869__B net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11078__B net1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10184_ _05153_ _05154_ _05155_ _05156_ vssd1 vssd1 vccd1 vccd1 _05157_ sky130_fd_sc_hd__a22o_1
Xfanout1202 net1203 vssd1 vssd1 vccd1 vccd1 net1202 sky130_fd_sc_hd__buf_4
Xfanout1213 net1214 vssd1 vssd1 vccd1 vccd1 net1213 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_33_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1224 net1225 vssd1 vssd1 vccd1 vccd1 net1224 sky130_fd_sc_hd__clkbuf_8
Xfanout1235 net1238 vssd1 vssd1 vccd1 vccd1 net1235 sky130_fd_sc_hd__buf_4
X_16800_ net365 net363 _02478_ vssd1 vssd1 vccd1 vccd1 _02479_ sky130_fd_sc_hd__and3_1
Xfanout1246 net1250 vssd1 vssd1 vccd1 vccd1 net1246 sky130_fd_sc_hd__clkbuf_4
X_17780_ obsg2.obsNeeded\[0\] _04399_ _03458_ vssd1 vssd1 vccd1 vccd1 _03459_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_22_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09771__B net1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1257 net1263 vssd1 vssd1 vccd1 vccd1 net1257 sky130_fd_sc_hd__clkbuf_4
X_14992_ net2203 net158 _01549_ control.body\[1007\] vssd1 vssd1 vccd1 vccd1 _00329_
+ sky130_fd_sc_hd__a22o_1
Xfanout270 _04307_ vssd1 vssd1 vccd1 vccd1 net270 sky130_fd_sc_hd__buf_2
Xfanout1268 net1269 vssd1 vssd1 vccd1 vccd1 net1268 sky130_fd_sc_hd__clkbuf_4
Xfanout1279 net1280 vssd1 vssd1 vccd1 vccd1 net1279 sky130_fd_sc_hd__clkbuf_2
Xfanout281 net282 vssd1 vssd1 vccd1 vccd1 net281 sky130_fd_sc_hd__clkbuf_4
X_16731_ obsg2.obstacleArray\[99\] net500 net481 obsg2.obstacleArray\[97\] vssd1 vssd1
+ vccd1 vccd1 _02410_ sky130_fd_sc_hd__a22o_1
Xfanout292 net293 vssd1 vssd1 vccd1 vccd1 net292 sky130_fd_sc_hd__clkbuf_4
X_13943_ ag2.body\[85\] net197 _08154_ ag2.body\[77\] vssd1 vssd1 vccd1 vccd1 _00166_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11806__B net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14957__X _01547_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19450_ clknet_leaf_110_clk _00394_ net1416 vssd1 vssd1 vccd1 vccd1 control.body\[936\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__17242__B1 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16662_ _02336_ _02337_ _02340_ net359 net357 vssd1 vssd1 vccd1 vccd1 _02341_ sky130_fd_sc_hd__o221a_1
XFILLER_0_72_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13874_ _04903_ net56 vssd1 vssd1 vccd1 vccd1 _08147_ sky130_fd_sc_hd__nor2_2
XANTENNA__17793__A1 net1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16596__A2 net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18401_ _08139_ _03826_ vssd1 vssd1 vccd1 vccd1 _03891_ sky130_fd_sc_hd__nand2_1
X_15613_ ag2.body\[462\] net123 _01620_ ag2.body\[454\] vssd1 vssd1 vccd1 vccd1 _00880_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12606__A1 net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12825_ net240 _07613_ _07614_ net1759 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[168\]
+ sky130_fd_sc_hd__a22o_1
X_19381_ clknet_leaf_112_clk _00325_ net1425 vssd1 vssd1 vccd1 vccd1 control.body\[1011\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12067__C1 net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16593_ obsg2.obstacleArray\[72\] obsg2.obstacleArray\[73\] net443 vssd1 vssd1 vccd1
+ vccd1 _02272_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10617__B1 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18332_ net906 _04641_ _06173_ _08027_ _08140_ vssd1 vssd1 vccd1 vccd1 _03828_ sky130_fd_sc_hd__a311o_1
X_15544_ ag2.body\[514\] net187 _01580_ ag2.body\[506\] vssd1 vssd1 vccd1 vccd1 _00820_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12082__A2 net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12756_ net305 _07581_ vssd1 vssd1 vccd1 vccd1 _07582_ sky130_fd_sc_hd__nor2_1
XFILLER_0_84_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18263_ net530 _03770_ vssd1 vssd1 vccd1 vccd1 _01379_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_13_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11707_ img_gen.tracker.frame\[290\] net624 net607 img_gen.tracker.frame\[293\] vssd1
+ vssd1 vccd1 vccd1 _06679_ sky130_fd_sc_hd__o22a_1
XFILLER_0_127_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15475_ ag2.body\[580\] net111 _01604_ ag2.body\[572\] vssd1 vssd1 vccd1 vccd1 _00758_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_96_3238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12687_ net388 net384 net382 _07306_ vssd1 vssd1 vccd1 vccd1 _07549_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_96_3249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17214_ ag2.body\[50\] net722 net929 _03994_ _02889_ vssd1 vssd1 vccd1 vccd1 _02893_
+ sky130_fd_sc_hd__a221o_1
X_14426_ net980 ag2.body\[554\] vssd1 vssd1 vccd1 vccd1 _08587_ sky130_fd_sc_hd__xor2_1
XFILLER_0_65_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18194_ _01703_ _03638_ _03703_ vssd1 vssd1 vccd1 vccd1 _03736_ sky130_fd_sc_hd__and3_1
X_11638_ _06511_ _06571_ _06584_ _06529_ vssd1 vssd1 vccd1 vccd1 _06611_ sky130_fd_sc_hd__a31o_1
XFILLER_0_21_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_1327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17145_ _02820_ _02821_ _02822_ _02823_ vssd1 vssd1 vccd1 vccd1 _02824_ sky130_fd_sc_hd__or4_1
XFILLER_0_68_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14357_ net977 _04144_ _04147_ net1013 vssd1 vssd1 vccd1 vccd1 _08518_ sky130_fd_sc_hd__a22o_1
XFILLER_0_107_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10263__A2_N _05222_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_1473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11569_ obsg2.obstacleArray\[88\] obsg2.obstacleArray\[89\] obsg2.obstacleArray\[92\]
+ obsg2.obstacleArray\[93\] net1125 net512 vssd1 vssd1 vccd1 vccd1 _06542_ sky130_fd_sc_hd__mux4_1
XFILLER_0_97_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold707 control.body\[922\] vssd1 vssd1 vccd1 vccd1 net2269 sky130_fd_sc_hd__dlygate4sd3_1
Xhold718 _00382_ vssd1 vssd1 vccd1 vccd1 net2280 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13308_ net384 net338 net331 _07486_ vssd1 vssd1 vccd1 vccd1 _07837_ sky130_fd_sc_hd__or4_2
X_17076_ _02747_ _02752_ _02753_ _02754_ vssd1 vssd1 vccd1 vccd1 _02755_ sky130_fd_sc_hd__or4_1
Xhold729 control.body\[936\] vssd1 vssd1 vccd1 vccd1 net2291 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14288_ net988 ag2.body\[473\] vssd1 vssd1 vccd1 vccd1 _08449_ sky130_fd_sc_hd__xor2_1
XANTENNA__09538__A1 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16027_ _01689_ _01704_ vssd1 vssd1 vccd1 vccd1 _01706_ sky130_fd_sc_hd__nand2_1
XFILLER_0_106_1647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_872 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13239_ net238 _07808_ _07809_ net1909 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[387\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__17508__X _03187_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16808__B1 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16284__A1 net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_127_Right_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17978_ obsg2.obstacleArray\[14\] _03599_ net522 vssd1 vssd1 vccd1 vccd1 _01265_
+ sky130_fd_sc_hd__o21a_1
XANTENNA__10901__A net1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13098__A1 net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18644__CLK clknet_leaf_15_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16929_ ag2.body\[369\] net733 net724 ag2.body\[370\] vssd1 vssd1 vccd1 vccd1 _02608_
+ sky130_fd_sc_hd__o22a_1
X_19717_ clknet_leaf_134_clk net2442 net1303 vssd1 vssd1 vccd1 vccd1 control.body\[675\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12845__A1 net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_2920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10620__B net1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17233__B1 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_2330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19648_ clknet_leaf_128_clk _00592_ net1329 vssd1 vssd1 vccd1 vccd1 control.body\[750\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_66_2341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_2806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09401_ net273 _04343_ _04384_ vssd1 vssd1 vccd1 vccd1 _01402_ sky130_fd_sc_hd__nor3_1
XFILLER_0_137_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14598__A1 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_2205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14598__B2 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18794__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19579_ clknet_leaf_117_clk _00523_ net1386 vssd1 vssd1 vccd1 vccd1 control.body\[809\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_62_2216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17403__B net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_2227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09332_ net2122 _04335_ vssd1 vssd1 vccd1 vccd1 _01430_ sky130_fd_sc_hd__xor2_1
XANTENNA__17897__Y _03533_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09474__B1 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13270__A1 net236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12073__A2 net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_1331 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09263_ _04287_ vssd1 vssd1 vccd1 vccd1 sound_gen.osc1.timer_nxt\[12\] sky130_fd_sc_hd__inv_2
XANTENNA__09202__A net1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout233_A net247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11820__A2 net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_2724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_2735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_1386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_2746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13022__A1 net240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09194_ ag2.body\[602\] vssd1 vssd1 vccd1 vccd1 _04219_ sky130_fd_sc_hd__inv_2
XFILLER_0_117_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18234__B net35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13659__A net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20423_ clknet_leaf_37_clk _01310_ net1350 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[59\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_47_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14107__X _08268_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12563__A net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16035__A net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1415 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1142_A net1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20354_ clknet_leaf_140_clk _01245_ net1291 vssd1 vssd1 vccd1 vccd1 img_gen.updater.commands.rR1.rainbowRNG\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_105_1135 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20285_ clknet_leaf_35_clk control.divider.next_count\[6\] net1348 vssd1 vssd1 vccd1
+ vccd1 control.divider.count\[6\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_101_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18250__A _03691_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1028_X net1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19147__RESET_B net1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout390_X net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17698__S1 net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11887__A2 net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout488_X net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16275__A1 net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold12 control.button2.Q\[1\] vssd1 vssd1 vccd1 vccd1 net1574 sky130_fd_sc_hd__dlygate4sd3_1
Xhold23 control.button4.Q\[0\] vssd1 vssd1 vccd1 vccd1 net1585 sky130_fd_sc_hd__dlygate4sd3_1
X_08978_ ag2.body\[72\] vssd1 vssd1 vccd1 vccd1 _04003_ sky130_fd_sc_hd__inv_2
XANTENNA__10811__A net1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold34 img_gen.tracker.frame\[8\] vssd1 vssd1 vccd1 vccd1 net1596 sky130_fd_sc_hd__dlygate4sd3_1
Xhold45 img_gen.tracker.frame\[543\] vssd1 vssd1 vccd1 vccd1 net1607 sky130_fd_sc_hd__dlygate4sd3_1
Xhold56 img_gen.tracker.frame\[407\] vssd1 vssd1 vccd1 vccd1 net1618 sky130_fd_sc_hd__dlygate4sd3_1
Xhold67 _01207_ vssd1 vssd1 vccd1 vccd1 net1629 sky130_fd_sc_hd__dlygate4sd3_1
Xhold78 img_gen.tracker.frame\[522\] vssd1 vssd1 vccd1 vccd1 net1640 sky130_fd_sc_hd__dlygate4sd3_1
Xhold89 img_gen.tracker.frame\[492\] vssd1 vssd1 vccd1 vccd1 net1651 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__17224__B1 net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10940_ ag2.body\[296\] net1237 vssd1 vssd1 vccd1 vccd1 _05913_ sky130_fd_sc_hd__xor2_1
XFILLER_0_98_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14589__A1 net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13841__B net223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14589__B2 _03965_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout822_X net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10871_ _05840_ _05841_ _05842_ _05843_ vssd1 vssd1 vccd1 vccd1 _05844_ sky130_fd_sc_hd__a22o_1
XANTENNA__12738__A net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12610_ net231 _07506_ _07507_ net1832 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[60\]
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_26_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13590_ _07953_ _07964_ _07963_ vssd1 vssd1 vccd1 vccd1 _07965_ sky130_fd_sc_hd__o21a_1
XANTENNA__09465__B1 net1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13261__A1 net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_26_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14027__A1_N net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12541_ net313 _07468_ vssd1 vssd1 vccd1 vccd1 _07469_ sky130_fd_sc_hd__or2_1
XFILLER_0_137_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_4_6__f_clk_X clknet_4_6__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13013__A1 net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15260_ net2621 net97 net50 net2213 vssd1 vssd1 vccd1 vccd1 _00568_ sky130_fd_sc_hd__a22o_1
X_12472_ net385 net382 _07306_ _06724_ vssd1 vssd1 vccd1 vccd1 _07427_ sky130_fd_sc_hd__a31o_1
XFILLER_0_129_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16750__A2 net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14211_ net1000 ag2.body\[408\] vssd1 vssd1 vccd1 vccd1 _08372_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_91_3102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11423_ net1226 control.body\[848\] vssd1 vssd1 vccd1 vccd1 _06396_ sky130_fd_sc_hd__xor2_1
XANTENNA__14761__A1 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_3113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15191_ _05559_ net58 vssd1 vssd1 vccd1 vccd1 _01573_ sky130_fd_sc_hd__nor2_4
XFILLER_0_85_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_9 _03446_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14142_ net998 _04052_ _04053_ net1017 _08302_ vssd1 vssd1 vccd1 vccd1 _08303_ sky130_fd_sc_hd__a221o_1
X_11354_ _06319_ _06320_ _06321_ _06326_ vssd1 vssd1 vccd1 vccd1 _06327_ sky130_fd_sc_hd__or4_4
XTAP_TAPCELL_ROW_39_1517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10264__Y _05237_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10705__B net1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10305_ net1096 control.body\[701\] vssd1 vssd1 vccd1 vccd1 _05278_ sky130_fd_sc_hd__nand2_1
XANTENNA__14513__A1 net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15710__B1 _01629_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14513__B2 net1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14073_ _08227_ _08229_ _08231_ _08232_ vssd1 vssd1 vccd1 vccd1 _08234_ sky130_fd_sc_hd__or4_1
X_18950_ clknet_leaf_5_clk img_gen.tracker.next_frame\[388\] net1268 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[388\] sky130_fd_sc_hd__dfrtp_1
X_11285_ net1112 control.body\[1109\] vssd1 vssd1 vccd1 vccd1 _06258_ sky130_fd_sc_hd__nand2_1
X_10236_ ag2.body\[326\] net1090 vssd1 vssd1 vccd1 vccd1 _05209_ sky130_fd_sc_hd__nand2_1
X_17901_ _01691_ _03533_ net48 obsg2.obstacleArray\[0\] vssd1 vssd1 vccd1 vccd1 _03537_
+ sky130_fd_sc_hd__a31o_1
XANTENNA__09782__A net1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13024_ _07707_ net262 _07705_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[274\]
+ sky130_fd_sc_hd__mux2_1
X_18881_ clknet_leaf_11_clk img_gen.tracker.next_frame\[319\] net1281 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[319\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_101_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_89_3031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_3042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1010 net1011 vssd1 vssd1 vccd1 vccd1 net1010 sky130_fd_sc_hd__buf_4
XANTENNA__12920__B net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16266__A1 net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1021 net1024 vssd1 vssd1 vccd1 vccd1 net1021 sky130_fd_sc_hd__buf_4
X_17832_ net971 ag2.apple_cord\[3\] net224 vssd1 vssd1 vccd1 vccd1 _03493_ sky130_fd_sc_hd__mux2_1
Xfanout1032 ag2.randCord\[5\] vssd1 vssd1 vccd1 vccd1 net1032 sky130_fd_sc_hd__clkbuf_8
X_10167_ ag2.body\[578\] net1173 vssd1 vssd1 vccd1 vccd1 _05140_ sky130_fd_sc_hd__xor2_1
Xfanout1043 ag2.body\[1\] vssd1 vssd1 vccd1 vccd1 net1043 sky130_fd_sc_hd__clkbuf_4
XANTENNA__20404__RESET_B net1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1054 net1055 vssd1 vssd1 vccd1 vccd1 net1054 sky130_fd_sc_hd__clkbuf_4
Xfanout1065 net1068 vssd1 vssd1 vccd1 vccd1 net1065 sky130_fd_sc_hd__buf_4
X_17763_ _02966_ _02970_ _02971_ _03441_ _02950_ vssd1 vssd1 vccd1 vccd1 _03442_ sky130_fd_sc_hd__o311a_2
Xfanout1076 net1077 vssd1 vssd1 vccd1 vccd1 net1076 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_83_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10098_ net1084 control.body\[942\] vssd1 vssd1 vccd1 vccd1 _05071_ sky130_fd_sc_hd__xor2_1
XANTENNA__12827__A1 net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1087 net1093 vssd1 vssd1 vccd1 vccd1 net1087 sky130_fd_sc_hd__buf_4
X_14975_ _04614_ net59 vssd1 vssd1 vccd1 vccd1 _01549_ sky130_fd_sc_hd__nor2_2
Xfanout1098 net1106 vssd1 vssd1 vccd1 vccd1 net1098 sky130_fd_sc_hd__buf_2
X_16714_ obsg2.obstacleArray\[127\] net501 net487 obsg2.obstacleArray\[126\] vssd1
+ vssd1 vccd1 vccd1 _02393_ sky130_fd_sc_hd__a22o_1
XFILLER_0_117_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17063__X _02742_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17215__B1 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19502_ clknet_leaf_115_clk _00446_ net1396 vssd1 vssd1 vccd1 vccd1 control.body\[892\]
+ sky130_fd_sc_hd__dfrtp_1
X_13926_ ag2.body\[70\] net134 _08152_ ag2.body\[62\] vssd1 vssd1 vccd1 vccd1 _00151_
+ sky130_fd_sc_hd__a22o_1
X_17694_ ag2.body\[153\] net734 net963 _04047_ _03368_ vssd1 vssd1 vccd1 vccd1 _03373_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_107_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14847__B _08447_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19433_ clknet_leaf_108_clk _00377_ net1434 vssd1 vssd1 vccd1 vccd1 control.body\[967\]
+ sky130_fd_sc_hd__dfrtp_1
X_16645_ obsg2.obstacleArray\[48\] obsg2.obstacleArray\[49\] net444 vssd1 vssd1 vccd1
+ vccd1 _02324_ sky130_fd_sc_hd__mux2_1
X_13857_ ag2.body\[20\] net116 _08134_ ag2.body\[12\] vssd1 vssd1 vccd1 vccd1 _00100_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12648__A net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11552__A net1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12808_ net232 _07605_ _07606_ net1922 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[159\]
+ sky130_fd_sc_hd__a22o_1
X_19364_ clknet_leaf_102_clk _00308_ net1428 vssd1 vssd1 vccd1 vccd1 control.body\[1026\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_128_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16576_ obsg2.obstacleArray\[116\] obsg2.obstacleArray\[117\] net445 vssd1 vssd1
+ vccd1 vccd1 _02255_ sky130_fd_sc_hd__mux2_1
XANTENNA__12055__A2 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13788_ img_gen.updater.commands.count\[13\] _08091_ img_gen.updater.commands.count\[14\]
+ vssd1 vssd1 vccd1 vccd1 _08095_ sky130_fd_sc_hd__a21o_1
XFILLER_0_29_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18315_ _08137_ _03810_ vssd1 vssd1 vccd1 vccd1 _03811_ sky130_fd_sc_hd__and2_1
XANTENNA__11271__B net1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15527_ ag2.body\[530\] net157 _01610_ ag2.body\[522\] vssd1 vssd1 vccd1 vccd1 _00804_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_84_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12739_ net683 _07573_ vssd1 vssd1 vccd1 vccd1 _07574_ sky130_fd_sc_hd__nor2_1
X_19295_ clknet_leaf_98_clk _00239_ net1446 vssd1 vssd1 vccd1 vccd1 control.body\[1101\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__16726__C1 net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_0_clk_A clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18246_ _03687_ net35 vssd1 vssd1 vccd1 vccd1 _03762_ sky130_fd_sc_hd__nor2_1
X_15458_ ag2.body\[597\] net87 _01602_ ag2.body\[589\] vssd1 vssd1 vccd1 vccd1 _00743_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_5_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16741__A2 net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18054__B _03570_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14409_ net1017 net924 vssd1 vssd1 vccd1 vccd1 _08570_ sky130_fd_sc_hd__nand2_1
X_18177_ obsg2.obstacleArray\[85\] _03727_ net532 vssd1 vssd1 vccd1 vccd1 _01336_
+ sky130_fd_sc_hd__o21a_1
XANTENNA__09676__B net1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15389_ net2601 net70 _01595_ net2333 vssd1 vssd1 vccd1 vccd1 _00681_ sky130_fd_sc_hd__a22o_1
XFILLER_0_53_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold504 img_gen.tracker.frame\[429\] vssd1 vssd1 vccd1 vccd1 net2066 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17128_ _02801_ _02802_ _02803_ _02804_ _02806_ vssd1 vssd1 vccd1 vccd1 _02807_ sky130_fd_sc_hd__a221o_1
XFILLER_0_4_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold515 img_gen.tracker.frame\[390\] vssd1 vssd1 vccd1 vccd1 net2077 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold526 img_gen.tracker.frame\[380\] vssd1 vssd1 vccd1 vccd1 net2088 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10615__B _04758_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold537 img_gen.tracker.frame\[198\] vssd1 vssd1 vccd1 vccd1 net2099 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__17238__X _02917_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15694__A _04430_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold548 control.body\[911\] vssd1 vssd1 vccd1 vccd1 net2110 sky130_fd_sc_hd__dlygate4sd3_1
X_17059_ _04004_ net877 net865 _04005_ _02737_ vssd1 vssd1 vccd1 vccd1 _02738_ sky130_fd_sc_hd__a221o_1
Xhold559 img_gen.tracker.frame\[556\] vssd1 vssd1 vccd1 vccd1 net2121 sky130_fd_sc_hd__dlygate4sd3_1
X_09950_ control.body\[738\] net1170 vssd1 vssd1 vccd1 vccd1 _04923_ sky130_fd_sc_hd__nand2b_1
XANTENNA__18070__A net42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_1590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09692__A ag2.body\[65\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20070_ clknet_leaf_73_clk _01014_ net1501 vssd1 vssd1 vccd1 vccd1 ag2.body\[324\]
+ sky130_fd_sc_hd__dfrtp_1
X_09881_ ag2.body\[162\] net1178 vssd1 vssd1 vccd1 vccd1 _04854_ sky130_fd_sc_hd__xor2_1
XFILLER_0_0_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkload18_A clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10631__A net1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__20145__RESET_B net1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_68_2403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout183_A net219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17757__A1 _01742_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17133__B net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout350_A net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1092_A net1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout448_A _02214_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12046__A2 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13243__A1 net238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16980__A2 net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_1459 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11181__B net1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09315_ _04319_ _04324_ _04331_ net272 sound_gen.osc1.count\[4\] vssd1 vssd1 vccd1
+ vccd1 _01439_ sky130_fd_sc_hd__a32o_1
XFILLER_0_118_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16464__S net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18245__A net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16317__X _01996_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout236_X net236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout615_A net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1357_A net1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09246_ score_detect.N\[0\] vssd1 vssd1 vccd1 vccd1 _04271_ sky130_fd_sc_hd__inv_2
XFILLER_0_134_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15588__B net56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16732__A2 net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14743__A1 net993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09177_ ag2.body\[549\] vssd1 vssd1 vccd1 vccd1 _04202_ sky130_fd_sc_hd__inv_2
XFILLER_0_105_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout403_X net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1145_X net1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20406_ clknet_leaf_34_clk _01293_ net1346 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[42\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_32_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout984_A ag2.randCord\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20337_ clknet_leaf_21_clk _01228_ net1363 vssd1 vssd1 vccd1 vccd1 ag2.apple_cord\[5\]
+ sky130_fd_sc_hd__dfrtp_1
Xoutput13 net13 vssd1 vssd1 vccd1 vccd1 gpio_out[12] sky130_fd_sc_hd__buf_2
XFILLER_0_47_1387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput24 net24 vssd1 vssd1 vccd1 vccd1 gpio_out[22] sky130_fd_sc_hd__buf_2
XANTENNA__12580__X _07490_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout96_A net100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11070_ ag2.body\[362\] net776 net785 ag2.body\[360\] vssd1 vssd1 vccd1 vccd1 _06043_
+ sky130_fd_sc_hd__a2bb2o_1
X_20268_ clknet_leaf_37_clk net1582 net1349 vssd1 vssd1 vccd1 vccd1 control.detect2.Q\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__17308__B net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout772_X net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16248__A1 _01912_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10021_ ag2.body\[264\] net1237 vssd1 vssd1 vccd1 vccd1 _04994_ sky130_fd_sc_hd__xor2_1
XANTENNA__17445__B1 net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20199_ clknet_leaf_54_clk _01143_ net1454 vssd1 vssd1 vccd1 vccd1 ag2.body\[197\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_19_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13852__A _05671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14760_ net970 _03989_ ag2.body\[46\] net798 vssd1 vssd1 vccd1 vccd1 _08921_ sky130_fd_sc_hd__o22a_1
XANTENNA__13482__A1 net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout51_X net51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11972_ img_gen.tracker.frame\[526\] net583 net544 img_gen.tracker.frame\[523\] _06943_
+ vssd1 vssd1 vccd1 vccd1 _06944_ sky130_fd_sc_hd__o221a_1
XANTENNA__08946__A net1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13711_ track.highScore\[1\] _04636_ _08050_ vssd1 vssd1 vccd1 vccd1 track.nextHighScore\[1\]
+ sky130_fd_sc_hd__mux2_4
XANTENNA_clkbuf_leaf_2_clk_A clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10923_ ag2.body\[457\] net782 net754 ag2.body\[461\] vssd1 vssd1 vccd1 vccd1 _05896_
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_98_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14691_ _08847_ _08851_ vssd1 vssd1 vccd1 vccd1 _08852_ sky130_fd_sc_hd__nand2_1
XFILLER_0_85_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_19_Right_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13063__S _07723_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16430_ obsg2.obstacleArray\[72\] obsg2.obstacleArray\[73\] net453 vssd1 vssd1 vccd1
+ vccd1 _02109_ sky130_fd_sc_hd__mux2_1
X_13642_ _08002_ net222 _08000_ vssd1 vssd1 vccd1 vccd1 control.divider.next_count\[14\]
+ sky130_fd_sc_hd__and3b_1
XFILLER_0_131_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13234__A1 net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10854_ _04603_ _04758_ net643 _04571_ vssd1 vssd1 vccd1 vccd1 _05827_ sky130_fd_sc_hd__o211ai_4
XANTENNA__12037__A2 net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16882__B net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09989__A1 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16361_ obsg2.obstacleArray\[10\] net409 vssd1 vssd1 vccd1 vccd1 _02040_ sky130_fd_sc_hd__or2_1
XFILLER_0_32_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13573_ _07934_ _07948_ _04282_ vssd1 vssd1 vccd1 vccd1 net24 sky130_fd_sc_hd__mux2_1
XANTENNA__09989__B2 _04943_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12755__X _07581_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10785_ net1195 control.body\[625\] vssd1 vssd1 vccd1 vccd1 _05758_ sky130_fd_sc_hd__nand2_1
XFILLER_0_52_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18100_ obsg2.obstacleArray\[53\] _03682_ net524 vssd1 vssd1 vccd1 vccd1 _01304_
+ sky130_fd_sc_hd__o21a_1
XANTENNA__11796__A1 net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15312_ control.body\[721\] net77 _01588_ net2470 vssd1 vssd1 vccd1 vccd1 _00611_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_32_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19080_ clknet_leaf_29_clk img_gen.tracker.next_frame\[518\] net1334 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[518\] sky130_fd_sc_hd__dfrtp_1
X_12524_ img_gen.tracker.frame\[23\] net649 _07458_ vssd1 vssd1 vccd1 vccd1 _07459_
+ sky130_fd_sc_hd__and3_1
X_16292_ obsg2.obstacleArray\[118\] obsg2.obstacleArray\[119\] net408 vssd1 vssd1
+ vccd1 vccd1 _01971_ sky130_fd_sc_hd__mux2_1
X_18031_ obsg2.obstacleArray\[29\] _03637_ net531 vssd1 vssd1 vccd1 vccd1 _01280_
+ sky130_fd_sc_hd__o21a_1
XANTENNA__17994__A net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15243_ control.body\[790\] net97 _01578_ net2287 vssd1 vssd1 vccd1 vccd1 _00552_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__13299__A net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12455_ _07325_ _07351_ _07413_ _07414_ _07412_ vssd1 vssd1 vccd1 vccd1 _07415_ sky130_fd_sc_hd__a311o_1
XFILLER_0_129_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20607__1539 vssd1 vssd1 vccd1 vccd1 _20607__1539/HI net1539 sky130_fd_sc_hd__conb_1
XFILLER_0_62_591 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11406_ ag2.body\[570\] net1172 vssd1 vssd1 vccd1 vccd1 _06379_ sky130_fd_sc_hd__xor2_1
X_15174_ net2652 net103 _01571_ net2207 vssd1 vssd1 vccd1 vccd1 _00490_ sky130_fd_sc_hd__a22o_1
X_12386_ _07251_ _07254_ _07287_ vssd1 vssd1 vccd1 vccd1 _07351_ sky130_fd_sc_hd__nor3_2
XPHY_EDGE_ROW_28_Right_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16487__A1 net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14125_ net1009 ag2.body\[375\] vssd1 vssd1 vccd1 vccd1 _08286_ sky130_fd_sc_hd__or2_1
XANTENNA__17684__B1 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11337_ _06303_ _06304_ _06309_ vssd1 vssd1 vccd1 vccd1 _06310_ sky130_fd_sc_hd__a21o_1
X_19982_ clknet_leaf_64_clk _00926_ net1474 vssd1 vssd1 vccd1 vccd1 ag2.body\[412\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_103_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18228__A2 _03703_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14056_ net1034 ag2.body\[36\] vssd1 vssd1 vccd1 vccd1 _08217_ sky130_fd_sc_hd__xor2_1
X_18933_ clknet_leaf_140_clk img_gen.tracker.next_frame\[371\] net1294 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[371\] sky130_fd_sc_hd__dfrtp_1
X_11268_ ag2.body\[124\] net1142 vssd1 vssd1 vccd1 vccd1 _06241_ sky130_fd_sc_hd__xor2_1
XFILLER_0_94_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17436__B1 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13007_ net288 _07697_ _07698_ net1883 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[266\]
+ sky130_fd_sc_hd__a22o_1
X_10219_ _04571_ _04758_ net643 vssd1 vssd1 vccd1 vccd1 _05192_ sky130_fd_sc_hd__o21ai_2
X_11199_ net762 control.body\[876\] control.body\[877\] net754 _06171_ vssd1 vssd1
+ vccd1 vccd1 _06172_ sky130_fd_sc_hd__a221o_1
XANTENNA__13465__C net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18864_ clknet_leaf_26_clk img_gen.tracker.next_frame\[302\] net1344 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[302\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17815_ net924 _08124_ vssd1 vssd1 vccd1 vccd1 _03482_ sky130_fd_sc_hd__nor2_1
X_18795_ clknet_leaf_22_clk img_gen.tracker.next_frame\[233\] net1358 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[233\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_94_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15462__A2 net90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17746_ _02516_ _02519_ _03070_ _03424_ vssd1 vssd1 vccd1 vccd1 _03425_ sky130_fd_sc_hd__o211a_1
X_14958_ net2260 net172 _01547_ control.body\[1024\] vssd1 vssd1 vccd1 vccd1 _00298_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__17739__A1 _02844_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13473__A1 net250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_37_Right_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18049__B _03562_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13909_ ag2.body\[55\] net119 _08150_ ag2.body\[47\] vssd1 vssd1 vccd1 vccd1 _00136_
+ sky130_fd_sc_hd__a22o_1
X_17677_ ag2.body\[472\] net737 net947 _04170_ vssd1 vssd1 vccd1 vccd1 _03356_ sky130_fd_sc_hd__a22o_1
X_14889_ control.body\[1099\] net180 _01539_ net2186 vssd1 vssd1 vccd1 vccd1 _00237_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_58_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16411__A1 net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11282__A net1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16628_ _02304_ _02305_ _02306_ net394 net361 vssd1 vssd1 vccd1 vccd1 _02307_ sky130_fd_sc_hd__a221o_1
X_19416_ clknet_leaf_103_clk _00360_ net1427 vssd1 vssd1 vccd1 vccd1 control.body\[982\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_134_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19839__RESET_B net1414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16559_ obsg2.obstacleArray\[104\] obsg2.obstacleArray\[105\] net442 vssd1 vssd1
+ vccd1 vccd1 _02238_ sky130_fd_sc_hd__mux2_1
X_19347_ clknet_leaf_101_clk _00291_ net1439 vssd1 vssd1 vccd1 vccd1 control.body\[1041\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14593__A net1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09100_ ag2.body\[351\] vssd1 vssd1 vccd1 vccd1 _04125_ sky130_fd_sc_hd__inv_2
XANTENNA__18832__CLK clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19278_ clknet_leaf_97_clk _00222_ net1450 vssd1 vssd1 vccd1 vccd1 control.body\[1116\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__16714__A2 net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11882__S1 net1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09031_ ag2.body\[178\] vssd1 vssd1 vccd1 vccd1 _04056_ sky130_fd_sc_hd__inv_2
X_18229_ net519 _03753_ vssd1 vssd1 vccd1 vccd1 _01362_ sky130_fd_sc_hd__nor2_1
XFILLER_0_26_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_46_Right_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_1641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18467__A2 net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold301 img_gen.tracker.frame\[336\] vssd1 vssd1 vccd1 vccd1 net1863 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09601__B1 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20397__RESET_B net1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold312 img_gen.tracker.frame\[372\] vssd1 vssd1 vccd1 vccd1 net1874 sky130_fd_sc_hd__dlygate4sd3_1
Xhold323 img_gen.tracker.frame\[47\] vssd1 vssd1 vccd1 vccd1 net1885 sky130_fd_sc_hd__dlygate4sd3_1
Xhold334 img_gen.tracker.frame\[471\] vssd1 vssd1 vccd1 vccd1 net1896 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18982__CLK clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12841__A _07431_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold345 img_gen.tracker.frame\[143\] vssd1 vssd1 vccd1 vccd1 net1907 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__20326__RESET_B net1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold356 img_gen.tracker.frame\[354\] vssd1 vssd1 vccd1 vccd1 net1918 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold367 img_gen.tracker.frame\[77\] vssd1 vssd1 vccd1 vccd1 net1929 sky130_fd_sc_hd__dlygate4sd3_1
X_20122_ clknet_leaf_81_clk _01066_ net1485 vssd1 vssd1 vccd1 vccd1 ag2.body\[264\]
+ sky130_fd_sc_hd__dfrtp_4
Xhold378 img_gen.tracker.frame\[388\] vssd1 vssd1 vccd1 vccd1 net1940 sky130_fd_sc_hd__dlygate4sd3_1
X_09933_ ag2.body\[30\] net1078 vssd1 vssd1 vccd1 vccd1 _04906_ sky130_fd_sc_hd__xor2_1
Xhold389 toggle1.bcd_tens\[3\] vssd1 vssd1 vccd1 vccd1 net1951 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout803 net804 vssd1 vssd1 vccd1 vccd1 net803 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_106_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12560__B _06638_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout814 net816 vssd1 vssd1 vccd1 vccd1 net814 sky130_fd_sc_hd__clkbuf_4
Xfanout825 net827 vssd1 vssd1 vccd1 vccd1 net825 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_0_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout398_A net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17427__B1 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20053_ clknet_leaf_72_clk _00997_ net1501 vssd1 vssd1 vccd1 vccd1 ag2.body\[339\]
+ sky130_fd_sc_hd__dfrtp_4
Xfanout836 _03965_ vssd1 vssd1 vccd1 vccd1 net836 sky130_fd_sc_hd__buf_2
XFILLER_0_110_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout847 _03963_ vssd1 vssd1 vccd1 vccd1 net847 sky130_fd_sc_hd__clkbuf_4
X_09864_ ag2.body\[159\] net1065 vssd1 vssd1 vccd1 vccd1 _04837_ sky130_fd_sc_hd__nand2_1
XANTENNA__10361__A _04983_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout858 net859 vssd1 vssd1 vccd1 vccd1 net858 sky130_fd_sc_hd__buf_4
XANTENNA_fanout1105_A net1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout869 obsg2.randCord\[1\] vssd1 vssd1 vccd1 vccd1 net869 sky130_fd_sc_hd__clkbuf_8
Xhold1001 control.body\[676\] vssd1 vssd1 vccd1 vccd1 net2563 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__16967__B net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1012 control.body\[673\] vssd1 vssd1 vccd1 vccd1 net2574 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1023 control.body\[724\] vssd1 vssd1 vccd1 vccd1 net2585 sky130_fd_sc_hd__dlygate4sd3_1
X_09795_ net1161 control.body\[963\] vssd1 vssd1 vccd1 vccd1 _04768_ sky130_fd_sc_hd__xor2_1
Xhold1034 control.body\[661\] vssd1 vssd1 vccd1 vccd1 net2596 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14768__A net1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1045 control.body\[719\] vssd1 vssd1 vccd1 vccd1 net2607 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_55_Right_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout565_A net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13672__A net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1056 control.body\[1031\] vssd1 vssd1 vccd1 vccd1 net2618 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1067 control.body\[773\] vssd1 vssd1 vccd1 vccd1 net2629 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1078 control.body\[881\] vssd1 vssd1 vccd1 vccd1 net2640 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13464__A1 net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1089 control.body\[976\] vssd1 vssd1 vccd1 vccd1 net2651 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_36_1011 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19488__CLK clknet_leaf_113_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout732_A net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1095_X net1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11192__A net1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12019__A2 net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17798__B net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_1256 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout618_X net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19509__RESET_B net1403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10570_ net641 _04519_ vssd1 vssd1 vccd1 vccd1 _05543_ sky130_fd_sc_hd__nor2_2
XFILLER_0_88_1443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_64_Right_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_295 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09229_ control.body\[1084\] vssd1 vssd1 vccd1 vccd1 _04254_ sky130_fd_sc_hd__inv_2
XFILLER_0_106_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15913__B1 _01652_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19162__RESET_B net1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12240_ _07187_ _07208_ _07209_ _07204_ _04274_ vssd1 vssd1 vccd1 vccd1 _07210_ sky130_fd_sc_hd__a32o_1
XFILLER_0_115_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout987_X net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16469__B2 net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12171_ net560 _07139_ _07140_ _07142_ vssd1 vssd1 vccd1 vccd1 _07143_ sky130_fd_sc_hd__a22o_1
XANTENNA__12751__A net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17130__A2 net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11122_ net1202 control.body\[865\] vssd1 vssd1 vccd1 vccd1 _06095_ sky130_fd_sc_hd__or2_1
XFILLER_0_120_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold890 control.body\[750\] vssd1 vssd1 vccd1 vccd1 net2452 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__17418__B1 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15930_ ag2.body\[168\] net126 _01655_ ag2.body\[160\] vssd1 vssd1 vccd1 vccd1 _01162_
+ sky130_fd_sc_hd__a22o_1
X_11053_ ag2.body\[387\] net1154 vssd1 vssd1 vccd1 vccd1 _06026_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_73_Right_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10004_ net1074 control.body\[734\] vssd1 vssd1 vccd1 vccd1 _04977_ sky130_fd_sc_hd__nand2_1
XANTENNA__18091__B1 net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15861_ ag2.body\[236\] net175 _01646_ ag2.body\[228\] vssd1 vssd1 vccd1 vccd1 _01102_
+ sky130_fd_sc_hd__a22o_1
X_17600_ ag2.body\[419\] net852 vssd1 vssd1 vccd1 vccd1 _03279_ sky130_fd_sc_hd__xor2_1
XFILLER_0_56_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14812_ net833 ag2.body\[377\] ag2.body\[379\] net818 vssd1 vssd1 vccd1 vccd1 _01483_
+ sky130_fd_sc_hd__a2bb2o_1
X_18580_ clknet_leaf_14_clk img_gen.tracker.next_frame\[18\] net1279 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[18\] sky130_fd_sc_hd__dfrtp_1
X_15792_ ag2.body\[302\] net208 _01639_ ag2.body\[294\] vssd1 vssd1 vccd1 vccd1 _01040_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_54_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17531_ ag2.body\[273\] net873 vssd1 vssd1 vccd1 vccd1 _03210_ sky130_fd_sc_hd__or2_1
XANTENNA__17989__A net45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14743_ net993 _04114_ _08897_ _08899_ _08903_ vssd1 vssd1 vccd1 vccd1 _08904_ sky130_fd_sc_hd__a2111o_4
XFILLER_0_59_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11955_ net563 _06904_ _06906_ net467 vssd1 vssd1 vccd1 vccd1 _06927_ sky130_fd_sc_hd__a31o_1
XFILLER_0_59_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12198__A _07169_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_120_3971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10906_ net1145 control.body\[675\] vssd1 vssd1 vccd1 vccd1 _05879_ sky130_fd_sc_hd__xor2_1
X_17462_ ag2.body\[531\] net853 vssd1 vssd1 vccd1 vccd1 _03141_ sky130_fd_sc_hd__xor2_1
XFILLER_0_135_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14674_ net1000 ag2.body\[384\] vssd1 vssd1 vccd1 vccd1 _08835_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_120_3982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13207__A1 net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11886_ img_gen.tracker.frame\[28\] net606 net590 img_gen.tracker.frame\[34\] _06857_
+ vssd1 vssd1 vccd1 vccd1 _06858_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_120_3993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16413_ obsg2.obstacleArray\[103\] _02059_ net397 _02091_ vssd1 vssd1 vccd1 vccd1
+ _02092_ sky130_fd_sc_hd__o211a_1
X_19201_ clknet_leaf_86_clk _00145_ net1461 vssd1 vssd1 vccd1 vccd1 ag2.body\[64\]
+ sky130_fd_sc_hd__dfrtp_4
X_13625_ _07990_ _07991_ net220 vssd1 vssd1 vccd1 vccd1 control.divider.next_count\[8\]
+ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_101_3392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_1218 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10837_ _05806_ _05807_ _05808_ _05809_ vssd1 vssd1 vccd1 vccd1 _05810_ sky130_fd_sc_hd__a22o_1
X_17393_ ag2.body\[507\] net853 vssd1 vssd1 vccd1 vccd1 _03072_ sky130_fd_sc_hd__xor2_1
XANTENNA__17501__B net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_82_Right_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_17_Left_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11769__A1 net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19132_ clknet_leaf_141_clk img_gen.tracker.next_frame\[570\] net1294 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[570\] sky130_fd_sc_hd__dfrtp_1
X_16344_ _02021_ _02022_ net418 vssd1 vssd1 vccd1 vccd1 _02023_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16157__B1 _01729_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13556_ ssdec1.in\[1\] ssdec1.in\[0\] vssd1 vssd1 vccd1 vccd1 _07938_ sky130_fd_sc_hd__nand2_1
XFILLER_0_125_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10768_ ag2.body\[216\] net1237 vssd1 vssd1 vccd1 vccd1 _05741_ sky130_fd_sc_hd__xor2_1
XFILLER_0_89_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12507_ net315 _07449_ vssd1 vssd1 vccd1 vccd1 _07450_ sky130_fd_sc_hd__or2_1
X_19063_ clknet_leaf_8_clk img_gen.tracker.next_frame\[501\] net1270 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[501\] sky130_fd_sc_hd__dfrtp_1
X_16275_ net419 _01953_ _01952_ net370 vssd1 vssd1 vccd1 vccd1 _01954_ sky130_fd_sc_hd__a211o_1
XANTENNA__15021__B net66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_max_cap363_A _02076_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13487_ net2095 net644 _07906_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[538\]
+ sky130_fd_sc_hd__and3_1
X_10699_ ag2.body\[23\] net1054 vssd1 vssd1 vccd1 vccd1 _05672_ sky130_fd_sc_hd__nand2_1
X_18014_ net351 _03624_ vssd1 vssd1 vccd1 vccd1 _03625_ sky130_fd_sc_hd__nand2_1
X_15226_ net2208 net93 _01576_ control.body\[799\] vssd1 vssd1 vccd1 vccd1 _00537_
+ sky130_fd_sc_hd__a22o_1
X_12438_ net748 _06629_ vssd1 vssd1 vccd1 vccd1 _07399_ sky130_fd_sc_hd__and2_1
XFILLER_0_2_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_114_3786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10165__B net1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_114_3797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15157_ control.body\[857\] net105 _01569_ net2545 vssd1 vssd1 vccd1 vccd1 _00475_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_65_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12369_ _06634_ _07301_ vssd1 vssd1 vccd1 vccd1 _07335_ sky130_fd_sc_hd__nor2_2
XANTENNA__12661__A net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14108_ net997 ag2.body\[568\] vssd1 vssd1 vccd1 vccd1 _08269_ sky130_fd_sc_hd__nand2_1
X_19965_ clknet_leaf_62_clk _00909_ net1469 vssd1 vssd1 vccd1 vccd1 ag2.body\[427\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_120_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15088_ net2242 net148 _01562_ net2463 vssd1 vssd1 vccd1 vccd1 _00413_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_91_Right_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_26_Left_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14039_ _08198_ _08199_ vssd1 vssd1 vccd1 vccd1 _08200_ sky130_fd_sc_hd__nand2_1
X_18916_ clknet_leaf_142_clk img_gen.tracker.next_frame\[354\] net1253 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[354\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__20338__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19896_ clknet_leaf_85_clk _00840_ net1462 vssd1 vssd1 vccd1 vccd1 ag2.body\[502\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__17890__C _03529_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18847_ clknet_leaf_4_clk img_gen.tracker.next_frame\[285\] net1277 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[285\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__16279__S net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09580_ _04471_ _04550_ net892 vssd1 vssd1 vccd1 vccd1 _04553_ sky130_fd_sc_hd__a21oi_4
X_18778_ clknet_leaf_17_clk img_gen.tracker.next_frame\[216\] net1318 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[216\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17899__A net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17729_ obsg2.obstacleArray\[136\] net493 net484 obsg2.obstacleArray\[137\] _03407_
+ vssd1 vssd1 vccd1 vccd1 _03408_ sky130_fd_sc_hd__a221o_1
XFILLER_0_78_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20098__Q ag2.body\[288\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_35_Left_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19780__CLK clknet_leaf_127_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkload85_A clknet_leaf_102_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19673__RESET_B net1386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17411__B net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12836__A net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout146_A net183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_560 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12555__B _07476_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09210__A net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1055_A net1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09014_ ag2.body\[142\] vssd1 vssd1 vccd1 vccd1 _04039_ sky130_fd_sc_hd__inv_2
XANTENNA__16794__S1 net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18242__B net35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold120 img_gen.tracker.frame\[116\] vssd1 vssd1 vccd1 vccd1 net1682 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09864__B net1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold131 img_gen.tracker.frame\[79\] vssd1 vssd1 vccd1 vccd1 net1693 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_48_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold142 img_gen.tracker.frame\[306\] vssd1 vssd1 vccd1 vccd1 net1704 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1222_A net1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold153 img_gen.tracker.frame\[353\] vssd1 vssd1 vccd1 vccd1 net1715 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_44_Left_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10735__A2 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold164 obsg2.obsNeeded\[3\] vssd1 vssd1 vccd1 vccd1 net1726 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1060 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold175 img_gen.tracker.frame\[279\] vssd1 vssd1 vccd1 vccd1 net1737 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout682_A net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold186 img_gen.tracker.frame\[296\] vssd1 vssd1 vccd1 vccd1 net1748 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10803__B net1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18728__CLK clknet_leaf_142_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold197 img_gen.tracker.frame\[168\] vssd1 vssd1 vccd1 vccd1 net1759 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout600 net602 vssd1 vssd1 vccd1 vccd1 net600 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_106_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20105_ clknet_leaf_79_clk _01049_ net1489 vssd1 vssd1 vccd1 vccd1 ag2.body\[295\]
+ sky130_fd_sc_hd__dfrtp_4
Xfanout611 _06475_ vssd1 vssd1 vccd1 vccd1 net611 sky130_fd_sc_hd__clkbuf_4
X_09916_ _04882_ _04883_ _04884_ _04888_ vssd1 vssd1 vccd1 vccd1 _04889_ sky130_fd_sc_hd__or4_1
Xfanout622 net625 vssd1 vssd1 vccd1 vccd1 net622 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout1010_X net1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10091__A net1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout644 net645 vssd1 vssd1 vccd1 vccd1 net644 sky130_fd_sc_hd__buf_2
XANTENNA__13685__A1 net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_6_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_15_clk_X clknet_leaf_15_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1108_X net1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout655 net656 vssd1 vssd1 vccd1 vccd1 net655 sky130_fd_sc_hd__clkbuf_2
X_20036_ clknet_leaf_67_clk _00980_ net1495 vssd1 vssd1 vccd1 vccd1 ag2.body\[354\]
+ sky130_fd_sc_hd__dfrtp_4
Xfanout666 net674 vssd1 vssd1 vccd1 vccd1 net666 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout677 net681 vssd1 vssd1 vccd1 vccd1 net677 sky130_fd_sc_hd__buf_2
X_09847_ net1133 control.body\[972\] vssd1 vssd1 vccd1 vccd1 _04820_ sky130_fd_sc_hd__nand2_1
XANTENNA__11696__B1 _06661_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16189__S net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout688 net695 vssd1 vssd1 vccd1 vccd1 net688 sky130_fd_sc_hd__buf_4
XANTENNA_fanout947_A net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout699 net700 vssd1 vssd1 vccd1 vccd1 net699 sky130_fd_sc_hd__clkbuf_4
XANTENNA__14498__A net1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16084__C1 net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout568_X net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_4093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13437__A1 net235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09778_ ag2.body\[235\] net770 net1111 _04073_ _04742_ vssd1 vssd1 vccd1 vccd1 _04751_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_77_1188 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout59_A net62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20606__1538 vssd1 vssd1 vccd1 vccd1 _20606__1538/HI net1538 sky130_fd_sc_hd__conb_1
XFILLER_0_115_1318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_1_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17179__A2 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout735_X net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1477_X net1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_53_Left_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_1415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11740_ img_gen.tracker.frame\[23\] net590 vssd1 vssd1 vccd1 vccd1 _06712_ sky130_fd_sc_hd__or2_1
XFILLER_0_132_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10671__A1 _04418_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11671_ _06628_ _06642_ vssd1 vssd1 vccd1 vccd1 _06643_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout902_X net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10671__B2 _05643_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16218__A net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_137_4487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11650__A _06497_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13410_ _07558_ net303 vssd1 vssd1 vccd1 vccd1 _07876_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_137_4498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10622_ ag2.body\[51\] net1150 vssd1 vssd1 vccd1 vccd1 _05595_ sky130_fd_sc_hd__xor2_1
X_14390_ net830 ag2.body\[298\] ag2.body\[303\] net795 _08550_ vssd1 vssd1 vccd1 vccd1
+ _08551_ sky130_fd_sc_hd__o221a_1
XFILLER_0_119_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11620__B1 net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13341_ net274 _07848_ _07849_ net1622 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[449\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__10423__B2 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10553_ _05515_ _05516_ _05520_ _05521_ _05525_ vssd1 vssd1 vccd1 vccd1 _05526_ sky130_fd_sc_hd__a221o_1
XANTENNA__10266__A _05237_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16652__S net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_703 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17975__C net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_580 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16060_ _01726_ _01738_ vssd1 vssd1 vccd1 vccd1 _01739_ sky130_fd_sc_hd__nor2_1
XANTENNA__15776__B net60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19503__CLK clknet_leaf_113_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13272_ net282 _07821_ _07822_ net1618 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[407\]
+ sky130_fd_sc_hd__a22o_1
X_10484_ ag2.body\[587\] net767 net743 ag2.body\[591\] _05456_ vssd1 vssd1 vccd1 vccd1
+ _05457_ sky130_fd_sc_hd__o221a_1
XFILLER_0_20_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15011_ _05573_ net58 vssd1 vssd1 vccd1 vccd1 _01553_ sky130_fd_sc_hd__nor2_4
X_12223_ img_gen.updater.commands.count\[10\] img_gen.updater.commands.count\[11\]
+ img_gen.updater.commands.count\[12\] vssd1 vssd1 vccd1 vccd1 _07193_ sky130_fd_sc_hd__a21o_1
XANTENNA__09774__B net1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17103__A2 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12912__C _07638_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12154_ img_gen.tracker.frame\[474\] net540 vssd1 vssd1 vccd1 vccd1 _07126_ sky130_fd_sc_hd__or2_1
XFILLER_0_124_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11105_ net1160 control.body\[1099\] vssd1 vssd1 vccd1 vccd1 _06078_ sky130_fd_sc_hd__and2_1
XFILLER_0_100_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19750_ clknet_leaf_129_clk _00694_ net1325 vssd1 vssd1 vccd1 vccd1 control.body\[644\]
+ sky130_fd_sc_hd__dfrtp_1
X_16962_ _02639_ _02640_ _02638_ vssd1 vssd1 vccd1 vccd1 _02641_ sky130_fd_sc_hd__a21o_1
X_12085_ img_gen.tracker.frame\[324\] net629 net556 img_gen.tracker.frame\[330\] _07056_
+ vssd1 vssd1 vccd1 vccd1 _07057_ sky130_fd_sc_hd__a221o_1
XANTENNA__09790__A net1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18701_ clknet_leaf_9_clk img_gen.tracker.next_frame\[139\] net1274 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[139\] sky130_fd_sc_hd__dfrtp_1
X_15913_ ag2.body\[186\] net130 _01652_ ag2.body\[178\] vssd1 vssd1 vccd1 vccd1 _01148_
+ sky130_fd_sc_hd__a22o_1
X_11036_ control.body\[1043\] net1159 vssd1 vssd1 vccd1 vccd1 _06009_ sky130_fd_sc_hd__nand2b_1
XANTENNA__16099__S net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16893_ _02569_ _02570_ _02571_ _02568_ vssd1 vssd1 vccd1 vccd1 _02572_ sky130_fd_sc_hd__a211o_1
X_19681_ clknet_leaf_117_clk _00625_ net1385 vssd1 vssd1 vccd1 vccd1 control.body\[719\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18632_ clknet_leaf_145_clk img_gen.tracker.next_frame\[70\] net1242 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[70\] sky130_fd_sc_hd__dfrtp_1
X_15844_ ag2.body\[253\] net176 _01644_ ag2.body\[245\] vssd1 vssd1 vccd1 vccd1 _01087_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11502__A_N net1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_3590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15775_ ag2.body\[319\] net209 _01637_ ag2.body\[311\] vssd1 vssd1 vccd1 vccd1 _01025_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_91_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18563_ clknet_leaf_15_clk img_gen.tracker.next_frame\[1\] net1312 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[1\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_103_3454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12987_ net233 _07688_ _07689_ net1719 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[255\]
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_103_3465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_3476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14726_ net1023 ag2.body\[118\] vssd1 vssd1 vccd1 vccd1 _08887_ sky130_fd_sc_hd__xor2_1
XFILLER_0_87_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17514_ ag2.body\[585\] net730 net848 _04215_ _03192_ vssd1 vssd1 vccd1 vccd1 _03193_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_59_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18494_ net1516 net1510 vssd1 vssd1 vccd1 vccd1 _00025_ sky130_fd_sc_hd__or2_1
X_11938_ img_gen.tracker.frame\[145\] net621 net603 img_gen.tracker.frame\[148\] vssd1
+ vssd1 vccd1 vccd1 _06910_ sky130_fd_sc_hd__o22a_1
XFILLER_0_59_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17445_ ag2.body\[380\] net709 net949 _04137_ _03123_ vssd1 vssd1 vccd1 vccd1 _03124_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_68_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14657_ net1040 _04042_ ag2.body\[150\] net802 _08811_ vssd1 vssd1 vccd1 vccd1 _08818_
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_89_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18119__A1 net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12656__A net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11869_ img_gen.tracker.frame\[286\] net581 net574 vssd1 vssd1 vccd1 vccd1 _06841_
+ sky130_fd_sc_hd__o21a_1
XANTENNA__17590__A2 net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13608_ control.divider.count\[1\] net2159 _07981_ vssd1 vssd1 vccd1 vccd1 control.divider.next_count\[1\]
+ sky130_fd_sc_hd__a21oi_1
X_17376_ _03018_ _03052_ _03051_ vssd1 vssd1 vccd1 vccd1 _03055_ sky130_fd_sc_hd__mux2_1
X_14588_ net994 _04012_ ag2.body\[83\] net822 _08748_ vssd1 vssd1 vccd1 vccd1 _08749_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_27_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_116_3848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16327_ obsg2.obstacleArray\[73\] net413 _02005_ net418 vssd1 vssd1 vccd1 vccd1 _02006_
+ sky130_fd_sc_hd__o211a_1
X_19115_ clknet_leaf_141_clk img_gen.tracker.next_frame\[553\] net1295 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[553\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__10414__A1 _05364_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12806__D _07508_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13539_ _06821_ net309 _07630_ vssd1 vssd1 vccd1 vccd1 _07927_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_116_3859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19183__CLK clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19046_ clknet_leaf_8_clk img_gen.tracker.next_frame\[484\] net1273 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[484\] sky130_fd_sc_hd__dfrtp_1
X_16258_ net417 _01934_ _01936_ net369 vssd1 vssd1 vccd1 vccd1 _01937_ sky130_fd_sc_hd__a211o_1
XFILLER_0_109_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15209_ _06331_ net53 vssd1 vssd1 vccd1 vccd1 _01575_ sky130_fd_sc_hd__nor2_2
XFILLER_0_23_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09684__B net1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16189_ _01866_ _01867_ net373 vssd1 vssd1 vccd1 vccd1 _01868_ sky130_fd_sc_hd__mux2_1
XANTENNA__12391__A net1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10904__A net1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10717__A2 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_1568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10623__B net1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15656__A2 net139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09971__Y _04944_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_2476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19948_ clknet_leaf_45_clk _00892_ net1382 vssd1 vssd1 vccd1 vccd1 ag2.body\[442\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_71_2487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_2498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09701_ _04670_ _04671_ _04672_ _04673_ vssd1 vssd1 vccd1 vccd1 _04674_ sky130_fd_sc_hd__a22o_1
XFILLER_0_4_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17406__B net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19879_ clknet_leaf_91_clk _00823_ net1415 vssd1 vssd1 vccd1 vccd1 ag2.body\[517\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__11182__A_N net1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11294__X _06267_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09632_ net897 _04602_ _04492_ vssd1 vssd1 vccd1 vccd1 _04605_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_74_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13419__A1 net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14111__A net1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_2995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09205__A net1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09563_ _04495_ _04496_ _04503_ _04535_ _04484_ vssd1 vssd1 vccd1 vccd1 _04536_ sky130_fd_sc_hd__o311a_1
XANTENNA_fanout263_A net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11525__S0 net1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09494_ ag2.body\[374\] net1081 vssd1 vssd1 vccd1 vccd1 _04467_ sky130_fd_sc_hd__xor2_1
XANTENNA__16369__B1 _01919_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16908__A2 net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17141__B net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout430_A _01734_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_42_clk_A clknet_4_7__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16038__A net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1172_A net1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout528_A net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17581__A2 net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_1226 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11828__S1 net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_132_4340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_4351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20585_ clknet_leaf_107_clk _01442_ _00049_ vssd1 vssd1 vccd1 vccd1 sound_gen.osc1.count\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10086__A net1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout316_X net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14781__A net1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_132_4362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_1435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1058_X net1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1437_A net1442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09875__A ag2.body\[163\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_57_clk_A clknet_4_12__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18550__CLK clknet_leaf_132_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout897_A net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15895__A2 net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_100_clk_A clknet_4_11__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1225_X net1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12732__C _07460_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09574__A2 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_1491 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout685_X net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1406 net1409 vssd1 vssd1 vccd1 vccd1 net1406 sky130_fd_sc_hd__clkbuf_4
Xfanout1417 net1419 vssd1 vssd1 vccd1 vccd1 net1417 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_54_1962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout430 _01734_ vssd1 vssd1 vccd1 vccd1 net430 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_79_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1428 net1430 vssd1 vssd1 vccd1 vccd1 net1428 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_54_1973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_1490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout441 net443 vssd1 vssd1 vccd1 vccd1 net441 sky130_fd_sc_hd__buf_2
Xfanout1439 net1442 vssd1 vssd1 vccd1 vccd1 net1439 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_54_1984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout452 net453 vssd1 vssd1 vccd1 vccd1 net452 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_126_4177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout463 _01709_ vssd1 vssd1 vccd1 vccd1 net463 sky130_fd_sc_hd__buf_8
XANTENNA_clkbuf_leaf_115_clk_A clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout852_X net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17316__B net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_1394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout474 _06647_ vssd1 vssd1 vccd1 vccd1 net474 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_50_1848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout485 _02373_ vssd1 vssd1 vccd1 vccd1 net485 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_50_1859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20019_ clknet_leaf_58_clk _00963_ net1471 vssd1 vssd1 vccd1 vccd1 ag2.body\[369\]
+ sky130_fd_sc_hd__dfrtp_4
Xfanout496 _01712_ vssd1 vssd1 vccd1 vccd1 net496 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_6_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12910_ _07315_ net227 vssd1 vssd1 vccd1 vccd1 _07653_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_31_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14021__A net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13890_ ag2.body\[38\] net115 _08148_ ag2.body\[30\] vssd1 vssd1 vccd1 vccd1 _00119_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_31_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10341__B1 net1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_61_Left_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12841_ _07431_ _07621_ vssd1 vssd1 vccd1 vccd1 _07622_ sky130_fd_sc_hd__nor2_1
XANTENNA__19056__CLK clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16647__S net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14083__A1 net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_520 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14083__B2 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1130 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15560_ _04687_ net61 vssd1 vssd1 vccd1 vccd1 _01614_ sky130_fd_sc_hd__nor2_2
XFILLER_0_55_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12772_ net281 _07588_ _07589_ net1941 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[140\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_51_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14511_ _08664_ _08665_ _08667_ _08668_ vssd1 vssd1 vccd1 vccd1 _08672_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_48_1777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11723_ img_gen.tracker.frame\[233\] net608 net592 img_gen.tracker.frame\[239\] _06694_
+ vssd1 vssd1 vccd1 vccd1 _06695_ sky130_fd_sc_hd__o221a_1
X_15491_ ag2.body\[562\] net109 _01606_ ag2.body\[554\] vssd1 vssd1 vccd1 vccd1 _00772_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11841__B1 net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09769__B net1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_48_1799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17230_ _04156_ net883 net851 _04157_ vssd1 vssd1 vccd1 vccd1 _02909_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_29_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14442_ net1010 ag2.body\[231\] vssd1 vssd1 vccd1 vccd1 _08603_ sky130_fd_sc_hd__xor2_1
XFILLER_0_65_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11654_ net758 net748 vssd1 vssd1 vccd1 vccd1 _06627_ sky130_fd_sc_hd__nor2_1
XANTENNA__10708__B net1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16890__B net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout70 net91 vssd1 vssd1 vccd1 vccd1 net70 sky130_fd_sc_hd__buf_1
XFILLER_0_126_349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout81 net83 vssd1 vssd1 vccd1 vccd1 net81 sky130_fd_sc_hd__buf_2
XFILLER_0_107_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout92 net100 vssd1 vssd1 vccd1 vccd1 net92 sky130_fd_sc_hd__buf_2
X_10605_ net1060 control.body\[991\] vssd1 vssd1 vccd1 vccd1 _05578_ sky130_fd_sc_hd__nand2_1
X_17161_ ag2.body\[599\] net928 vssd1 vssd1 vccd1 vccd1 _02840_ sky130_fd_sc_hd__or2_1
X_14373_ net981 ag2.body\[418\] vssd1 vssd1 vccd1 vccd1 _08534_ sky130_fd_sc_hd__xor2_1
XFILLER_0_68_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11585_ net1192 net1144 vssd1 vssd1 vccd1 vccd1 _06558_ sky130_fd_sc_hd__or2_1
XFILLER_0_101_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16112_ obsg2.obstacleArray\[68\] obsg2.obstacleArray\[69\] net426 vssd1 vssd1 vccd1
+ vccd1 _01791_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13324_ net229 _07842_ _07843_ net2009 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[438\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_52_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_94_3177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17092_ ag2.body\[301\] net955 vssd1 vssd1 vccd1 vccd1 _02771_ sky130_fd_sc_hd__xor2_1
XFILLER_0_80_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10536_ _05501_ _05506_ _05507_ _05508_ vssd1 vssd1 vccd1 vccd1 _05509_ sky130_fd_sc_hd__or4_2
XFILLER_0_68_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_3701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_3712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_3188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_3723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_3199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12923__B net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16043_ net350 _01720_ net355 vssd1 vssd1 vccd1 vccd1 _01722_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_108_Right_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13255_ net234 _07815_ _07816_ net1601 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[396\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_126_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10467_ net1059 control.body\[1015\] vssd1 vssd1 vccd1 vccd1 _05440_ sky130_fd_sc_hd__nand2_1
X_12206_ _07177_ _04259_ img_gen.control.current\[0\] vssd1 vssd1 vccd1 vccd1 _07178_
+ sky130_fd_sc_hd__and3b_1
XFILLER_0_62_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13100__A net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_1288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13186_ net675 _07783_ vssd1 vssd1 vccd1 vccd1 _07784_ sky130_fd_sc_hd__nor2_1
X_10398_ net1230 control.body\[1056\] vssd1 vssd1 vccd1 vccd1 _05371_ sky130_fd_sc_hd__xor2_1
XANTENNA__16296__C1 net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11372__A2 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19802_ clknet_leaf_125_clk _00746_ net1410 vssd1 vssd1 vccd1 vccd1 ag2.body\[584\]
+ sky130_fd_sc_hd__dfrtp_4
X_12137_ img_gen.tracker.frame\[492\] net616 vssd1 vssd1 vccd1 vccd1 _07109_ sky130_fd_sc_hd__or2_1
XFILLER_0_40_1530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17994_ net381 _01737_ _03561_ vssd1 vssd1 vccd1 vccd1 _03610_ sky130_fd_sc_hd__or3b_1
XFILLER_0_19_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_109_3641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19733_ clknet_leaf_129_clk _00677_ net1327 vssd1 vssd1 vccd1 vccd1 control.body\[659\]
+ sky130_fd_sc_hd__dfrtp_1
X_16945_ ag2.body\[389\] net949 vssd1 vssd1 vccd1 vccd1 _02624_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_109_3652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12068_ net1225 net1199 img_gen.tracker.frame\[117\] vssd1 vssd1 vccd1 vccd1 _07040_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_105_3516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_3527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11019_ ag2.body\[593\] net1196 vssd1 vssd1 vccd1 vccd1 _05992_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_105_3538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19664_ clknet_leaf_134_clk _00608_ net1309 vssd1 vssd1 vccd1 vccd1 control.body\[734\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_56_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16876_ _02546_ _02547_ _02548_ _02554_ vssd1 vssd1 vccd1 vccd1 _02555_ sky130_fd_sc_hd__a211o_1
XANTENNA__18052__A3 net39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1014 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09025__A ag2.body\[161\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11274__B net1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18615_ clknet_leaf_146_clk img_gen.tracker.next_frame\[53\] net1241 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[53\] sky130_fd_sc_hd__dfrtp_1
X_15827_ ag2.body\[269\] net205 _01643_ ag2.body\[261\] vssd1 vssd1 vccd1 vccd1 _01071_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__14074__A1 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19595_ clknet_leaf_119_clk net2448 net1390 vssd1 vssd1 vccd1 vccd1 control.body\[793\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14074__B2 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14866__A net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19265__RESET_B net1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15758_ _05212_ net60 vssd1 vssd1 vccd1 vccd1 _01636_ sky130_fd_sc_hd__nor2_2
X_18546_ clknet_leaf_135_clk _00072_ net1299 vssd1 vssd1 vccd1 vccd1 img_gen.updater.commands.count\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12085__B1 net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19549__CLK clknet_leaf_115_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18057__B _03574_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11832__B1 net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14709_ net1030 _04073_ _04074_ net1010 _08864_ vssd1 vssd1 vccd1 vccd1 _08870_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_64_2280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15689_ ag2.body\[387\] net140 _01616_ ag2.body\[379\] vssd1 vssd1 vccd1 vccd1 _00949_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_75_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18477_ net1512 net1506 vssd1 vssd1 vccd1 vccd1 _00008_ sky130_fd_sc_hd__or2_1
XANTENNA__15023__B1 _01555_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12817__C net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_2144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17428_ ag2.body\[117\] net707 net713 ag2.body\[116\] vssd1 vssd1 vccd1 vccd1 _03107_
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_12_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_2155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16771__B1 net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_962 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_2166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10618__B net1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18573__CLK clknet_leaf_15_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16292__S net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17359_ net1044 net1043 _03006_ _03037_ vssd1 vssd1 vccd1 vccd1 _03038_ sky130_fd_sc_hd__o31ai_1
XANTENNA__18073__A net42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09695__A ag2.body\[71\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20370_ clknet_leaf_22_clk _01257_ net1361 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[6\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_77_2663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_77_2674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload40 clknet_leaf_127_clk vssd1 vssd1 vccd1 vccd1 clkload40/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload51 clknet_leaf_33_clk vssd1 vssd1 vccd1 vccd1 clkload51/Y sky130_fd_sc_hd__inv_12
XTAP_TAPCELL_ROW_77_2685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19029_ clknet_leaf_2_clk img_gen.tracker.next_frame\[467\] net1247 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[467\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_101_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkload62 clknet_leaf_51_clk vssd1 vssd1 vccd1 vccd1 clkload62/Y sky130_fd_sc_hd__inv_6
XANTENNA__11548__A_N _06511_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20605__1537 vssd1 vssd1 vccd1 vccd1 _20605__1537/HI net1537 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_73_2538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload73 clknet_leaf_114_clk vssd1 vssd1 vccd1 vccd1 clkload73/Y sky130_fd_sc_hd__inv_8
XANTENNA__10634__A net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_2084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_2095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload84 clknet_leaf_125_clk vssd1 vssd1 vccd1 vccd1 clkload84/Y sky130_fd_sc_hd__inv_8
XFILLER_0_11_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkload95 clknet_leaf_91_clk vssd1 vssd1 vccd1 vccd1 clkload95/Y sky130_fd_sc_hd__inv_12
XFILLER_0_41_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10353__B net1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18520__B net9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08994_ ag2.body\[91\] vssd1 vssd1 vccd1 vccd1 _04019_ sky130_fd_sc_hd__inv_2
XANTENNA__14837__B1 _08852_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10571__B1 _05543_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1018_A net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout380_A net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09859__A3 _04420_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16975__B net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11184__B net1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09615_ net1049 control.body\[807\] vssd1 vssd1 vccd1 vccd1 _04588_ sky130_fd_sc_hd__xor2_1
XANTENNA_fanout645_A net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14776__A net1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11752__X _06724_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13680__A _04238_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09546_ net909 net904 vssd1 vssd1 vccd1 vccd1 _04519_ sky130_fd_sc_hd__and2_4
XANTENNA__12076__B1 net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11823__B1 net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_4560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout812_A net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09477_ ag2.body\[466\] net1175 vssd1 vssd1 vccd1 vccd1 _04450_ sky130_fd_sc_hd__xor2_1
XANTENNA__18916__CLK clknet_leaf_142_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_4571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_4402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15014__B1 _01553_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10809__A net1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_134_4413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1175_X net1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_134_4424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_1181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_1630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_24_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_24_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload1 clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clkload1/Y sky130_fd_sc_hd__clkinvlp_4
X_20637_ net1554 vssd1 vssd1 vccd1 vccd1 gpio_out[32] sky130_fd_sc_hd__buf_2
XANTENNA_fanout600_X net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16055__X _01734_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_24_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11370_ _06267_ _06289_ _06313_ _06342_ vssd1 vssd1 vccd1 vccd1 _06343_ sky130_fd_sc_hd__and4_1
XFILLER_0_46_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20568_ clknet_leaf_107_clk sound_gen.osc1.keepCounting_nxt _00032_ vssd1 vssd1 vccd1
+ vccd1 sound_gen.osc1.keepCounting sky130_fd_sc_hd__dfrtp_1
XFILLER_0_132_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10321_ _05290_ _05291_ _05292_ _05293_ vssd1 vssd1 vccd1 vccd1 _05294_ sky130_fd_sc_hd__a22o_1
XFILLER_0_61_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20499_ clknet_leaf_23_clk _01386_ net1360 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[135\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_128_4217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13040_ img_gen.tracker.frame\[283\] net646 vssd1 vssd1 vccd1 vccd1 _07715_ sky130_fd_sc_hd__and2_1
XANTENNA__09547__A2 _04519_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10252_ net1226 control.body\[784\] vssd1 vssd1 vccd1 vccd1 _05225_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_128_4228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_128_4239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16278__C1 net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1604 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_1456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10183_ ag2.body\[419\] net1156 vssd1 vssd1 vccd1 vccd1 _05156_ sky130_fd_sc_hd__or2_1
XFILLER_0_121_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17327__A ag2.body\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1203 net1214 vssd1 vssd1 vccd1 vccd1 net1203 sky130_fd_sc_hd__buf_4
Xfanout1214 ag2.y\[1\] vssd1 vssd1 vccd1 vccd1 net1214 sky130_fd_sc_hd__clkbuf_4
Xfanout1225 ag2.y\[0\] vssd1 vssd1 vccd1 vccd1 net1225 sky130_fd_sc_hd__clkbuf_4
Xfanout1236 net1237 vssd1 vssd1 vccd1 vccd1 net1236 sky130_fd_sc_hd__clkbuf_2
X_14991_ control.body\[1014\] net151 _01549_ control.body\[1006\] vssd1 vssd1 vccd1
+ vccd1 _00328_ sky130_fd_sc_hd__a22o_1
Xfanout1247 net1250 vssd1 vssd1 vccd1 vccd1 net1247 sky130_fd_sc_hd__buf_2
Xfanout1258 net1260 vssd1 vssd1 vccd1 vccd1 net1258 sky130_fd_sc_hd__clkbuf_4
Xfanout260 net269 vssd1 vssd1 vccd1 vccd1 net260 sky130_fd_sc_hd__buf_2
Xfanout271 _04307_ vssd1 vssd1 vccd1 vccd1 net271 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout1269 net1287 vssd1 vssd1 vccd1 vccd1 net1269 sky130_fd_sc_hd__clkbuf_4
Xfanout282 _07335_ vssd1 vssd1 vccd1 vccd1 net282 sky130_fd_sc_hd__buf_2
X_16730_ _02404_ _02405_ _02408_ net432 vssd1 vssd1 vccd1 vccd1 _02409_ sky130_fd_sc_hd__o211a_1
X_13942_ ag2.body\[84\] net191 _08154_ ag2.body\[76\] vssd1 vssd1 vccd1 vccd1 _00165_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_57_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10314__B1 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout293 net294 vssd1 vssd1 vccd1 vccd1 net293 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11094__B net1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16661_ _02338_ _02339_ net394 vssd1 vssd1 vccd1 vccd1 _02340_ sky130_fd_sc_hd__mux2_1
X_13873_ _07181_ _08138_ _08146_ vssd1 vssd1 vccd1 vccd1 _00104_ sky130_fd_sc_hd__a21o_1
XFILLER_0_9_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15612_ ag2.body\[461\] net124 _01620_ ag2.body\[453\] vssd1 vssd1 vccd1 vccd1 _00879_
+ sky130_fd_sc_hd__a22o_1
X_18400_ _04636_ _04638_ _03827_ vssd1 vssd1 vccd1 vccd1 _03890_ sky130_fd_sc_hd__o21ai_4
X_12824_ net676 _07613_ vssd1 vssd1 vccd1 vccd1 _07614_ sky130_fd_sc_hd__nor2_1
X_16592_ obsg2.obstacleArray\[74\] obsg2.obstacleArray\[75\] net443 vssd1 vssd1 vccd1
+ vccd1 _02271_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20549__CLK clknet_leaf_105_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19380_ clknet_leaf_112_clk _00324_ net1426 vssd1 vssd1 vccd1 vccd1 control.body\[1010\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13803__A1 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13803__B2 net1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18331_ net915 _04636_ vssd1 vssd1 vccd1 vccd1 _03827_ sky130_fd_sc_hd__nand2_1
XANTENNA__11822__B net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15543_ ag2.body\[513\] net160 _01580_ ag2.body\[505\] vssd1 vssd1 vccd1 vccd1 _00819_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11814__B1 net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12755_ net334 _07475_ vssd1 vssd1 vccd1 vccd1 _07581_ sky130_fd_sc_hd__or2_2
XANTENNA__15005__B1 _01552_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18262_ _03410_ _03533_ net48 obsg2.obstacleArray\[128\] vssd1 vssd1 vccd1 vccd1
+ _03770_ sky130_fd_sc_hd__a31o_1
XFILLER_0_84_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11706_ img_gen.tracker.frame\[305\] net606 net551 img_gen.tracker.frame\[308\] _06677_
+ vssd1 vssd1 vccd1 vccd1 _06678_ sky130_fd_sc_hd__o221a_1
XFILLER_0_84_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15474_ ag2.body\[579\] net108 _01604_ ag2.body\[571\] vssd1 vssd1 vccd1 vccd1 _00757_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__16753__B1 net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12686_ net292 _07547_ _07548_ net1732 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[95\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_56_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_96_3239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17213_ ag2.body\[51\] net848 vssd1 vssd1 vccd1 vccd1 _02892_ sky130_fd_sc_hd__xor2_1
X_14425_ net1025 ag2.body\[557\] vssd1 vssd1 vccd1 vccd1 _08586_ sky130_fd_sc_hd__xor2_1
X_18193_ obsg2.obstacleArray\[93\] _03735_ net526 vssd1 vssd1 vccd1 vccd1 _01344_
+ sky130_fd_sc_hd__o21a_1
X_11637_ _06511_ _06596_ _06609_ vssd1 vssd1 vccd1 vccd1 _06610_ sky130_fd_sc_hd__and3b_1
XANTENNA__09786__Y _04759_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16406__A net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17144_ ag2.body\[269\] net707 net699 ag2.body\[270\] _02817_ vssd1 vssd1 vccd1 vccd1
+ _02823_ sky130_fd_sc_hd__a221o_1
XANTENNA__15310__A _04522_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14356_ net982 _04143_ ag2.body\[407\] net792 _08512_ vssd1 vssd1 vccd1 vccd1 _08517_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_123_820 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11568_ _06485_ _06532_ _06535_ _06540_ _06497_ vssd1 vssd1 vccd1 vccd1 _06541_ sky130_fd_sc_hd__a311o_1
XFILLER_0_107_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold708 control.body\[1103\] vssd1 vssd1 vccd1 vccd1 net2270 sky130_fd_sc_hd__dlygate4sd3_1
X_13307_ net280 net297 _07836_ net1989 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[428\]
+ sky130_fd_sc_hd__a22o_1
X_17075_ ag2.body\[28\] net959 vssd1 vssd1 vccd1 vccd1 _02754_ sky130_fd_sc_hd__xor2_1
X_10519_ ag2.body\[96\] net788 net781 ag2.body\[97\] vssd1 vssd1 vccd1 vccd1 _05492_
+ sky130_fd_sc_hd__o22a_1
Xhold719 control.body\[925\] vssd1 vssd1 vccd1 vccd1 net2281 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_126_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14287_ net979 ag2.body\[474\] vssd1 vssd1 vccd1 vccd1 _08448_ sky130_fd_sc_hd__xor2_1
XFILLER_0_0_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11499_ net1217 net1167 vssd1 vssd1 vccd1 vccd1 _06472_ sky130_fd_sc_hd__or2_1
XFILLER_0_123_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16026_ _01683_ _01688_ vssd1 vssd1 vccd1 vccd1 _01705_ sky130_fd_sc_hd__xor2_1
XANTENNA__11269__B net1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13238_ net672 _07808_ vssd1 vssd1 vccd1 vccd1 _07809_ sky130_fd_sc_hd__nor2_1
XANTENNA__15964__B net60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11837__X _06809_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16808__B2 ag2.body\[71\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09962__B net1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13169_ net668 _07775_ vssd1 vssd1 vccd1 vccd1 _07776_ sky130_fd_sc_hd__nor2_1
XANTENNA__14295__A1 net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17977_ net45 _03598_ vssd1 vssd1 vccd1 vccd1 _03599_ sky130_fd_sc_hd__nor2_1
XFILLER_0_40_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11285__A net1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19716_ clknet_leaf_133_clk net2337 net1308 vssd1 vssd1 vccd1 vccd1 control.body\[674\]
+ sky130_fd_sc_hd__dfrtp_1
X_16928_ _04132_ net862 net691 ag2.body\[375\] vssd1 vssd1 vccd1 vccd1 _02607_ sky130_fd_sc_hd__o22a_1
XFILLER_0_46_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_2910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19371__CLK clknet_leaf_102_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_2921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19647_ clknet_leaf_128_clk _00591_ net1329 vssd1 vssd1 vccd1 vccd1 control.body\[749\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__16287__S net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12668__X _07539_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_2331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16859_ _02534_ _02535_ _02536_ _02537_ vssd1 vssd1 vccd1 vccd1 _02538_ sky130_fd_sc_hd__or4_1
XANTENNA__15244__B1 _01578_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_2342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_2807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09400_ sound_gen.osc1.stayCount\[2\] _04342_ net2366 vssd1 vssd1 vccd1 vccd1 _04384_
+ sky130_fd_sc_hd__a21oi_1
XANTENNA__12058__B1 net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15795__A1 ag2.body\[288\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19578_ clknet_leaf_118_clk _00522_ net1388 vssd1 vssd1 vccd1 vccd1 control.body\[808\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_62_2206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_9_Left_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_2217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_2228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_372 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09331_ _04336_ _04339_ vssd1 vssd1 vccd1 vccd1 _01431_ sky130_fd_sc_hd__nor2_1
X_18529_ clknet_leaf_137_clk _00055_ net1298 vssd1 vssd1 vccd1 vccd1 img_gen.updater.commands.cmd_num\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_48_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09474__A1 _04427_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10629__A net1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17536__A2 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17700__A net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09262_ sound_gen.osc1.timer\[1\] _04284_ _04286_ sound_gen.posDetector1.N\[0\] vssd1
+ vssd1 vccd1 vccd1 _04287_ sky130_fd_sc_hd__o22ai_4
XFILLER_0_117_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16744__B1 net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10348__B net1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_79_2725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_79_2736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09193_ ag2.body\[593\] vssd1 vssd1 vccd1 vccd1 _04218_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_79_2747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_1473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout226_A net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20422_ clknet_leaf_35_clk _01309_ net1350 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[58\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__13659__B net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14867__A_N _04947_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16035__B net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12781__A1 net239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20353_ clknet_leaf_139_clk _01244_ net1289 vssd1 vssd1 vccd1 vccd1 img_gen.updater.commands.rR1.rainbowRNG\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1135_A net1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20284_ clknet_leaf_35_clk control.divider.next_count\[5\] net1348 vssd1 vssd1 vccd1
+ vccd1 control.divider.count\[5\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__15874__B net65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18250__B net35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11894__S net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1302_A net1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold13 control.divider.detect.Q\[0\] vssd1 vssd1 vccd1 vccd1 net1575 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold24 control.button3.Q\[0\] vssd1 vssd1 vccd1 vccd1 net1586 sky130_fd_sc_hd__dlygate4sd3_1
X_08977_ ag2.body\[71\] vssd1 vssd1 vccd1 vccd1 _04002_ sky130_fd_sc_hd__inv_2
Xhold35 img_gen.tracker.frame\[377\] vssd1 vssd1 vccd1 vccd1 net1597 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout762_A net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout383_X net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15483__B1 _01605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold46 img_gen.tracker.frame\[100\] vssd1 vssd1 vccd1 vccd1 net1608 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__16680__C1 _02228_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold57 img_gen.tracker.frame\[373\] vssd1 vssd1 vccd1 vccd1 net1619 sky130_fd_sc_hd__dlygate4sd3_1
Xhold68 img_gen.tracker.frame\[6\] vssd1 vssd1 vccd1 vccd1 net1630 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold79 sound_gen.osc1.stayCount\[5\] vssd1 vssd1 vccd1 vccd1 net1641 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_19_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16197__S net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14038__A1 net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout550_X net550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14038__B2 net1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1292_X net1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11482__X _06455_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout648_X net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12049__B1 net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10870_ ag2.body\[534\] net1084 vssd1 vssd1 vccd1 vccd1 _05843_ sky130_fd_sc_hd__or2_1
XFILLER_0_97_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15786__B2 ag2.body\[288\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout41_A _03702_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12738__B _07572_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_1703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09529_ _04487_ _04488_ _04499_ _04500_ vssd1 vssd1 vccd1 vccd1 _04502_ sky130_fd_sc_hd__a22o_1
XFILLER_0_39_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout815_X net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12540_ net338 net329 _07467_ vssd1 vssd1 vccd1 vccd1 _07468_ sky130_fd_sc_hd__or3_1
XFILLER_0_87_1327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10480__C1 net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12471_ _06724_ net382 _07307_ vssd1 vssd1 vccd1 vccd1 _07426_ sky130_fd_sc_hd__and3_1
XFILLER_0_136_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16226__A net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14210_ net1028 ag2.body\[413\] vssd1 vssd1 vccd1 vccd1 _08371_ sky130_fd_sc_hd__xor2_1
XFILLER_0_129_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11422_ net1077 control.body\[854\] vssd1 vssd1 vccd1 vccd1 _06395_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_91_3103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15190_ net2401 net101 _01572_ control.body\[831\] vssd1 vssd1 vccd1 vccd1 _00505_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_65_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11575__A2 net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12772__A1 net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14141_ net981 ag2.body\[170\] vssd1 vssd1 vccd1 vccd1 _08302_ sky130_fd_sc_hd__xor2_1
X_11353_ _06322_ _06323_ _06324_ _06325_ vssd1 vssd1 vccd1 vccd1 _06326_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_39_1507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16660__S net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10304_ net1096 control.body\[701\] vssd1 vssd1 vccd1 vccd1 _05277_ sky130_fd_sc_hd__or2_1
X_14072_ net984 ag2.body\[210\] vssd1 vssd1 vccd1 vccd1 _08233_ sky130_fd_sc_hd__xor2_1
XANTENNA__11089__B net1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11284_ net1111 control.body\[1109\] vssd1 vssd1 vccd1 vccd1 _06257_ sky130_fd_sc_hd__or2_1
XANTENNA__16232__Y _01911_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18160__B net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17900_ net355 _03535_ vssd1 vssd1 vccd1 vccd1 _03536_ sky130_fd_sc_hd__and2_1
X_13023_ img_gen.tracker.frame\[274\] net646 vssd1 vssd1 vccd1 vccd1 _07707_ sky130_fd_sc_hd__and2_1
X_10235_ ag2.body\[326\] net1090 vssd1 vssd1 vccd1 vccd1 _05208_ sky130_fd_sc_hd__or2_1
X_18880_ clknet_leaf_11_clk img_gen.tracker.next_frame\[318\] net1283 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[318\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_89_3032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1000 net1005 vssd1 vssd1 vccd1 vccd1 net1000 sky130_fd_sc_hd__buf_4
XFILLER_0_105_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19394__CLK clknet_leaf_103_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1011 net1014 vssd1 vssd1 vccd1 vccd1 net1011 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_89_3043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1022 net1024 vssd1 vssd1 vccd1 vccd1 net1022 sky130_fd_sc_hd__buf_2
X_17831_ ag2.apple_cord\[2\] net224 _03492_ net685 vssd1 vssd1 vccd1 vccd1 _01225_
+ sky130_fd_sc_hd__a211o_1
Xfanout1033 ag2.randCord\[5\] vssd1 vssd1 vccd1 vccd1 net1033 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_100_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10280__Y _05253_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10166_ ag2.body\[576\] net1220 vssd1 vssd1 vccd1 vccd1 _05139_ sky130_fd_sc_hd__xor2_1
Xfanout1044 ag2.body\[0\] vssd1 vssd1 vccd1 vccd1 net1044 sky130_fd_sc_hd__clkbuf_4
Xfanout1055 net1069 vssd1 vssd1 vccd1 vccd1 net1055 sky130_fd_sc_hd__buf_4
Xfanout1066 net1068 vssd1 vssd1 vccd1 vccd1 net1066 sky130_fd_sc_hd__buf_4
Xfanout1077 net1082 vssd1 vssd1 vccd1 vccd1 net1077 sky130_fd_sc_hd__buf_4
X_17762_ _03084_ _03087_ _03088_ _03110_ vssd1 vssd1 vccd1 vccd1 _03441_ sky130_fd_sc_hd__o31a_4
Xfanout1088 net1092 vssd1 vssd1 vccd1 vccd1 net1088 sky130_fd_sc_hd__buf_4
X_10097_ net1133 control.body\[940\] vssd1 vssd1 vccd1 vccd1 _05070_ sky130_fd_sc_hd__xor2_1
X_14974_ net637 net54 vssd1 vssd1 vccd1 vccd1 _01548_ sky130_fd_sc_hd__nor2_1
X_19501_ clknet_leaf_113_clk _00445_ net1396 vssd1 vssd1 vccd1 vccd1 control.body\[891\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1099 net1101 vssd1 vssd1 vccd1 vccd1 net1099 sky130_fd_sc_hd__buf_4
X_16713_ _02390_ _02391_ net496 vssd1 vssd1 vccd1 vccd1 _02392_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13925_ ag2.body\[69\] net134 _08152_ ag2.body\[61\] vssd1 vssd1 vccd1 vccd1 _00150_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__14029__A1 net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17693_ _03366_ _03367_ _03369_ _03371_ vssd1 vssd1 vccd1 vccd1 _03372_ sky130_fd_sc_hd__a211o_1
XANTENNA__14029__B2 net1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12929__A net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkload4_A clknet_4_9__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19432_ clknet_leaf_111_clk _00376_ net1422 vssd1 vssd1 vccd1 vccd1 control.body\[966\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_134_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16644_ obsg2.obstacleArray\[51\] net450 net391 vssd1 vssd1 vccd1 vccd1 _02323_ sky130_fd_sc_hd__o21a_1
X_13856_ ag2.body\[19\] net116 _08134_ ag2.body\[11\] vssd1 vssd1 vccd1 vccd1 _00099_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__09571__A2_N net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1028 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20604__1536 vssd1 vssd1 vccd1 vccd1 _20604__1536/HI net1536 sky130_fd_sc_hd__conb_1
XFILLER_0_97_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_18_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12807_ net667 _07605_ vssd1 vssd1 vccd1 vccd1 _07606_ sky130_fd_sc_hd__nor2_1
XANTENNA__11552__B net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19363_ clknet_leaf_102_clk _00307_ net1438 vssd1 vssd1 vccd1 vccd1 control.body\[1025\]
+ sky130_fd_sc_hd__dfrtp_1
X_16575_ obsg2.obstacleArray\[119\] net450 net391 _02253_ vssd1 vssd1 vccd1 vccd1
+ _02254_ sky130_fd_sc_hd__o211a_1
X_13787_ img_gen.updater.commands.count\[13\] _08091_ _08094_ _08070_ vssd1 vssd1
+ vccd1 vccd1 _00070_ sky130_fd_sc_hd__o211a_1
X_10999_ _05965_ _05968_ _05970_ _05971_ vssd1 vssd1 vccd1 vccd1 _05972_ sky130_fd_sc_hd__or4_1
XANTENNA__17775__D_N _03453_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11799__C1 net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18314_ net324 track.nextHighScore\[7\] _03798_ vssd1 vssd1 vccd1 vccd1 _03810_ sky130_fd_sc_hd__or3_1
XFILLER_0_123_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12738_ net305 _07572_ vssd1 vssd1 vccd1 vccd1 _07573_ sky130_fd_sc_hd__nor2_1
X_15526_ ag2.body\[529\] net158 _01610_ ag2.body\[521\] vssd1 vssd1 vccd1 vccd1 _00803_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__16726__B1 net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11263__B2 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19294_ clknet_leaf_99_clk _00238_ net1447 vssd1 vssd1 vccd1 vccd1 control.body\[1100\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10168__B net1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18245_ net519 _03761_ vssd1 vssd1 vccd1 vccd1 _01370_ sky130_fd_sc_hd__nor2_1
X_15457_ ag2.body\[596\] net87 _01602_ net2528 vssd1 vssd1 vccd1 vccd1 _00742_ sky130_fd_sc_hd__a22o_1
XANTENNA__14201__A1 net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12669_ net307 _07539_ vssd1 vssd1 vccd1 vccd1 _07540_ sky130_fd_sc_hd__nor2_1
XFILLER_0_115_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14201__B2 net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14408_ net998 _03964_ _08564_ _08565_ _08568_ vssd1 vssd1 vccd1 vccd1 _08569_ sky130_fd_sc_hd__a221o_1
XFILLER_0_113_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18176_ _03614_ net41 vssd1 vssd1 vccd1 vccd1 _03727_ sky130_fd_sc_hd__nor2_1
XFILLER_0_128_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15388_ net2572 net69 _01595_ net2210 vssd1 vssd1 vccd1 vccd1 _00680_ sky130_fd_sc_hd__a22o_1
XFILLER_0_26_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xwire480 _04415_ vssd1 vssd1 vccd1 vccd1 net480 sky130_fd_sc_hd__buf_2
XFILLER_0_0_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14339_ net1015 ag2.body\[614\] vssd1 vssd1 vccd1 vccd1 _08500_ sky130_fd_sc_hd__xor2_1
X_17127_ _04188_ net874 net727 ag2.body\[514\] _02805_ vssd1 vssd1 vccd1 vccd1 _02806_
+ sky130_fd_sc_hd__a221o_1
Xhold505 img_gen.tracker.frame\[541\] vssd1 vssd1 vccd1 vccd1 net2067 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16423__X _02102_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold516 toggle1.bcd_ones\[3\] vssd1 vssd1 vccd1 vccd1 net2078 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_55_2010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold527 img_gen.tracker.frame\[129\] vssd1 vssd1 vccd1 vccd1 net2089 sky130_fd_sc_hd__dlygate4sd3_1
Xhold538 img_gen.tracker.frame\[427\] vssd1 vssd1 vccd1 vccd1 net2100 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17058_ ag2.body\[73\] net734 net855 _04006_ vssd1 vssd1 vccd1 vccd1 _02737_ sky130_fd_sc_hd__a22o_1
XANTENNA__19737__CLK clknet_leaf_132_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15694__B net64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold549 _00425_ vssd1 vssd1 vccd1 vccd1 net2111 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18070__B _03662_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16009_ _01686_ _01687_ vssd1 vssd1 vccd1 vccd1 _01688_ sky130_fd_sc_hd__xnor2_1
XANTENNA__13495__A net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09880_ _04848_ _04849_ _04851_ _04852_ vssd1 vssd1 vccd1 vccd1 _04853_ sky130_fd_sc_hd__a22o_1
XANTENNA__09692__B net1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16257__A2 net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18761__CLK clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15465__B1 _01603_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16662__C1 net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1529 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_2404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18069__Y _03662_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout176_A net183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19117__CLK clknet_leaf_131_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12558__B net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16745__S net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14440__A1 net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout343_A net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14440__B2 net1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1085_A net1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09314_ sound_gen.osc1.count\[4\] _04323_ vssd1 vssd1 vccd1 vccd1 _04331_ sky130_fd_sc_hd__or2_1
XANTENNA__16717__B1 net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09245_ control.body_update.direction\[0\] vssd1 vssd1 vccd1 vccd1 _04270_ sky130_fd_sc_hd__inv_2
XFILLER_0_8_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09867__B net1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout510_A net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16046__A net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_403 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout608_A _06476_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11006__A1 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11006__B2 net1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15940__A1 ag2.body\[162\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09176_ ag2.body\[547\] vssd1 vssd1 vccd1 vccd1 _04201_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10806__B net1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_784 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12754__A1 net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20405_ clknet_leaf_30_clk _01292_ net1338 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[41\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA_fanout1040_X net1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18261__A net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1138_X net1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1517_A net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20336_ clknet_leaf_21_clk _01227_ net1364 vssd1 vssd1 vccd1 vccd1 ag2.apple_cord\[4\]
+ sky130_fd_sc_hd__dfrtp_1
Xoutput14 net14 vssd1 vssd1 vccd1 vccd1 gpio_out[13] sky130_fd_sc_hd__buf_2
Xoutput25 net25 vssd1 vssd1 vccd1 vccd1 gpio_out[23] sky130_fd_sc_hd__buf_2
XANTENNA_fanout977_A ag2.randCord\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout598_X net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20267_ clknet_leaf_36_clk net1574 net1349 vssd1 vssd1 vccd1 vccd1 control.detect2.Q\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10517__B1 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_399 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10020_ ag2.body\[266\] net776 net1066 _04092_ _04992_ vssd1 vssd1 vccd1 vccd1 _04993_
+ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout89_A net90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09922__A2 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11637__B _06596_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20198_ clknet_leaf_54_clk _01142_ net1454 vssd1 vssd1 vccd1 vccd1 ag2.body\[196\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__14259__A1 net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout765_X net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10541__B net1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14259__B2 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15456__B1 _01602_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16653__C1 net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13852__B net55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout932_X net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11971_ img_gen.tracker.frame\[520\] net599 vssd1 vssd1 vccd1 vccd1 _06943_ sky130_fd_sc_hd__or2_1
XANTENNA__17324__B net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15208__B1 _01574_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11653__A net1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13710_ net2398 _04239_ _08050_ vssd1 vssd1 vccd1 vccd1 track.nextHighScore\[0\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10296__A2 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10922_ ag2.body\[461\] net754 net778 ag2.body\[457\] vssd1 vssd1 vccd1 vccd1 _05895_
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_98_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14690_ _08845_ _08849_ _08850_ vssd1 vssd1 vccd1 vccd1 _08851_ sky130_fd_sc_hd__and3_1
XANTENNA__16956__B1 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout44_X net44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13641_ control.divider.count\[14\] control.divider.count\[13\] _07997_ vssd1 vssd1
+ vccd1 vccd1 _08002_ sky130_fd_sc_hd__and3_1
X_10853_ net1096 control.body\[693\] vssd1 vssd1 vccd1 vccd1 _05826_ sky130_fd_sc_hd__xor2_1
XANTENNA__16655__S net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17340__A net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16360_ obsg2.obstacleArray\[8\] obsg2.obstacleArray\[9\] net409 vssd1 vssd1 vccd1
+ vccd1 _02039_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_1061 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13572_ _07933_ _07943_ _07934_ vssd1 vssd1 vccd1 vccd1 _07948_ sky130_fd_sc_hd__a21bo_1
XANTENNA__09989__A2 _04947_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16708__B1 net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10784_ net1169 control.body\[626\] vssd1 vssd1 vccd1 vccd1 _05757_ sky130_fd_sc_hd__xor2_1
XFILLER_0_93_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15311_ net2538 net77 _01588_ control.body\[712\] vssd1 vssd1 vccd1 vccd1 _00610_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12993__A1 net233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12523_ net2032 net650 _07458_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[22\]
+ sky130_fd_sc_hd__and3_1
X_16291_ _01966_ _01969_ net371 vssd1 vssd1 vccd1 vccd1 _01970_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12484__A net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18030_ net45 _03636_ vssd1 vssd1 vccd1 vccd1 _03637_ sky130_fd_sc_hd__nor2_1
XANTENNA__14195__B1 ag2.body\[162\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15242_ net2216 net98 _01578_ control.body\[781\] vssd1 vssd1 vccd1 vccd1 _00551_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__18634__CLK clknet_leaf_131_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12454_ net777 net1167 _07355_ _07380_ vssd1 vssd1 vccd1 vccd1 _07414_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_35_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15931__B2 ag2.body\[161\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10716__B net1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11405_ ag2.body\[569\] net1203 vssd1 vssd1 vccd1 vccd1 _06378_ sky130_fd_sc_hd__xor2_1
XANTENNA__13867__X _08141_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_1478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15173_ _06180_ _06182_ net63 vssd1 vssd1 vccd1 vccd1 _01571_ sky130_fd_sc_hd__o21a_2
XFILLER_0_50_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12385_ img_gen.updater.commands.rR1.rainbowRNG\[2\] net248 _07333_ vssd1 vssd1 vccd1
+ vccd1 _07350_ sky130_fd_sc_hd__a21o_1
XFILLER_0_1_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14124_ net1009 ag2.body\[375\] vssd1 vssd1 vccd1 vccd1 _08285_ sky130_fd_sc_hd__nand2_1
XFILLER_0_65_1466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11336_ net1045 control.body\[663\] vssd1 vssd1 vccd1 vccd1 _06309_ sky130_fd_sc_hd__xor2_1
X_19981_ clknet_leaf_64_clk _00925_ net1475 vssd1 vssd1 vccd1 vccd1 ag2.body\[411\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__09617__A1_N net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12490__Y _07439_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18932_ clknet_leaf_141_clk img_gen.tracker.next_frame\[370\] net1294 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[370\] sky130_fd_sc_hd__dfrtp_1
X_14055_ net970 ag2.body\[35\] vssd1 vssd1 vccd1 vccd1 _08216_ sky130_fd_sc_hd__xor2_1
X_11267_ net640 net634 vssd1 vssd1 vccd1 vccd1 _06240_ sky130_fd_sc_hd__nor2_2
XANTENNA__14204__A net1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13180__C_N _07515_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13170__A1 net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13006_ net262 _07697_ _07698_ net1627 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[265\]
+ sky130_fd_sc_hd__a22o_1
X_10218_ _05180_ _05185_ _05188_ _05190_ vssd1 vssd1 vccd1 vccd1 _05191_ sky130_fd_sc_hd__or4b_2
XFILLER_0_98_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18863_ clknet_leaf_12_clk img_gen.tracker.next_frame\[301\] net1286 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[301\] sky130_fd_sc_hd__dfrtp_1
X_11198_ net1172 control.body\[874\] vssd1 vssd1 vccd1 vccd1 _06171_ sky130_fd_sc_hd__xor2_1
XANTENNA__15447__B1 _01601_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13465__D net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11720__A2 net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17814_ _03477_ _03479_ vssd1 vssd1 vccd1 vccd1 _03481_ sky130_fd_sc_hd__nand2_1
XFILLER_0_20_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10149_ ag2.body\[58\] net1177 vssd1 vssd1 vccd1 vccd1 _05122_ sky130_fd_sc_hd__nand2_1
X_18794_ clknet_leaf_22_clk img_gen.tracker.next_frame\[232\] net1358 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[232\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17745_ _02671_ _02673_ _03151_ vssd1 vssd1 vccd1 vccd1 _03424_ sky130_fd_sc_hd__o21a_1
X_14957_ net893 _04646_ net65 vssd1 vssd1 vccd1 vccd1 _01547_ sky130_fd_sc_hd__and3_2
XANTENNA__17739__A2 _02849_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13908_ ag2.body\[54\] net90 _08150_ ag2.body\[46\] vssd1 vssd1 vccd1 vccd1 _00135_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__16947__B1 net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17676_ _03347_ _03354_ _03348_ _03352_ vssd1 vssd1 vccd1 vccd1 _03355_ sky130_fd_sc_hd__or4b_4
X_14888_ control.body\[1098\] net179 _01539_ net2392 vssd1 vssd1 vccd1 vccd1 _00236_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_134_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19415_ clknet_leaf_103_clk _00359_ net1432 vssd1 vssd1 vccd1 vccd1 control.body\[981\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__17458__A2_N net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16627_ obsg2.obstacleArray\[32\] obsg2.obstacleArray\[33\] net441 vssd1 vssd1 vccd1
+ vccd1 _02306_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13839_ net1045 _08103_ _08105_ _07413_ vssd1 vssd1 vccd1 vccd1 _00087_ sky130_fd_sc_hd__o211a_1
XANTENNA__14422__A1 net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14422__B2 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19346_ clknet_leaf_101_clk net2261 net1443 vssd1 vssd1 vccd1 vccd1 control.body\[1040\]
+ sky130_fd_sc_hd__dfrtp_1
X_16558_ obsg2.obstacleArray\[106\] obsg2.obstacleArray\[107\] net442 vssd1 vssd1
+ vccd1 vccd1 _02237_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18164__A2 net37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_99_Left_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11787__A2 net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12984__A1 net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15509_ ag2.body\[546\] net155 _01608_ ag2.body\[538\] vssd1 vssd1 vccd1 vccd1 _00788_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_45_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19277_ clknet_leaf_97_clk _00221_ net1450 vssd1 vssd1 vccd1 vccd1 control.body\[1115\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_112_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16489_ net401 _02155_ _02154_ net364 vssd1 vssd1 vccd1 vccd1 _02168_ sky130_fd_sc_hd__a211o_1
XANTENNA__10907__A net1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09030_ ag2.body\[177\] vssd1 vssd1 vccd1 vccd1 _04055_ sky130_fd_sc_hd__inv_2
X_18228_ _03670_ _03703_ obsg2.obstacleArray\[111\] vssd1 vssd1 vccd1 vccd1 _03753_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_5_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19879__RESET_B net1415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_1500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_122 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12736__A1 net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17249__X _02928_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18159_ obsg2.obstacleArray\[76\] _03718_ net522 vssd1 vssd1 vccd1 vccd1 _01327_
+ sky130_fd_sc_hd__o21a_1
XANTENNA__12681__X _07546_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09974__Y _04947_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold302 img_gen.tracker.frame\[185\] vssd1 vssd1 vccd1 vccd1 net1864 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09601__A1 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold313 img_gen.tracker.frame\[197\] vssd1 vssd1 vccd1 vccd1 net1875 sky130_fd_sc_hd__dlygate4sd3_1
Xhold324 img_gen.tracker.frame\[547\] vssd1 vssd1 vccd1 vccd1 net1886 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13937__B net61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold335 img_gen.tracker.frame\[264\] vssd1 vssd1 vccd1 vccd1 net1897 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold346 img_gen.tracker.frame\[42\] vssd1 vssd1 vccd1 vccd1 net1908 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14489__A1 net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold357 img_gen.tracker.frame\[487\] vssd1 vssd1 vccd1 vccd1 net1919 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14489__B2 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09932_ ag2.body\[24\] net1222 vssd1 vssd1 vccd1 vccd1 _04905_ sky130_fd_sc_hd__and2b_1
X_20121_ clknet_leaf_80_clk _01065_ net1487 vssd1 vssd1 vccd1 vccd1 ag2.body\[279\]
+ sky130_fd_sc_hd__dfrtp_2
Xhold368 img_gen.tracker.frame\[470\] vssd1 vssd1 vccd1 vccd1 net1930 sky130_fd_sc_hd__dlygate4sd3_1
Xhold379 img_gen.tracker.frame\[140\] vssd1 vssd1 vccd1 vccd1 net1941 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14114__A net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout804 net805 vssd1 vssd1 vccd1 vccd1 net804 sky130_fd_sc_hd__buf_4
Xfanout815 net816 vssd1 vssd1 vccd1 vccd1 net815 sky130_fd_sc_hd__buf_4
XANTENNA__12560__C net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout826 net827 vssd1 vssd1 vccd1 vccd1 net826 sky130_fd_sc_hd__clkbuf_4
X_20052_ clknet_leaf_72_clk _00996_ net1503 vssd1 vssd1 vccd1 vccd1 ag2.body\[338\]
+ sky130_fd_sc_hd__dfrtp_4
X_09863_ ag2.body\[157\] net1113 vssd1 vssd1 vccd1 vccd1 _04836_ sky130_fd_sc_hd__or2_1
Xfanout837 net839 vssd1 vssd1 vccd1 vccd1 net837 sky130_fd_sc_hd__buf_4
XANTENNA__11457__B net1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout848 net857 vssd1 vssd1 vccd1 vccd1 net848 sky130_fd_sc_hd__buf_4
XANTENNA_fanout293_A net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout859 net867 vssd1 vssd1 vccd1 vccd1 net859 sky130_fd_sc_hd__buf_2
Xhold1002 control.body\[806\] vssd1 vssd1 vccd1 vccd1 net2564 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11711__A2 net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1013 control.body\[944\] vssd1 vssd1 vccd1 vccd1 net2575 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1000_A net1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15989__A1 ag2.body\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1024 control.body\[882\] vssd1 vssd1 vccd1 vccd1 net2586 sky130_fd_sc_hd__dlygate4sd3_1
X_09794_ net1110 control.body\[965\] vssd1 vssd1 vccd1 vccd1 _04767_ sky130_fd_sc_hd__xor2_1
Xhold1035 control.body\[931\] vssd1 vssd1 vccd1 vccd1 net2597 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_119_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1046 control.body\[838\] vssd1 vssd1 vccd1 vccd1 net2608 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_84_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1057 control.body\[1065\] vssd1 vssd1 vccd1 vccd1 net2619 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1068 control.body\[955\] vssd1 vssd1 vccd1 vccd1 net2630 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1079 sound_gen.dac1.dacCount\[3\] vssd1 vssd1 vccd1 vccd1 net2641 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout558_A net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_1504 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__20559__Q net26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09214__Y _04239_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16938__B1 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17431__Y _03110_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout725_A _04264_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17798__C net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15610__B1 _01620_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout346_X net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1088_X net1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09878__A ag2.body\[166\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18657__CLK clknet_leaf_131_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11227__B2 net1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_1268 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11778__A2 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_2_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16166__A1 net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10817__A net1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09228_ control.body\[1051\] vssd1 vssd1 vccd1 vccd1 _04253_ sky130_fd_sc_hd__inv_2
XFILLER_0_90_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09159_ ag2.body\[504\] vssd1 vssd1 vccd1 vccd1 _04184_ sky130_fd_sc_hd__inv_2
XANTENNA__16063__X _01742_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_9_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12170_ img_gen.tracker.frame\[420\] net617 net544 img_gen.tracker.frame\[426\] _07141_
+ vssd1 vssd1 vccd1 vccd1 _07142_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_9_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17319__B net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout882_X net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20603__1535 vssd1 vssd1 vccd1 vccd1 _20603__1535/HI net1535 sky130_fd_sc_hd__conb_1
X_11121_ net1171 control.body\[866\] vssd1 vssd1 vccd1 vccd1 _06094_ sky130_fd_sc_hd__or2_1
XANTENNA__11950__A2 net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20319_ clknet_leaf_44_clk _01215_ net1378 vssd1 vssd1 vccd1 vccd1 obsg2.randCord\[4\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_25_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_1330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14024__A net980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold880 _00661_ vssd1 vssd1 vccd1 vccd1 net2442 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11000__X _05973_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold891 control.body\[673\] vssd1 vssd1 vccd1 vccd1 net2453 sky130_fd_sc_hd__dlygate4sd3_1
X_11052_ ag2.body\[384\] net784 net763 ag2.body\[388\] _06021_ vssd1 vssd1 vccd1 vccd1
+ _06025_ sky130_fd_sc_hd__a221o_1
XANTENNA__10271__B net1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10003_ net1072 control.body\[734\] vssd1 vssd1 vccd1 vccd1 _04976_ sky130_fd_sc_hd__or2_1
XANTENNA__11702__A2 _06644_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15860_ ag2.body\[235\] net175 _01646_ ag2.body\[227\] vssd1 vssd1 vccd1 vccd1 _01101_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__20036__RESET_B net1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16641__A2 net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14811_ net1037 ag2.body\[380\] vssd1 vssd1 vccd1 vccd1 _01482_ sky130_fd_sc_hd__xor2_1
X_15791_ ag2.body\[301\] net209 _01639_ ag2.body\[293\] vssd1 vssd1 vccd1 vccd1 _01039_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__14652__A1 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19432__CLK clknet_leaf_111_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12112__C1 _06647_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14652__B2 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17530_ ag2.body\[273\] net873 vssd1 vssd1 vccd1 vccd1 _03209_ sky130_fd_sc_hd__nand2_1
X_14742_ net1012 _04117_ _08900_ _08901_ _08902_ vssd1 vssd1 vccd1 vccd1 _08903_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_98_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11954_ net572 _06925_ _06923_ net473 vssd1 vssd1 vccd1 vccd1 _06926_ sky130_fd_sc_hd__a211o_1
XANTENNA__16929__B1 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10905_ net1095 control.body\[677\] vssd1 vssd1 vccd1 vccd1 _05878_ sky130_fd_sc_hd__xor2_1
X_17461_ _03134_ _03139_ vssd1 vssd1 vccd1 vccd1 _03140_ sky130_fd_sc_hd__or2_1
X_14673_ net1000 ag2.body\[384\] vssd1 vssd1 vccd1 vccd1 _08834_ sky130_fd_sc_hd__nand2_1
XFILLER_0_19_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_120_3972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11885_ net1216 net1191 img_gen.tracker.frame\[25\] vssd1 vssd1 vccd1 vccd1 _06857_
+ sky130_fd_sc_hd__or3_1
XFILLER_0_135_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_120_3983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_120_3994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15601__B1 _01619_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19200_ clknet_leaf_53_clk _00144_ net1455 vssd1 vssd1 vccd1 vccd1 ag2.body\[63\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__13802__S net1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13624_ control.divider.count\[7\] control.divider.count\[6\] _07985_ control.divider.count\[8\]
+ vssd1 vssd1 vccd1 vccd1 _07991_ sky130_fd_sc_hd__a31o_1
X_16412_ obsg2.obstacleArray\[102\] net452 vssd1 vssd1 vccd1 vccd1 _02091_ sky130_fd_sc_hd__or2_1
X_10836_ ag2.body\[304\] net1236 vssd1 vssd1 vccd1 vccd1 _05809_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_101_3393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17392_ ag2.body\[505\] net874 vssd1 vssd1 vccd1 vccd1 _03071_ sky130_fd_sc_hd__xor2_1
XANTENNA__19582__CLK clknet_leaf_118_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18146__A2 _03570_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19131_ clknet_leaf_140_clk img_gen.tracker.next_frame\[569\] net1297 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[569\] sky130_fd_sc_hd__dfrtp_1
X_16343_ obsg2.obstacleArray\[92\] obsg2.obstacleArray\[93\] net408 vssd1 vssd1 vccd1
+ vccd1 _02022_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16157__A1 _01742_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13555_ ssdec1.in\[2\] ssdec1.in\[3\] _07931_ vssd1 vssd1 vccd1 vccd1 _07937_ sky130_fd_sc_hd__and3_1
XFILLER_0_137_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10767_ _04238_ _04946_ _05517_ vssd1 vssd1 vccd1 vccd1 _05740_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_109_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12506_ net387 net339 _07448_ vssd1 vssd1 vccd1 vccd1 _07449_ sky130_fd_sc_hd__or3_1
XANTENNA__19972__RESET_B net1470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16274_ obsg2.obstacleArray\[24\] obsg2.obstacleArray\[25\] net411 vssd1 vssd1 vccd1
+ vccd1 _01953_ sky130_fd_sc_hd__mux2_1
X_19062_ clknet_leaf_9_clk img_gen.tracker.next_frame\[500\] net1274 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[500\] sky130_fd_sc_hd__dfrtp_1
X_13486_ net2087 net644 _07906_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[537\]
+ sky130_fd_sc_hd__and3_1
XFILLER_0_129_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10698_ _04471_ net634 vssd1 vssd1 vccd1 vccd1 _05671_ sky130_fd_sc_hd__nor2_2
XANTENNA__12718__A1 net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18013_ net432 net462 net495 net482 vssd1 vssd1 vccd1 vccd1 _03624_ sky130_fd_sc_hd__and4_1
X_15225_ net2564 net93 _01576_ control.body\[798\] vssd1 vssd1 vccd1 vccd1 _00536_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__19901__RESET_B net1464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12437_ net1192 _07380_ _06490_ vssd1 vssd1 vccd1 vccd1 _07398_ sky130_fd_sc_hd__a21oi_1
XANTENNA__17106__B1 net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10729__B1 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_114_3787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_114_3798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19219__RESET_B net1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15156_ net2276 net105 _01569_ control.body\[848\] vssd1 vssd1 vccd1 vccd1 _00474_
+ sky130_fd_sc_hd__a22o_1
X_12368_ img_gen.updater.commands.rR1.rainbowRNG\[1\] net248 _07333_ vssd1 vssd1 vccd1
+ vccd1 _07334_ sky130_fd_sc_hd__a21o_1
XFILLER_0_61_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17229__B net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12661__B net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14107_ _08263_ _08265_ _08267_ vssd1 vssd1 vccd1 vccd1 _08268_ sky130_fd_sc_hd__or3b_2
XANTENNA__11941__A2 net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11319_ ag2.body\[553\] net778 net768 ag2.body\[555\] _06291_ vssd1 vssd1 vccd1 vccd1
+ _06292_ sky130_fd_sc_hd__a221o_1
X_19964_ clknet_leaf_62_clk _00908_ net1469 vssd1 vssd1 vccd1 vccd1 ag2.body\[426\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__10462__A _04686_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15087_ net2269 net147 _01562_ net2390 vssd1 vssd1 vccd1 vccd1 _00412_ sky130_fd_sc_hd__a22o_1
XANTENNA__15132__A2 net107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12299_ _07223_ _07263_ vssd1 vssd1 vccd1 vccd1 _07266_ sky130_fd_sc_hd__and2b_1
XANTENNA__13143__A1 net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14038_ net991 _04180_ _04183_ net1011 vssd1 vssd1 vccd1 vccd1 _08199_ sky130_fd_sc_hd__o22a_1
X_18915_ clknet_leaf_3_clk img_gen.tracker.next_frame\[353\] net1258 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[353\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__11277__B net1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10181__B net1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19895_ clknet_leaf_86_clk _00839_ net1462 vssd1 vssd1 vccd1 vccd1 ag2.body\[501\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_38_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16617__C1 net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18846_ clknet_leaf_4_clk img_gen.tracker.next_frame\[284\] net1259 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[284\] sky130_fd_sc_hd__dfrtp_1
X_18777_ clknet_leaf_16_clk img_gen.tracker.next_frame\[215\] net1320 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[215\] sky130_fd_sc_hd__dfrtp_1
X_15989_ ag2.body\[2\] _01659_ _01662_ _01672_ vssd1 vssd1 vccd1 vccd1 _01204_ sky130_fd_sc_hd__o22a_1
XANTENNA__15840__B1 _01644_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17728_ obsg2.obstacleArray\[139\] net502 net488 obsg2.obstacleArray\[138\] vssd1
+ vssd1 vccd1 vccd1 _03407_ sky130_fd_sc_hd__a22o_1
XFILLER_0_76_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17899__B _03533_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19925__CLK clknet_leaf_51_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12539__D net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17659_ ag2.body\[106\] net866 vssd1 vssd1 vccd1 vccd1 _03338_ sky130_fd_sc_hd__or2_1
XANTENNA__18076__A net43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11209__A1 _04446_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12957__A1 net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19329_ clknet_leaf_103_clk _00273_ net1433 vssd1 vssd1 vccd1 vccd1 control.body\[1071\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11740__B net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16148__A1 net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_572 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14109__A net997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout139_A net144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17896__B2 _03519_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09013_ ag2.body\[141\] vssd1 vssd1 vccd1 vccd1 _04038_ sky130_fd_sc_hd__inv_2
XFILLER_0_85_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10924__X _05897_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout306_A net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14580__A1_N net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11917__C1 net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1048_A net1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold110 img_gen.tracker.frame\[126\] vssd1 vssd1 vccd1 vccd1 net1672 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_130_4290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold121 img_gen.tracker.frame\[469\] vssd1 vssd1 vccd1 vccd1 net1683 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__17139__B net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold132 img_gen.tracker.frame\[219\] vssd1 vssd1 vccd1 vccd1 net1694 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_1_clk_A clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold143 img_gen.tracker.frame\[496\] vssd1 vssd1 vccd1 vccd1 net1705 sky130_fd_sc_hd__dlygate4sd3_1
Xhold154 img_gen.tracker.frame\[139\] vssd1 vssd1 vccd1 vccd1 net1716 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_125_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold165 img_gen.tracker.frame\[348\] vssd1 vssd1 vccd1 vccd1 net1727 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09209__Y _04234_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold176 img_gen.tracker.frame\[421\] vssd1 vssd1 vccd1 vccd1 net1738 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1215_A net1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout601 net602 vssd1 vssd1 vccd1 vccd1 net601 sky130_fd_sc_hd__clkbuf_4
Xhold187 img_gen.tracker.frame\[53\] vssd1 vssd1 vccd1 vccd1 net1749 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_1612 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16978__B net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20104_ clknet_leaf_79_clk _01048_ net1489 vssd1 vssd1 vccd1 vccd1 ag2.body\[294\]
+ sky130_fd_sc_hd__dfrtp_4
Xhold198 img_gen.tracker.frame\[237\] vssd1 vssd1 vccd1 vccd1 net1760 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout612 _06475_ vssd1 vssd1 vccd1 vccd1 net612 sky130_fd_sc_hd__clkbuf_4
X_09915_ _04885_ _04886_ _04887_ net634 vssd1 vssd1 vccd1 vccd1 _04888_ sky130_fd_sc_hd__or4b_1
XFILLER_0_121_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16209__A_N net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout623 net625 vssd1 vssd1 vccd1 vccd1 net623 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11145__B1 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout634 _04697_ vssd1 vssd1 vccd1 vccd1 net634 sky130_fd_sc_hd__buf_4
XANTENNA__14779__A net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout645 net654 vssd1 vssd1 vccd1 vccd1 net645 sky130_fd_sc_hd__buf_2
XANTENNA_fanout675_A net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13685__A2 net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout656 net657 vssd1 vssd1 vccd1 vccd1 net656 sky130_fd_sc_hd__buf_1
XANTENNA__13683__A _04944_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20035_ clknet_leaf_67_clk _00979_ net1495 vssd1 vssd1 vccd1 vccd1 ag2.body\[353\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_95_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout667 net669 vssd1 vssd1 vccd1 vccd1 net667 sky130_fd_sc_hd__clkbuf_4
X_09846_ net1133 control.body\[972\] vssd1 vssd1 vccd1 vccd1 _04819_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout1003_X net1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout678 net681 vssd1 vssd1 vccd1 vccd1 net678 sky130_fd_sc_hd__clkbuf_4
Xfanout689 net695 vssd1 vssd1 vccd1 vccd1 net689 sky130_fd_sc_hd__buf_2
X_09777_ _04745_ _04746_ _04748_ _04749_ vssd1 vssd1 vccd1 vccd1 _04750_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_124_4094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout463_X net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout842_A net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14634__A1 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14634__B2 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_1_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09510__B1 net1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17602__B net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout630_X net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout728_X net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17584__B1 obsg2.randCord\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_1043 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11670_ net1122 net1070 net1094 vssd1 vssd1 vccd1 vccd1 _06642_ sky130_fd_sc_hd__o21a_4
XFILLER_0_49_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10671__A2 _04984_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_347 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12948__A1 net246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_137_4488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10621_ ag2.body\[52\] net1121 vssd1 vssd1 vccd1 vccd1 _05594_ sky130_fd_sc_hd__or2_1
XFILLER_0_119_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_4499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_712 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09813__A1 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09813__B2 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13340_ net249 _07848_ _07849_ net1599 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[448\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_134_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10552_ _05513_ _05514_ _05522_ _05523_ vssd1 vssd1 vccd1 vccd1 _05525_ sky130_fd_sc_hd__a22o_1
XANTENNA__17887__A1 _03521_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10266__B _05238_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17975__D net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_715 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_592 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13271_ net257 _07821_ _07822_ net1814 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[406\]
+ sky130_fd_sc_hd__a22o_1
X_10483_ ag2.body\[588\] net1120 vssd1 vssd1 vccd1 vccd1 _05456_ sky130_fd_sc_hd__xnor2_1
XANTENNA__12762__A net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14306__X _08467_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15010_ control.body\[999\] net166 _01552_ control.body\[991\] vssd1 vssd1 vccd1
+ vccd1 _00345_ sky130_fd_sc_hd__a22o_1
XFILLER_0_121_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12222_ img_gen.updater.commands.count\[6\] img_gen.updater.commands.count\[5\] _07191_
+ img_gen.updater.commands.count\[9\] img_gen.updater.commands.count\[8\] vssd1 vssd1
+ vccd1 vccd1 _07192_ sky130_fd_sc_hd__a311o_1
X_20301__1519 vssd1 vssd1 vccd1 vccd1 _20301__1519/HI net1519 sky130_fd_sc_hd__conb_1
XFILLER_0_66_1572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_1545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12481__B net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_735 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13069__S _07726_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12153_ net558 _07124_ _07122_ vssd1 vssd1 vccd1 vccd1 _07125_ sky130_fd_sc_hd__a21o_1
XANTENNA__16311__A1 net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13125__A1 net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11104_ _06067_ _06073_ _06074_ _06076_ vssd1 vssd1 vccd1 vccd1 _06077_ sky130_fd_sc_hd__and4_1
XANTENNA__11097__B net1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16961_ ag2.body\[293\] net952 vssd1 vssd1 vccd1 vccd1 _02640_ sky130_fd_sc_hd__or2_1
X_12084_ img_gen.tracker.frame\[327\] net611 net594 img_gen.tracker.frame\[333\] vssd1
+ vssd1 vccd1 vccd1 _07056_ sky130_fd_sc_hd__a22o_1
XANTENNA__16240__Y _01919_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1171 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18700_ clknet_leaf_9_clk img_gen.tracker.next_frame\[138\] net1274 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[138\] sky130_fd_sc_hd__dfrtp_1
X_15912_ ag2.body\[185\] net131 _01652_ ag2.body\[177\] vssd1 vssd1 vccd1 vccd1 _01147_
+ sky130_fd_sc_hd__a22o_1
X_11035_ net1159 control.body\[1043\] vssd1 vssd1 vccd1 vccd1 _06008_ sky130_fd_sc_hd__nand2b_1
X_19680_ clknet_leaf_136_clk _00624_ net1384 vssd1 vssd1 vccd1 vccd1 control.body\[718\]
+ sky130_fd_sc_hd__dfrtp_1
X_16892_ ag2.body\[214\] net942 vssd1 vssd1 vccd1 vccd1 _02571_ sky130_fd_sc_hd__xor2_1
XFILLER_0_99_1392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16075__B1 net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18631_ clknet_leaf_145_clk img_gen.tracker.next_frame\[69\] net1242 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[69\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15843_ ag2.body\[252\] net175 _01644_ ag2.body\[244\] vssd1 vssd1 vccd1 vccd1 _01086_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_107_3580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15822__B1 _01643_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_3591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18562_ clknet_leaf_15_clk img_gen.tracker.next_frame\[0\] net1278 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[0\] sky130_fd_sc_hd__dfrtp_1
X_15774_ ag2.body\[318\] net209 _01637_ ag2.body\[310\] vssd1 vssd1 vccd1 vccd1 _01024_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_99_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12986_ net665 _07688_ vssd1 vssd1 vccd1 vccd1 _07689_ sky130_fd_sc_hd__nor2_1
XFILLER_0_86_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_103_3455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12100__A2 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_103_3466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17513_ ag2.body\[587\] net715 net688 ag2.body\[591\] vssd1 vssd1 vccd1 vccd1 _03192_
+ sky130_fd_sc_hd__a22o_1
X_14725_ net1033 ag2.body\[117\] vssd1 vssd1 vccd1 vccd1 _08886_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_103_3477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_223 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18493_ net1516 net1510 vssd1 vssd1 vccd1 vccd1 _00024_ sky130_fd_sc_hd__or2_1
X_11937_ img_gen.tracker.frame\[187\] net548 _06908_ net574 vssd1 vssd1 vccd1 vccd1
+ _06909_ sky130_fd_sc_hd__o211a_1
XANTENNA__17512__B net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17444_ ag2.body\[376\] net884 vssd1 vssd1 vccd1 vccd1 _03123_ sky130_fd_sc_hd__xor2_1
X_14656_ net839 ag2.body\[145\] ag2.body\[146\] net829 _08816_ vssd1 vssd1 vccd1 vccd1
+ _08817_ sky130_fd_sc_hd__o221a_1
X_11868_ img_gen.tracker.frame\[268\] net604 net587 img_gen.tracker.frame\[274\] _06839_
+ vssd1 vssd1 vccd1 vccd1 _06840_ sky130_fd_sc_hd__o221a_1
XFILLER_0_55_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18119__A2 net38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12656__B _07532_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16128__B net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12939__A1 net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13607_ control.divider.count\[1\] control.divider.count\[0\] net220 vssd1 vssd1
+ vccd1 vccd1 _07981_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_83_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10819_ net751 control.body\[1094\] net742 vssd1 vssd1 vccd1 vccd1 _05792_ sky130_fd_sc_hd__a21o_1
XFILLER_0_55_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17375_ _03006_ _03046_ vssd1 vssd1 vccd1 vccd1 _03054_ sky130_fd_sc_hd__xor2_1
XFILLER_0_6_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14587_ net845 ag2.body\[80\] ag2.body\[84\] net815 vssd1 vssd1 vccd1 vccd1 _08748_
+ sky130_fd_sc_hd__a22o_1
X_11799_ _06661_ _06767_ _06768_ _06770_ net386 vssd1 vssd1 vccd1 vccd1 _06771_ sky130_fd_sc_hd__a311o_1
XFILLER_0_3_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10821__A_N net1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19114_ clknet_leaf_141_clk img_gen.tracker.next_frame\[552\] net1295 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[552\] sky130_fd_sc_hd__dfrtp_1
X_16326_ obsg2.obstacleArray\[72\] net406 vssd1 vssd1 vccd1 vccd1 _02005_ sky130_fd_sc_hd__or2_1
XFILLER_0_137_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_3849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13538_ net226 _07925_ _07926_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[569\]
+ sky130_fd_sc_hd__o21bai_1
XFILLER_0_55_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10176__B net1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19045_ clknet_leaf_10_clk img_gen.tracker.next_frame\[483\] net1275 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[483\] sky130_fd_sc_hd__dfrtp_1
X_16257_ obsg2.obstacleArray\[57\] net413 _01935_ net419 vssd1 vssd1 vccd1 vccd1 _01936_
+ sky130_fd_sc_hd__o211a_1
XANTENNA__09965__B net1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13469_ net281 _07898_ _07899_ net1656 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[527\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_113_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_11_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20305__CLK clknet_leaf_37_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12167__A2 net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15208_ net2345 net94 _01574_ control.body\[815\] vssd1 vssd1 vccd1 vccd1 _00521_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_45_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13487__B net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16188_ obsg2.obstacleArray\[48\] obsg2.obstacleArray\[49\] net422 vssd1 vssd1 vccd1
+ vccd1 _01867_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11914__A2 net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17527__X _03206_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11288__A net1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15139_ net2655 net105 _01567_ net2311 vssd1 vssd1 vccd1 vccd1 _00459_ sky130_fd_sc_hd__a22o_1
XANTENNA__09981__A net1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19947_ clknet_leaf_45_clk _00891_ net1382 vssd1 vssd1 vccd1 vccd1 ag2.body\[441\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__16853__A2 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_2477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_2488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09700_ ag2.body\[67\] net1162 vssd1 vssd1 vccd1 vccd1 _04673_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_71_2499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19878_ clknet_leaf_82_clk _00822_ net1479 vssd1 vssd1 vccd1 vccd1 ag2.body\[516\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__16066__B1 net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16605__A2 net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17802__A1 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09631_ net640 _04603_ _04572_ vssd1 vssd1 vccd1 vccd1 _04604_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_39_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18829_ clknet_leaf_141_clk img_gen.tracker.next_frame\[267\] net1261 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[267\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_88_2996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09562_ _04512_ _04518_ _04522_ _04534_ vssd1 vssd1 vccd1 vccd1 _04535_ sky130_fd_sc_hd__o22a_1
XANTENNA__13008__A net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17422__B net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09493_ ag2.body\[373\] net1104 vssd1 vssd1 vccd1 vccd1 _04466_ sky130_fd_sc_hd__xor2_1
XANTENNA__16369__A1 _01912_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12847__A _07431_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17566__B1 net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout256_A net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17030__A2 net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20602__1534 vssd1 vssd1 vccd1 vccd1 _20602__1534/HI net1534 sky130_fd_sc_hd__conb_1
XFILLER_0_110_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16038__B net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11470__B net1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_870 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout423_A net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_1238 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1165_A net1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_132_4341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20584_ clknet_leaf_107_clk _01441_ _00048_ vssd1 vssd1 vccd1 vccd1 sound_gen.osc1.count\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_132_4352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_132_4363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09875__B net1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_1580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12582__A net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16054__A net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout309_X net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1332_A net1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13355__A1 net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout792_A net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20381__RESET_B net1374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11905__A2 net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11198__A net1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17097__A2 net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1120_X net1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1218_X net1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13107__A1 net237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18845__CLK clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout580_X net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1407 net1409 vssd1 vssd1 vccd1 vccd1 net1407 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11118__B1 _06087_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout420 _01898_ vssd1 vssd1 vccd1 vccd1 net420 sky130_fd_sc_hd__clkbuf_2
Xfanout1418 net1419 vssd1 vssd1 vccd1 vccd1 net1418 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_1431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout431 _01734_ vssd1 vssd1 vccd1 vccd1 net431 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_100_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout678_X net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1429 net1430 vssd1 vssd1 vccd1 vccd1 net1429 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_54_1974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout442 net443 vssd1 vssd1 vccd1 vccd1 net442 sky130_fd_sc_hd__clkbuf_2
XANTENNA__11669__A1 _06639_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout453 net459 vssd1 vssd1 vccd1 vccd1 net453 sky130_fd_sc_hd__clkbuf_4
Xfanout464 net465 vssd1 vssd1 vccd1 vccd1 net464 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_35_1384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout486 net487 vssd1 vssd1 vccd1 vccd1 net486 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_1395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20018_ clknet_leaf_58_clk _00962_ net1471 vssd1 vssd1 vccd1 vccd1 ag2.body\[368\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_6_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout497 net499 vssd1 vssd1 vccd1 vccd1 net497 sky130_fd_sc_hd__buf_4
X_09829_ net1133 control.body\[924\] vssd1 vssd1 vccd1 vccd1 _04802_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout845_X net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18995__CLK clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15804__B1 _01641_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12840_ _06672_ _07531_ vssd1 vssd1 vccd1 vccd1 _07621_ sky130_fd_sc_hd__or2_1
XFILLER_0_69_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17332__B net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12771_ net256 _07588_ _07589_ net1716 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[139\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_69_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12757__A net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14510_ net833 ag2.body\[177\] ag2.body\[178\] net826 _08669_ vssd1 vssd1 vccd1 vccd1
+ _08671_ sky130_fd_sc_hd__a221o_1
X_11722_ img_gen.tracker.frame\[236\] net552 vssd1 vssd1 vccd1 vccd1 _06694_ sky130_fd_sc_hd__or2_1
XFILLER_0_138_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_48_1778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15490_ ag2.body\[561\] net110 _01606_ ag2.body\[553\] vssd1 vssd1 vccd1 vccd1 _00771_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_48_1789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12476__B net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14441_ _08596_ _08598_ _08600_ _08601_ vssd1 vssd1 vccd1 vccd1 _08602_ sky130_fd_sc_hd__or4b_1
XFILLER_0_83_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11653_ net1122 net1070 vssd1 vssd1 vccd1 vccd1 _06626_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_29_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16663__S net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout60 net61 vssd1 vssd1 vccd1 vccd1 net60 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_37_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout71 net79 vssd1 vssd1 vccd1 vccd1 net71 sky130_fd_sc_hd__buf_2
XANTENNA__20328__CLK clknet_leaf_105_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10604_ net1161 control.body\[987\] vssd1 vssd1 vccd1 vccd1 _05577_ sky130_fd_sc_hd__or2_1
XFILLER_0_65_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14372_ net1000 ag2.body\[416\] vssd1 vssd1 vccd1 vccd1 _08533_ sky130_fd_sc_hd__xor2_1
Xfanout82 net83 vssd1 vssd1 vccd1 vccd1 net82 sky130_fd_sc_hd__buf_2
X_17160_ ag2.body\[599\] net928 vssd1 vssd1 vccd1 vccd1 _02839_ sky130_fd_sc_hd__nand2_1
Xfanout93 net100 vssd1 vssd1 vccd1 vccd1 net93 sky130_fd_sc_hd__clkbuf_2
X_11584_ net1144 net595 vssd1 vssd1 vccd1 vccd1 _06557_ sky130_fd_sc_hd__nand2_1
XANTENNA__08970__A ag2.body\[57\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16111_ obsg2.obstacleArray\[70\] obsg2.obstacleArray\[71\] net426 vssd1 vssd1 vccd1
+ vccd1 _01790_ sky130_fd_sc_hd__mux2_1
X_13323_ net665 _07842_ vssd1 vssd1 vccd1 vccd1 _07843_ sky130_fd_sc_hd__nor2_1
XFILLER_0_101_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10535_ net1083 control.body\[918\] vssd1 vssd1 vccd1 vccd1 _05508_ sky130_fd_sc_hd__xor2_1
XFILLER_0_135_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17091_ ag2.body\[298\] net726 net964 _04099_ _02769_ vssd1 vssd1 vccd1 vccd1 _02770_
+ sky130_fd_sc_hd__o221a_1
XANTENNA__12492__A net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_3702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_3178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11600__S net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_94_3189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_3713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12149__A2 net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16042_ net355 net350 _01720_ vssd1 vssd1 vccd1 vccd1 _01721_ sky130_fd_sc_hd__and3_1
X_13254_ net671 _07815_ vssd1 vssd1 vccd1 vccd1 _07816_ sky130_fd_sc_hd__nor2_1
X_10466_ net1109 control.body\[1013\] vssd1 vssd1 vccd1 vccd1 _05439_ sky130_fd_sc_hd__nand2_1
XFILLER_0_126_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12205_ _06634_ _06825_ _06986_ _07147_ _07176_ vssd1 vssd1 vccd1 vccd1 _07177_ sky130_fd_sc_hd__a41o_1
XFILLER_0_86_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13185_ net337 net309 _07612_ vssd1 vssd1 vccd1 vccd1 _07783_ sky130_fd_sc_hd__and3_1
X_10397_ net1110 control.body\[1061\] vssd1 vssd1 vccd1 vccd1 _05370_ sky130_fd_sc_hd__or2_1
XANTENNA__20051__RESET_B net1504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19801_ clknet_leaf_124_clk _00745_ net1405 vssd1 vssd1 vccd1 vccd1 ag2.body\[599\]
+ sky130_fd_sc_hd__dfrtp_4
X_12136_ img_gen.tracker.frame\[495\] net602 net571 vssd1 vssd1 vccd1 vccd1 _07108_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_104_1554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17993_ obsg2.obstacleArray\[19\] _03609_ net533 vssd1 vssd1 vccd1 vccd1 _01270_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_62_1299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19732_ clknet_leaf_133_clk net2227 net1305 vssd1 vssd1 vccd1 vccd1 control.body\[658\]
+ sky130_fd_sc_hd__dfrtp_1
X_16944_ ag2.body\[391\] net931 vssd1 vssd1 vccd1 vccd1 _02623_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_109_3642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12067_ _07001_ _07015_ _07025_ _07038_ net386 vssd1 vssd1 vccd1 vccd1 _07039_ sky130_fd_sc_hd__o221ai_4
XTAP_TAPCELL_ROW_109_3653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11018_ ag2.body\[594\] net1169 vssd1 vssd1 vccd1 vccd1 _05991_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_105_3517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19663_ clknet_leaf_134_clk net2465 net1309 vssd1 vssd1 vccd1 vccd1 control.body\[733\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_105_3528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16875_ ag2.body\[465\] net730 net690 ag2.body\[471\] _02549_ vssd1 vssd1 vccd1 vccd1
+ _02554_ sky130_fd_sc_hd__a221o_1
XANTENNA__16599__A1 net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_3539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1075 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18614_ clknet_leaf_145_clk img_gen.tracker.next_frame\[52\] net1241 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[52\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_56_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15826_ ag2.body\[268\] net201 _01643_ ag2.body\[260\] vssd1 vssd1 vccd1 vccd1 _01070_
+ sky130_fd_sc_hd__a22o_1
X_19594_ clknet_leaf_118_clk _00538_ net1393 vssd1 vssd1 vccd1 vccd1 control.body\[792\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_56_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14074__A2 ag2.body\[213\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14866__B net59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18545_ clknet_leaf_135_clk _00071_ net1299 vssd1 vssd1 vccd1 vccd1 img_gen.updater.commands.count\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_15757_ ag2.body\[335\] net216 _01635_ ag2.body\[327\] vssd1 vssd1 vccd1 vccd1 _01009_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_87_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_138_clk clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_138_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_38_1471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17548__B1 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_83_2860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12667__A net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12969_ net341 _07498_ vssd1 vssd1 vccd1 vccd1 _07681_ sky130_fd_sc_hd__nor2_1
XFILLER_0_34_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19150__CLK clknet_leaf_51_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17012__A2 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14708_ net808 ag2.body\[237\] ag2.body\[239\] net795 _08868_ vssd1 vssd1 vccd1 vccd1
+ _08869_ sky130_fd_sc_hd__a221o_1
XFILLER_0_115_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18476_ net1514 net1508 vssd1 vssd1 vccd1 vccd1 _00007_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_64_2270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15688_ ag2.body\[386\] net136 _01616_ ag2.body\[378\] vssd1 vssd1 vccd1 vccd1 _00948_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_64_2281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17427_ ag2.body\[114\] net729 net720 ag2.body\[115\] _03105_ vssd1 vssd1 vccd1 vccd1
+ _03106_ sky130_fd_sc_hd__o221a_1
XANTENNA__18718__CLK clknet_leaf_142_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_2145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12817__D _07515_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_2156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14639_ net840 ag2.body\[576\] _04210_ net979 _08794_ vssd1 vssd1 vccd1 vccd1 _08800_
+ sky130_fd_sc_hd__a221o_1
XANTENNA__10187__A _05152_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15574__A2 net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_60_2167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09976__A net1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17358_ ag2.body\[4\] net925 _03017_ vssd1 vssd1 vccd1 vccd1 _03037_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_12_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16309_ obsg2.obstacleArray\[105\] net413 _01987_ net418 vssd1 vssd1 vccd1 vccd1
+ _01988_ sky130_fd_sc_hd__o211a_1
XANTENNA__09695__B net1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_372 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17289_ ag2.body\[305\] net736 net694 ag2.body\[311\] vssd1 vssd1 vccd1 vccd1 _02968_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_77_2664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload30 clknet_leaf_135_clk vssd1 vssd1 vccd1 vccd1 clkload30/Y sky130_fd_sc_hd__clkinv_4
XTAP_TAPCELL_ROW_77_2675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19028_ clknet_leaf_1_clk img_gen.tracker.next_frame\[466\] net1246 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[466\] sky130_fd_sc_hd__dfrtp_1
Xclkload41 clknet_leaf_128_clk vssd1 vssd1 vccd1 vccd1 clkload41/Y sky130_fd_sc_hd__clkinv_8
XFILLER_0_71_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_77_2686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_wire479_X net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_754 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload52 clknet_leaf_34_clk vssd1 vssd1 vccd1 vccd1 clkload52/Y sky130_fd_sc_hd__inv_16
Xclkload63 clknet_leaf_52_clk vssd1 vssd1 vccd1 vccd1 clkload63/Y sky130_fd_sc_hd__clkinv_4
XTAP_TAPCELL_ROW_73_2539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload74 clknet_leaf_115_clk vssd1 vssd1 vccd1 vccd1 clkload74/Y sky130_fd_sc_hd__inv_6
XFILLER_0_51_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_2085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18276__A1 net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload85 clknet_leaf_102_clk vssd1 vssd1 vccd1 vccd1 clkload85/X sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_58_2096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkload96 clknet_leaf_94_clk vssd1 vssd1 vccd1 vccd1 clkload96/Y sky130_fd_sc_hd__bufinv_16
XFILLER_0_122_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10020__B1 net1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08993_ ag2.body\[90\] vssd1 vssd1 vccd1 vccd1 _04018_ sky130_fd_sc_hd__inv_2
XFILLER_0_11_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14837__A1 _08475_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10571__A1 net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15218__A _04587_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14122__A net1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09713__B1 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11465__B net1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09859__A4 _04470_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_4020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout373_A net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09614_ net905 _04586_ net636 vssd1 vssd1 vccd1 vccd1 _04587_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_97_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18248__B net35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09545_ _04513_ _04514_ _04515_ _04516_ _04517_ vssd1 vssd1 vccd1 vccd1 _04518_ sky130_fd_sc_hd__a221o_2
X_20300__1518 vssd1 vssd1 vccd1 vccd1 _20300__1518/HI net1518 sky130_fd_sc_hd__conb_1
XFILLER_0_6_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_129_clk clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_129_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout540_A net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout161_X net161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16049__A net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout259_X net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout638_A _04470_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17003__A2 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09476_ ag2.body\[464\] net1223 vssd1 vssd1 vccd1 vccd1 _04449_ sky130_fd_sc_hd__xor2_1
XFILLER_0_91_1495 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_4550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_4403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_4414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_134_4425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10097__A net1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1070_X net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_1631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout426_X net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_1642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09886__A _04446_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20636_ net1553 vssd1 vssd1 vccd1 vccd1 gpio_out[31] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_24_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkload2 clknet_4_4__leaf_clk vssd1 vssd1 vccd1 vccd1 clkload2/X sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_24_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_24_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11051__A2 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20567_ clknet_leaf_43_clk _01426_ net1378 vssd1 vssd1 vccd1 vccd1 obsg2.randCord\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_1266 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10320_ ag2.body\[610\] net1169 vssd1 vssd1 vccd1 vccd1 _05293_ sky130_fd_sc_hd__or2_1
X_20498_ clknet_leaf_22_clk _01385_ net1361 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[134\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_131_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout795_X net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10544__B _04599_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10251_ net1170 control.body\[786\] vssd1 vssd1 vccd1 vccd1 _05224_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_128_4218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1502_X net1502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_4229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_37_1446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16817__A2 net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10182_ ag2.body\[419\] net1154 vssd1 vssd1 vccd1 vccd1 _05155_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_37_1457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17327__B net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_1616 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout962_X net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1204 net1205 vssd1 vssd1 vccd1 vccd1 net1204 sky130_fd_sc_hd__buf_4
Xfanout1215 net1221 vssd1 vssd1 vccd1 vccd1 net1215 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11656__A net1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1226 net1227 vssd1 vssd1 vccd1 vccd1 net1226 sky130_fd_sc_hd__buf_4
XANTENNA__15128__A _05634_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1237 net1238 vssd1 vssd1 vccd1 vccd1 net1237 sky130_fd_sc_hd__buf_4
XFILLER_0_121_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14032__A net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout250 net260 vssd1 vssd1 vccd1 vccd1 net250 sky130_fd_sc_hd__clkbuf_4
X_14990_ net2237 net158 _01549_ control.body\[1005\] vssd1 vssd1 vccd1 vccd1 _00327_
+ sky130_fd_sc_hd__a22o_1
Xfanout1248 net1250 vssd1 vssd1 vccd1 vccd1 net1248 sky130_fd_sc_hd__clkbuf_4
Xfanout261 net264 vssd1 vssd1 vccd1 vccd1 net261 sky130_fd_sc_hd__clkbuf_4
Xfanout1259 net1260 vssd1 vssd1 vccd1 vccd1 net1259 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11375__B net1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout272 _04306_ vssd1 vssd1 vccd1 vccd1 net272 sky130_fd_sc_hd__buf_2
X_13941_ ag2.body\[83\] net197 _08154_ ag2.body\[75\] vssd1 vssd1 vccd1 vccd1 _00164_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_96_1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout283 net285 vssd1 vssd1 vccd1 vccd1 net283 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10314__A1 _04421_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout294 net295 vssd1 vssd1 vccd1 vccd1 net294 sky130_fd_sc_hd__buf_2
XFILLER_0_96_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16660_ obsg2.obstacleArray\[12\] obsg2.obstacleArray\[13\] net443 vssd1 vssd1 vccd1
+ vccd1 _02339_ sky130_fd_sc_hd__mux2_1
XANTENNA__19173__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17242__A2 net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13872_ toggle1.bcd_hundreds\[0\] net434 _08144_ _08022_ vssd1 vssd1 vccd1 vccd1
+ _08146_ sky130_fd_sc_hd__a22o_1
XANTENNA__18158__B net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15611_ ag2.body\[460\] net123 _01620_ ag2.body\[452\] vssd1 vssd1 vccd1 vccd1 _00878_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_92_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_1600 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12823_ net383 net309 _07612_ vssd1 vssd1 vccd1 vccd1 _07613_ sky130_fd_sc_hd__and3_1
X_16591_ net396 _02269_ _02268_ net360 vssd1 vssd1 vccd1 vccd1 _02270_ sky130_fd_sc_hd__a211o_1
XFILLER_0_16_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13803__A2 net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11391__A net1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18330_ _04643_ _08026_ _08028_ vssd1 vssd1 vccd1 vccd1 _03826_ sky130_fd_sc_hd__or3_1
X_15542_ ag2.body\[512\] net188 _01580_ ag2.body\[504\] vssd1 vssd1 vccd1 vccd1 _00818_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__10617__A2 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12754_ net281 _07579_ _07580_ net1955 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[131\]
+ sky130_fd_sc_hd__a22o_1
X_18261_ net519 _03769_ vssd1 vssd1 vccd1 vccd1 _01378_ sky130_fd_sc_hd__nor2_1
X_11705_ img_gen.tracker.frame\[302\] net623 net591 img_gen.tracker.frame\[311\] vssd1
+ vssd1 vccd1 vccd1 _06677_ sky130_fd_sc_hd__o22a_1
XFILLER_0_132_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_117_3900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15556__A2 net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12685_ net267 _07547_ _07548_ net1729 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[94\]
+ sky130_fd_sc_hd__a22o_1
X_15473_ ag2.body\[578\] net111 _01604_ ag2.body\[570\] vssd1 vssd1 vccd1 vccd1 _00756_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_13_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17212_ _03991_ net869 net859 _03992_ vssd1 vssd1 vccd1 vccd1 _02891_ sky130_fd_sc_hd__a22o_1
XFILLER_0_126_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11636_ _06485_ _06605_ _06608_ _06497_ _06601_ vssd1 vssd1 vccd1 vccd1 _06609_ sky130_fd_sc_hd__a311o_1
XANTENNA__09796__A net1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14424_ net1035 ag2.body\[556\] vssd1 vssd1 vccd1 vccd1 _08585_ sky130_fd_sc_hd__xor2_1
X_18192_ _03636_ net41 vssd1 vssd1 vccd1 vccd1 _03735_ sky130_fd_sc_hd__nor2_1
XFILLER_0_65_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_1631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17143_ ag2.body\[269\] net707 net699 ag2.body\[270\] _02818_ vssd1 vssd1 vccd1 vccd1
+ _02822_ sky130_fd_sc_hd__o221ai_1
XFILLER_0_0_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14355_ net833 ag2.body\[401\] ag2.body\[402\] net826 _08515_ vssd1 vssd1 vccd1 vccd1
+ _08516_ sky130_fd_sc_hd__a221o_1
X_11567_ net506 _06536_ _06539_ net475 vssd1 vssd1 vccd1 vccd1 _06540_ sky130_fd_sc_hd__o211a_1
XANTENNA__15310__B net53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13111__A net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10518_ ag2.body\[96\] net788 net1164 _04024_ vssd1 vssd1 vccd1 vccd1 _05491_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_80_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13306_ net255 net297 _07836_ net2100 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[427\]
+ sky130_fd_sc_hd__a22o_1
X_14286_ _08443_ _08444_ _08446_ vssd1 vssd1 vccd1 vccd1 _08447_ sky130_fd_sc_hd__or3_1
X_17074_ ag2.body\[30\] net937 vssd1 vssd1 vccd1 vccd1 _02753_ sky130_fd_sc_hd__xor2_1
Xhold709 _00233_ vssd1 vssd1 vccd1 vccd1 net2271 sky130_fd_sc_hd__dlygate4sd3_1
X_11498_ _06469_ _06470_ net506 vssd1 vssd1 vccd1 vccd1 _06471_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10454__B net1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16025_ _01683_ _01688_ vssd1 vssd1 vccd1 vccd1 _01704_ sky130_fd_sc_hd__or2_1
XFILLER_0_0_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13237_ net382 _07425_ net314 vssd1 vssd1 vccd1 vccd1 _07808_ sky130_fd_sc_hd__and3_1
X_10449_ ag2.body\[455\] net1055 vssd1 vssd1 vccd1 vccd1 _05422_ sky130_fd_sc_hd__nand2_1
XFILLER_0_42_1604 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18627__RESET_B net1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10173__C _05119_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16808__A2 net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13168_ net336 net327 _07508_ vssd1 vssd1 vccd1 vccd1 _07775_ sky130_fd_sc_hd__and3_1
XFILLER_0_23_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20601__1533 vssd1 vssd1 vccd1 vccd1 _20601__1533/HI net1533 sky130_fd_sc_hd__conb_1
XANTENNA__14819__A1 net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14819__B2 net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_41_clk_A clknet_4_7__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11566__A net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12119_ net467 _07090_ net466 vssd1 vssd1 vccd1 vccd1 _07091_ sky130_fd_sc_hd__a21o_1
X_17976_ net298 _03597_ vssd1 vssd1 vccd1 vccd1 _03598_ sky130_fd_sc_hd__nand2_1
XANTENNA__10470__A net1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13099_ net344 _07572_ vssd1 vssd1 vccd1 vccd1 _07742_ sky130_fd_sc_hd__nor2_1
X_19715_ clknet_leaf_132_clk _00659_ net1303 vssd1 vssd1 vccd1 vccd1 control.body\[673\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_100_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16927_ ag2.body\[371\] net717 net691 ag2.body\[375\] vssd1 vssd1 vccd1 vccd1 _02606_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_79_1571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_85_2911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11853__X _06825_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17233__A2 net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19646_ clknet_leaf_128_clk _00590_ net1329 vssd1 vssd1 vccd1 vccd1 control.body\[748\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_66_2321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16858_ ag2.body\[203\] net853 vssd1 vssd1 vccd1 vccd1 _02537_ sky130_fd_sc_hd__xor2_1
XANTENNA_clkbuf_leaf_56_clk_A clknet_4_12__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_2332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_2343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_2808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15809_ ag2.body\[285\] net206 _01641_ ag2.body\[277\] vssd1 vssd1 vccd1 vccd1 _01055_
+ sky130_fd_sc_hd__a22o_1
X_19577_ clknet_leaf_116_clk _00521_ net1387 vssd1 vssd1 vccd1 vccd1 control.body\[823\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16789_ _01700_ _02463_ _02467_ net318 _02462_ vssd1 vssd1 vccd1 vccd1 _02468_ sky130_fd_sc_hd__o311a_1
XANTENNA__12397__A net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_2207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09330_ net2641 _04335_ net2117 vssd1 vssd1 vccd1 vccd1 _04339_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_62_2218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18528_ clknet_leaf_138_clk _00054_ net1292 vssd1 vssd1 vccd1 vccd1 img_gen.updater.commands.cmd_num\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_48_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_2229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1132 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_1300 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09474__A2 _04446_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_80_Left_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09261_ sound_gen.osc1.keepCounting sound_gen.posDetector1.N\[1\] vssd1 vssd1 vccd1
+ vccd1 _04286_ sky130_fd_sc_hd__nand2b_2
X_18459_ _03821_ _03947_ _08035_ vssd1 vssd1 vccd1 vccd1 _03948_ sky130_fd_sc_hd__o21ai_1
XANTENNA__15547__A2 net162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_462 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_2726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09192_ ag2.body\[591\] vssd1 vssd1 vccd1 vccd1 _04217_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_79_2737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_114_clk_A clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20421_ clknet_leaf_37_clk _01308_ net1353 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[57\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_12_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout121_A net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16035__C net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_1586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13021__A net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkload130 clknet_leaf_71_clk vssd1 vssd1 vccd1 vccd1 clkload130/Y sky130_fd_sc_hd__clkinv_8
XFILLER_0_86_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20352_ clknet_leaf_139_clk _01243_ net1289 vssd1 vssd1 vccd1 vccd1 img_gen.updater.commands.rR1.rainbowRNG\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__19046__CLK clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20283_ clknet_leaf_36_clk control.divider.next_count\[4\] net1348 vssd1 vssd1 vccd1
+ vccd1 control.divider.count\[4\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__12860__A net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_129_clk_A clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1030_A net1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1128_A net1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13675__B _07181_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17147__B net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout490_A net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11741__B1 net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout588_A net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold14 control.detect1.Q\[0\] vssd1 vssd1 vccd1 vccd1 net1576 sky130_fd_sc_hd__dlygate4sd3_1
X_08976_ ag2.body\[70\] vssd1 vssd1 vccd1 vccd1 _04001_ sky130_fd_sc_hd__inv_2
XANTENNA__19196__CLK clknet_leaf_53_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold25 sound_gen.dac1.dacCount\[7\] vssd1 vssd1 vccd1 vccd1 net1587 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold36 img_gen.tracker.frame\[225\] vssd1 vssd1 vccd1 vccd1 net1598 sky130_fd_sc_hd__dlygate4sd3_1
Xhold47 img_gen.tracker.frame\[99\] vssd1 vssd1 vccd1 vccd1 net1609 sky130_fd_sc_hd__dlygate4sd3_1
Xhold58 img_gen.tracker.frame\[62\] vssd1 vssd1 vccd1 vccd1 net1620 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__16478__S net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold69 img_gen.tracker.frame\[1\] vssd1 vssd1 vccd1 vccd1 net1631 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout376_X net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout755_A net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17224__A2 net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1508 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11923__B net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout922_A net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout543_X net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_119_Left_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09528_ _04485_ _04486_ _04497_ _04498_ _04490_ vssd1 vssd1 vccd1 vccd1 _04501_ sky130_fd_sc_hd__a221o_1
XFILLER_0_39_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_1704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18185__B1 net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09465__A2 net1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_26_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10539__B net1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09459_ net912 net920 net916 net907 vssd1 vssd1 vccd1 vccd1 _04432_ sky130_fd_sc_hd__a31o_1
XANTENNA_fanout710_X net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout808_X net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1452_X net1452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12470_ _07421_ net334 vssd1 vssd1 vccd1 vccd1 _07425_ sky130_fd_sc_hd__and2_2
XFILLER_0_30_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11421_ net637 _06391_ _06392_ _06393_ vssd1 vssd1 vccd1 vccd1 _06394_ sky130_fd_sc_hd__or4_1
X_20619_ net1562 vssd1 vssd1 vccd1 vccd1 gpio_oeb[31] sky130_fd_sc_hd__buf_2
XFILLER_0_129_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_3104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14140_ net842 ag2.body\[168\] ag2.body\[174\] net800 _08295_ vssd1 vssd1 vccd1 vccd1
+ _08301_ sky130_fd_sc_hd__a221o_1
X_11352_ ag2.body\[445\] net1103 vssd1 vssd1 vccd1 vccd1 _06325_ sky130_fd_sc_hd__or2_1
XFILLER_0_65_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_39_1508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10274__B net1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_128_Left_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_39_1519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11980__B1 net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10303_ net1121 control.body\[700\] vssd1 vssd1 vccd1 vccd1 _05276_ sky130_fd_sc_hd__xor2_1
X_14071_ net814 ag2.body\[212\] ag2.body\[215\] net794 vssd1 vssd1 vccd1 vccd1 _08232_
+ sky130_fd_sc_hd__a22o_1
X_11283_ net1085 control.body\[1110\] vssd1 vssd1 vccd1 vccd1 _06256_ sky130_fd_sc_hd__xor2_1
XANTENNA__14314__X _08475_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19539__CLK clknet_leaf_115_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13022_ net240 _07705_ _07706_ net1815 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[273\]
+ sky130_fd_sc_hd__a22o_1
X_10234_ ag2.body\[327\] net1067 vssd1 vssd1 vccd1 vccd1 _05207_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_89_3033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1001 net1002 vssd1 vssd1 vccd1 vccd1 net1001 sky130_fd_sc_hd__buf_4
Xfanout1012 net1013 vssd1 vssd1 vccd1 vccd1 net1012 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_89_3044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17830_ net824 net224 vssd1 vssd1 vccd1 vccd1 _03492_ sky130_fd_sc_hd__nor2_1
XANTENNA__11386__A net1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10165_ ag2.body\[580\] net1120 vssd1 vssd1 vccd1 vccd1 _05138_ sky130_fd_sc_hd__xor2_1
Xfanout1023 net1024 vssd1 vssd1 vccd1 vccd1 net1023 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_24_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1034 net1035 vssd1 vssd1 vccd1 vccd1 net1034 sky130_fd_sc_hd__buf_4
XANTENNA__20516__CLK clknet_leaf_113_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1045 net1046 vssd1 vssd1 vccd1 vccd1 net1045 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_41_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1056 net1057 vssd1 vssd1 vccd1 vccd1 net1056 sky130_fd_sc_hd__buf_4
X_17761_ _02683_ _02790_ _03120_ _03376_ vssd1 vssd1 vccd1 vccd1 _03440_ sky130_fd_sc_hd__and4_2
XANTENNA__19926__RESET_B net1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1067 net1068 vssd1 vssd1 vccd1 vccd1 net1067 sky130_fd_sc_hd__clkbuf_4
X_10096_ net1204 control.body\[937\] vssd1 vssd1 vccd1 vccd1 _05069_ sky130_fd_sc_hd__xor2_1
XANTENNA__18563__CLK clknet_leaf_15_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14973_ net2618 net157 net51 net2120 vssd1 vssd1 vccd1 vccd1 _00313_ sky130_fd_sc_hd__a22o_1
XFILLER_0_22_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1078 net1079 vssd1 vssd1 vccd1 vccd1 net1078 sky130_fd_sc_hd__buf_4
XFILLER_0_107_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19500_ clknet_leaf_115_clk _00444_ net1396 vssd1 vssd1 vccd1 vccd1 control.body\[890\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1089 net1092 vssd1 vssd1 vccd1 vccd1 net1089 sky130_fd_sc_hd__buf_4
XFILLER_0_136_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16712_ obsg2.obstacleArray\[88\] obsg2.obstacleArray\[89\] obsg2.obstacleArray\[90\]
+ obsg2.obstacleArray\[91\] net957 net537 vssd1 vssd1 vccd1 vccd1 _02391_ sky130_fd_sc_hd__mux4_1
XFILLER_0_92_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13924_ ag2.body\[68\] net133 _08152_ ag2.body\[60\] vssd1 vssd1 vccd1 vccd1 _00149_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__17215__A2 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17692_ _04045_ net865 net945 _04048_ _03370_ vssd1 vssd1 vccd1 vccd1 _03371_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_137_Left_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12929__B _07472_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19431_ clknet_leaf_108_clk net2376 net1434 vssd1 vssd1 vccd1 vccd1 control.body\[965\]
+ sky130_fd_sc_hd__dfrtp_1
X_16643_ obsg2.obstacleArray\[50\] net444 vssd1 vssd1 vccd1 vccd1 _02322_ sky130_fd_sc_hd__or2_1
XANTENNA__12527__C_N _07460_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13855_ ag2.body\[18\] net117 _08134_ ag2.body\[10\] vssd1 vssd1 vccd1 vccd1 _00098_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_18_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13106__A net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12806_ net342 net328 net309 _07508_ vssd1 vssd1 vccd1 vccd1 _07605_ sky130_fd_sc_hd__and4_1
X_19362_ clknet_leaf_102_clk _00306_ net1428 vssd1 vssd1 vccd1 vccd1 control.body\[1024\]
+ sky130_fd_sc_hd__dfrtp_1
X_16574_ obsg2.obstacleArray\[118\] net445 vssd1 vssd1 vccd1 vccd1 _02253_ sky130_fd_sc_hd__or2_1
XFILLER_0_97_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10998_ ag2.body\[336\] net789 net1090 _04121_ _05966_ vssd1 vssd1 vccd1 vccd1 _05971_
+ sky130_fd_sc_hd__a221o_1
X_13786_ img_gen.updater.commands.count\[13\] _08091_ vssd1 vssd1 vccd1 vccd1 _08094_
+ sky130_fd_sc_hd__nand2_1
XANTENNA__10449__B net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_855 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18313_ _03806_ _03808_ _03794_ vssd1 vssd1 vccd1 vccd1 _03809_ sky130_fd_sc_hd__o21bai_1
X_15525_ ag2.body\[528\] net158 _01610_ ag2.body\[520\] vssd1 vssd1 vccd1 vccd1 _00802_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__17520__B net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19293_ clknet_leaf_98_clk net2187 net1446 vssd1 vssd1 vccd1 vccd1 control.body\[1099\]
+ sky130_fd_sc_hd__dfrtp_1
X_12737_ net334 _07463_ vssd1 vssd1 vccd1 vccd1 _07572_ sky130_fd_sc_hd__or2_2
XANTENNA__12460__B2 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1398 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18244_ _03685_ net37 obsg2.obstacleArray\[119\] vssd1 vssd1 vccd1 vccd1 _03761_
+ sky130_fd_sc_hd__a21oi_1
X_15456_ ag2.body\[595\] net88 _01602_ ag2.body\[587\] vssd1 vssd1 vccd1 vccd1 _00741_
+ sky130_fd_sc_hd__a22o_1
X_12668_ _06671_ _07538_ vssd1 vssd1 vccd1 vccd1 _07539_ sky130_fd_sc_hd__or2_2
XFILLER_0_37_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14407_ net842 net1044 net792 ag2.body\[7\] vssd1 vssd1 vccd1 vccd1 _08568_ sky130_fd_sc_hd__a22o_1
XFILLER_0_5_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18175_ obsg2.obstacleArray\[84\] _03726_ net533 vssd1 vssd1 vccd1 vccd1 _01335_
+ sky130_fd_sc_hd__o21a_1
X_11619_ obsg2.obstacleArray\[53\] net509 vssd1 vssd1 vccd1 vccd1 _06592_ sky130_fd_sc_hd__or2_1
XANTENNA__12212__B2 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15387_ net2596 net70 _01595_ net2188 vssd1 vssd1 vccd1 vccd1 _00679_ sky130_fd_sc_hd__a22o_1
XANTENNA__10465__A net1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12599_ net277 _07499_ _07500_ net1847 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[56\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_114_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17126_ ag2.body\[512\] net886 vssd1 vssd1 vccd1 vccd1 _02805_ sky130_fd_sc_hd__xor2_1
X_14338_ _08494_ _08498_ vssd1 vssd1 vccd1 vccd1 _08499_ sky130_fd_sc_hd__or2_2
XANTENNA__15975__B net56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold506 img_gen.tracker.frame\[393\] vssd1 vssd1 vccd1 vccd1 net2068 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_55_2000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_2011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold517 img_gen.tracker.frame\[37\] vssd1 vssd1 vccd1 vccd1 net2079 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold528 img_gen.tracker.frame\[153\] vssd1 vssd1 vccd1 vccd1 net2090 sky130_fd_sc_hd__dlygate4sd3_1
X_17057_ _02733_ _02734_ _02735_ vssd1 vssd1 vccd1 vccd1 _02736_ sky130_fd_sc_hd__or3b_1
Xhold539 img_gen.tracker.frame\[564\] vssd1 vssd1 vccd1 vccd1 net2101 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09973__B _04420_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14269_ net1027 ag2.body\[13\] vssd1 vssd1 vccd1 vccd1 _08430_ sky130_fd_sc_hd__xor2_1
XANTENNA__12680__A net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16008_ net871 net861 vssd1 vssd1 vccd1 vccd1 _01687_ sky130_fd_sc_hd__nor2_1
XFILLER_0_21_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13495__B _07508_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18100__B1 net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11723__B1 net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18906__CLK clknet_leaf_144_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11296__A net1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1001 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__20196__CLK clknet_leaf_88_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17959_ net518 _03584_ vssd1 vssd1 vccd1 vccd1 _01261_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_68_2405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18079__A net42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18403__A1 _04493_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19629_ clknet_leaf_123_clk net2558 net1407 vssd1 vssd1 vccd1 vccd1 control.body\[763\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_75_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout169_A net171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09988__X _04961_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10359__B net1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09313_ _04319_ _04326_ _04330_ net272 net2228 vssd1 vssd1 vccd1 vccd1 _01440_ sky130_fd_sc_hd__a32o_1
XFILLER_0_91_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout336_A net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_60_clk clknet_4_13__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_60_clk
+ sky130_fd_sc_hd__clkbuf_8
X_09244_ net929 vssd1 vssd1 vccd1 vccd1 _04269_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout1078_A net1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12574__B _07486_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12203__A1 _06986_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09175_ ag2.body\[545\] vssd1 vssd1 vccd1 vccd1 _04200_ sky130_fd_sc_hd__inv_2
XFILLER_0_17_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15940__A2 net196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout503_A _01708_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout124_X net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1245_A net1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20404_ clknet_leaf_31_clk _01291_ net1338 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[40\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_82_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10765__A1 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11962__B1 net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_1_Right_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20335_ clknet_leaf_20_clk _01226_ net1364 vssd1 vssd1 vccd1 vccd1 ag2.apple_cord\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_4_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1033_X net1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16062__A net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput15 net15 vssd1 vssd1 vccd1 vccd1 gpio_out[14] sky130_fd_sc_hd__buf_2
Xoutput26 net26 vssd1 vssd1 vccd1 vccd1 gpio_out[24] sky130_fd_sc_hd__buf_2
XFILLER_0_124_1557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20266_ clknet_leaf_42_clk net1580 net1372 vssd1 vssd1 vccd1 vccd1 control.detect3.Q\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout872_A obsg2.randCord\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout493_X net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10822__B net1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11714__B1 net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17445__A2 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1200_X net1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19831__CLK clknet_leaf_124_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20197_ clknet_leaf_54_clk _01141_ net1455 vssd1 vssd1 vccd1 vccd1 ag2.body\[195\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_60_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08959_ ag2.body\[25\] vssd1 vssd1 vccd1 vccd1 _03984_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout660_X net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout758_X net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14948__C net65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14310__A net1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11970_ img_gen.tracker.frame\[517\] net620 vssd1 vssd1 vccd1 vccd1 _06942_ sky130_fd_sc_hd__or2_1
XFILLER_0_54_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10921_ _05891_ _05892_ _05893_ vssd1 vssd1 vccd1 vccd1 _05894_ sky130_fd_sc_hd__a21oi_1
XANTENNA__11653__B net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16956__A1 ag2.body\[294\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12690__A1 net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16956__B2 ag2.body\[295\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13640_ control.divider.count\[14\] control.divider.count\[13\] _07997_ vssd1 vssd1
+ vccd1 vccd1 _08001_ sky130_fd_sc_hd__and3_1
X_10852_ net1145 control.body\[691\] vssd1 vssd1 vccd1 vccd1 _05825_ sky130_fd_sc_hd__xor2_1
XANTENNA__14967__B1 net51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10269__B net1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout37_X net37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17340__B net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13571_ _07931_ _07944_ _07947_ _07932_ vssd1 vssd1 vccd1 vccd1 net23 sky130_fd_sc_hd__o22a_1
X_10783_ net1147 control.body\[627\] vssd1 vssd1 vccd1 vccd1 _05756_ sky130_fd_sc_hd__xor2_1
XFILLER_0_52_1073 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09989__A3 _04961_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20600__1532 vssd1 vssd1 vccd1 vccd1 _20600__1532/HI net1532 sky130_fd_sc_hd__conb_1
Xclkbuf_leaf_51_clk clknet_4_6__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_51_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_94_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15310_ _04522_ net53 vssd1 vssd1 vccd1 vccd1 _01588_ sky130_fd_sc_hd__nor2_2
XANTENNA__14719__B1 ag2.body\[337\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12522_ net2155 net649 _07458_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[21\]
+ sky130_fd_sc_hd__and3_1
X_16290_ _01967_ _01968_ net417 vssd1 vssd1 vccd1 vccd1 _01969_ sky130_fd_sc_hd__mux2_1
XANTENNA__20069__CLK clknet_leaf_73_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15241_ net2600 net98 _01578_ net2346 vssd1 vssd1 vccd1 vccd1 _00550_ sky130_fd_sc_hd__a22o_1
XFILLER_0_136_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16671__S net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14195__B2 net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12453_ net743 _07372_ vssd1 vssd1 vccd1 vccd1 _07413_ sky130_fd_sc_hd__nand2_1
XFILLER_0_129_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_379 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10205__B1 net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19361__CLK clknet_leaf_102_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11404_ ag2.body\[573\] net1101 vssd1 vssd1 vccd1 vccd1 _06377_ sky130_fd_sc_hd__xor2_1
X_15172_ control.body\[855\] net95 _01570_ control.body\[847\] vssd1 vssd1 vccd1 vccd1
+ _00489_ sky130_fd_sc_hd__a22o_1
X_12384_ _07275_ _07347_ _07348_ vssd1 vssd1 vccd1 vccd1 _07349_ sky130_fd_sc_hd__or3_1
XFILLER_0_65_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11953__B1 net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14123_ net973 ag2.body\[371\] vssd1 vssd1 vccd1 vccd1 _08284_ sky130_fd_sc_hd__xor2_1
X_11335_ net1194 control.body\[657\] vssd1 vssd1 vccd1 vccd1 _06308_ sky130_fd_sc_hd__xor2_1
XFILLER_0_50_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19980_ clknet_leaf_64_clk _00924_ net1474 vssd1 vssd1 vccd1 vccd1 ag2.body\[410\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__17684__A2 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18931_ clknet_leaf_141_clk img_gen.tracker.next_frame\[369\] net1294 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[369\] sky130_fd_sc_hd__dfrtp_1
X_11266_ _06152_ _06179_ _06208_ _06238_ vssd1 vssd1 vccd1 vccd1 _06239_ sky130_fd_sc_hd__and4_1
X_14054_ net1026 ag2.body\[37\] vssd1 vssd1 vccd1 vccd1 _08215_ sky130_fd_sc_hd__xor2_1
XANTENNA__10732__B net1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11705__B1 net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10217_ net750 control.body\[998\] control.body\[999\] net745 _05189_ vssd1 vssd1
+ vccd1 vccd1 _05190_ sky130_fd_sc_hd__o221a_1
X_13005_ net240 _07697_ _07698_ net1897 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[264\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__17436__A2 net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18862_ clknet_leaf_26_clk img_gen.tracker.next_frame\[300\] net1342 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[300\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_94_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11197_ net783 control.body\[872\] control.body\[878\] net748 vssd1 vssd1 vccd1 vccd1
+ _06170_ sky130_fd_sc_hd__a22o_1
XFILLER_0_20_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17813_ _03476_ _03479_ _03480_ _03474_ net925 vssd1 vssd1 vccd1 vccd1 _01220_ sky130_fd_sc_hd__a32o_1
XANTENNA__16644__B1 net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10148_ ag2.body\[58\] net1177 vssd1 vssd1 vccd1 vccd1 _05121_ sky130_fd_sc_hd__or2_1
XANTENNA__17841__C1 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18793_ clknet_leaf_22_clk img_gen.tracker.next_frame\[231\] net1359 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[231\] sky130_fd_sc_hd__dfrtp_1
X_17744_ _02508_ _02510_ _03286_ _03422_ vssd1 vssd1 vccd1 vccd1 _03423_ sky130_fd_sc_hd__o211a_1
X_10079_ _04420_ net638 _05051_ _04587_ vssd1 vssd1 vccd1 vccd1 _05052_ sky130_fd_sc_hd__o31a_1
X_14956_ net2141 net172 _01546_ control.body\[1039\] vssd1 vssd1 vccd1 vccd1 _00297_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__14220__A net1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12130__B1 net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13907_ ag2.body\[53\] net120 _08150_ ag2.body\[45\] vssd1 vssd1 vccd1 vccd1 _00134_
+ sky130_fd_sc_hd__a22o_1
X_17675_ _03345_ _03346_ _03349_ _03353_ vssd1 vssd1 vccd1 vccd1 _03354_ sky130_fd_sc_hd__a211o_1
XFILLER_0_77_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_1547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14887_ control.body\[1097\] net179 _01539_ net2178 vssd1 vssd1 vccd1 vccd1 _00235_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_134_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19414_ clknet_leaf_111_clk _00358_ net1427 vssd1 vssd1 vccd1 vccd1 control.body\[980\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10692__B1 net1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16626_ obsg2.obstacleArray\[35\] net449 net390 vssd1 vssd1 vccd1 vccd1 _02305_ sky130_fd_sc_hd__o21a_1
X_13838_ _06721_ _07372_ _08103_ _08129_ net1070 vssd1 vssd1 vccd1 vccd1 _00086_ sky130_fd_sc_hd__a32o_1
XANTENNA__14958__B1 _01547_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19345_ clknet_leaf_104_clk _00289_ net1431 vssd1 vssd1 vccd1 vccd1 control.body\[1055\]
+ sky130_fd_sc_hd__dfrtp_1
X_16557_ net394 _02235_ _02234_ net359 vssd1 vssd1 vccd1 vccd1 _02236_ sky130_fd_sc_hd__a211o_1
XANTENNA__09968__B net1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13769_ _08082_ vssd1 vssd1 vccd1 vccd1 _08083_ sky130_fd_sc_hd__inv_2
XANTENNA__12675__A net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_42_clk clknet_4_7__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_42_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_45_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15508_ ag2.body\[545\] net155 _01608_ ag2.body\[537\] vssd1 vssd1 vccd1 vccd1 _00787_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11641__C1 net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19276_ clknet_leaf_97_clk net2146 net1450 vssd1 vssd1 vccd1 vccd1 control.body\[1114\]
+ sky130_fd_sc_hd__dfrtp_1
X_16488_ net397 _02161_ _02163_ net366 vssd1 vssd1 vccd1 vccd1 _02167_ sky130_fd_sc_hd__a211o_1
XFILLER_0_45_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18227_ obsg2.obstacleArray\[110\] _03752_ net520 vssd1 vssd1 vccd1 vccd1 _01361_
+ sky130_fd_sc_hd__o21a_1
XANTENNA__15986__A ag2.body\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15439_ ag2.body\[612\] net85 _01600_ ag2.body\[604\] vssd1 vssd1 vccd1 vccd1 _00726_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__15922__A2 net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18362__A _07181_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09984__A net1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13933__B2 ag2.body\[68\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18158_ _03590_ net36 vssd1 vssd1 vccd1 vccd1 _03718_ sky130_fd_sc_hd__nor2_1
XFILLER_0_14_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold303 img_gen.tracker.frame\[288\] vssd1 vssd1 vccd1 vccd1 net1865 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11944__B1 net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17109_ _03977_ net850 net709 ag2.body\[12\] vssd1 vssd1 vccd1 vccd1 _02788_ sky130_fd_sc_hd__a22o_1
Xhold314 img_gen.tracker.frame\[67\] vssd1 vssd1 vccd1 vccd1 net1876 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold325 img_gen.tracker.frame\[109\] vssd1 vssd1 vccd1 vccd1 net1887 sky130_fd_sc_hd__dlygate4sd3_1
X_18089_ _03540_ net299 _03553_ vssd1 vssd1 vccd1 vccd1 _03675_ sky130_fd_sc_hd__or3_1
XANTENNA__19854__CLK clknet_leaf_93_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_492 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold336 img_gen.tracker.frame\[16\] vssd1 vssd1 vccd1 vccd1 net1898 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold347 img_gen.tracker.frame\[387\] vssd1 vssd1 vccd1 vccd1 net1909 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16883__B1 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold358 img_gen.tracker.frame\[150\] vssd1 vssd1 vccd1 vccd1 net1920 sky130_fd_sc_hd__dlygate4sd3_1
X_20120_ clknet_leaf_80_clk _01064_ net1487 vssd1 vssd1 vccd1 vccd1 ag2.body\[278\]
+ sky130_fd_sc_hd__dfrtp_4
X_09931_ net1054 ag2.body\[31\] vssd1 vssd1 vccd1 vccd1 _04904_ sky130_fd_sc_hd__and2b_1
Xhold369 img_gen.tracker.frame\[344\] vssd1 vssd1 vccd1 vccd1 net1931 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_4_3__f_clk clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_3__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_99_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkload23_A clknet_leaf_13_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout805 _03972_ vssd1 vssd1 vccd1 vccd1 net805 sky130_fd_sc_hd__buf_4
XFILLER_0_81_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout816 _03969_ vssd1 vssd1 vccd1 vccd1 net816 sky130_fd_sc_hd__buf_4
X_20051_ clknet_leaf_72_clk _00995_ net1504 vssd1 vssd1 vccd1 vccd1 ag2.body\[337\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA_clkbuf_4_7__f_clk_A clknet_3_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17427__A2 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12560__D net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout827 net831 vssd1 vssd1 vccd1 vccd1 net827 sky130_fd_sc_hd__buf_2
X_09862_ ag2.body\[157\] net1117 vssd1 vssd1 vccd1 vccd1 _04835_ sky130_fd_sc_hd__nand2_1
Xfanout838 net839 vssd1 vssd1 vccd1 vccd1 net838 sky130_fd_sc_hd__buf_2
Xfanout849 net857 vssd1 vssd1 vccd1 vccd1 net849 sky130_fd_sc_hd__buf_2
XANTENNA__16635__B1 net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1003 control.body\[906\] vssd1 vssd1 vccd1 vccd1 net2565 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1014 control.body\[716\] vssd1 vssd1 vccd1 vccd1 net2576 sky130_fd_sc_hd__dlygate4sd3_1
X_09793_ _04753_ _04761_ _04763_ _04765_ vssd1 vssd1 vccd1 vccd1 _04766_ sky130_fd_sc_hd__or4_1
Xhold1025 control.body\[786\] vssd1 vssd1 vccd1 vccd1 net2587 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout286_A net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1036 control.body\[636\] vssd1 vssd1 vccd1 vccd1 net2598 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1047 control.body\[934\] vssd1 vssd1 vccd1 vccd1 net2609 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1058 control.body\[875\] vssd1 vssd1 vccd1 vccd1 net2620 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_119_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1069 control.body\[952\] vssd1 vssd1 vccd1 vccd1 net2631 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1516 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout453_A net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1195_A net1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17060__B1 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14949__B1 _01546_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18256__B net35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09511__X _04484_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17160__B net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09878__B net1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout620_A net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout241_X net241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16057__A net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1362_A net1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout718_A _04265_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_33_clk clknet_4_5__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_33_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_14_1344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout339_X net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14195__A1_N net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11632__C1 net1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_916 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15374__B1 _01594_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09227_ control.body\[1039\] vssd1 vssd1 vccd1 vccd1 _04252_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout1150_X net1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout506_X net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__20361__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09158_ ag2.body\[503\] vssd1 vssd1 vccd1 vccd1 _04183_ sky130_fd_sc_hd__inv_2
XANTENNA__13924__A1 ag2.body\[68\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13924__B2 ag2.body\[60\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09089_ ag2.body\[329\] vssd1 vssd1 vccd1 vccd1 _04114_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_9_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_9_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1415_X net1415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11120_ net1171 control.body\[866\] vssd1 vssd1 vccd1 vccd1 _06093_ sky130_fd_sc_hd__nand2_1
X_20318_ clknet_leaf_44_clk _01214_ net1378 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleFlag
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__16874__B1 net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19589__RESET_B net1386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold870 control.body\[722\] vssd1 vssd1 vccd1 vccd1 net2432 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout875_X net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold881 control.body\[761\] vssd1 vssd1 vccd1 vccd1 net2443 sky130_fd_sc_hd__dlygate4sd3_1
X_11051_ ag2.body\[388\] net763 net749 ag2.body\[390\] _06019_ vssd1 vssd1 vccd1 vccd1
+ _06024_ sky130_fd_sc_hd__o221a_1
XANTENNA__17418__A2 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold892 control.body\[703\] vssd1 vssd1 vccd1 vccd1 net2454 sky130_fd_sc_hd__dlygate4sd3_1
X_20249_ clknet_leaf_70_clk _01193_ net1497 vssd1 vssd1 vccd1 vccd1 ag2.body\[151\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_25_1484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_1375 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16626__B1 net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10002_ net1170 control.body\[730\] vssd1 vssd1 vccd1 vccd1 _04975_ sky130_fd_sc_hd__nand2_1
XFILLER_0_99_1596 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14810_ net834 ag2.body\[377\] ag2.body\[378\] net826 _01479_ vssd1 vssd1 vccd1 vccd1
+ _01481_ sky130_fd_sc_hd__a221o_1
XANTENNA__11664__A net1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14040__A net1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15790_ ag2.body\[300\] net203 _01639_ ag2.body\[292\] vssd1 vssd1 vccd1 vccd1 _01038_
+ sky130_fd_sc_hd__a22o_1
X_14741_ net985 _04115_ ag2.body\[332\] net815 vssd1 vssd1 vccd1 vccd1 _08902_ sky130_fd_sc_hd__a22o_1
XFILLER_0_87_917 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11953_ img_gen.tracker.frame\[109\] net619 net547 img_gen.tracker.frame\[115\] _06924_
+ vssd1 vssd1 vccd1 vccd1 _06925_ sky130_fd_sc_hd__o221a_1
XANTENNA__13860__B1 _08134_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14778__A1_N net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20076__RESET_B net1492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17051__B1 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17460_ _03135_ _03136_ _03137_ _03138_ vssd1 vssd1 vccd1 vccd1 _03139_ sky130_fd_sc_hd__or4_1
X_10904_ net1072 control.body\[678\] vssd1 vssd1 vccd1 vccd1 _05877_ sky130_fd_sc_hd__xor2_1
X_14672_ net826 ag2.body\[386\] ag2.body\[385\] net834 vssd1 vssd1 vccd1 vccd1 _08833_
+ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__18601__CLK clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_3973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08973__A ag2.body\[63\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19727__CLK clknet_leaf_132_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11884_ _06853_ _06855_ net474 vssd1 vssd1 vccd1 vccd1 _06856_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_120_3984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16411_ net401 _02089_ _02088_ net364 vssd1 vssd1 vccd1 vccd1 _02090_ sky130_fd_sc_hd__a211o_1
XFILLER_0_19_1299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13623_ control.divider.count\[7\] control.divider.count\[8\] _07987_ vssd1 vssd1
+ vccd1 vccd1 _07990_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_120_3995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10835_ ag2.body\[304\] net1236 vssd1 vssd1 vccd1 vccd1 _05808_ sky130_fd_sc_hd__nand2_1
X_17391_ _03058_ _03061_ _03064_ _03069_ vssd1 vssd1 vccd1 vccd1 _03070_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_101_3394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_24_clk clknet_4_6__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_24_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_95_994 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19130_ clknet_leaf_141_clk img_gen.tracker.next_frame\[568\] net1296 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[568\] sky130_fd_sc_hd__dfrtp_1
X_16342_ obsg2.obstacleArray\[94\] obsg2.obstacleArray\[95\] net408 vssd1 vssd1 vccd1
+ vccd1 _02021_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13554_ ssdec1.in\[3\] _07931_ vssd1 vssd1 vccd1 vccd1 _07936_ sky130_fd_sc_hd__nand2_1
XFILLER_0_125_702 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10766_ _05727_ _05732_ _05734_ _05738_ vssd1 vssd1 vccd1 vccd1 _05739_ sky130_fd_sc_hd__or4_2
XFILLER_0_13_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10727__B net1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14168__A1 net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12505_ net606 _06638_ net439 net565 vssd1 vssd1 vccd1 vccd1 _07448_ sky130_fd_sc_hd__or4_1
X_19061_ clknet_leaf_9_clk img_gen.tracker.next_frame\[499\] net1271 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[499\] sky130_fd_sc_hd__dfrtp_1
X_16273_ obsg2.obstacleArray\[27\] net413 _01951_ net416 vssd1 vssd1 vccd1 vccd1 _01952_
+ sky130_fd_sc_hd__o211a_1
XANTENNA__14168__B2 net1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15365__B1 _01593_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15904__A2 net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10697_ _04470_ net634 vssd1 vssd1 vccd1 vccd1 _05670_ sky130_fd_sc_hd__nor2_2
X_13485_ net336 net332 net308 _07501_ vssd1 vssd1 vccd1 vccd1 _07906_ sky130_fd_sc_hd__or4_1
XFILLER_0_120_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18012_ obsg2.obstacleArray\[24\] _03623_ net532 vssd1 vssd1 vccd1 vccd1 _01275_
+ sky130_fd_sc_hd__o21a_1
XANTENNA__13915__A1 ag2.body\[60\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15224_ net2566 net92 _01576_ control.body\[797\] vssd1 vssd1 vccd1 vccd1 _00535_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_106_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12436_ img_gen.updater.commands.rR1.rainbowRNG\[6\] net248 _07377_ vssd1 vssd1 vccd1
+ vccd1 _07397_ sky130_fd_sc_hd__a21o_1
XFILLER_0_129_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15117__B1 _01554_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_114_3788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15155_ _06207_ net53 vssd1 vssd1 vccd1 vccd1 _01569_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_114_3799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16314__C1 net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12367_ _07172_ _07173_ _07302_ vssd1 vssd1 vccd1 vccd1 _07333_ sky130_fd_sc_hd__and3_1
XANTENNA__14215__A net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12661__C net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14106_ net840 ag2.body\[584\] _04213_ net987 _08266_ vssd1 vssd1 vccd1 vccd1 _08267_
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_65_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11318_ ag2.body\[559\] net1052 vssd1 vssd1 vccd1 vccd1 _06291_ sky130_fd_sc_hd__xor2_1
XFILLER_0_61_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19963_ clknet_leaf_62_clk _00907_ net1469 vssd1 vssd1 vccd1 vccd1 ag2.body\[425\]
+ sky130_fd_sc_hd__dfrtp_4
X_15086_ net2250 net147 _01562_ net2321 vssd1 vssd1 vccd1 vccd1 _00411_ sky130_fd_sc_hd__a22o_1
X_12298_ _07210_ _07263_ _07264_ vssd1 vssd1 vccd1 vccd1 _07265_ sky130_fd_sc_hd__and3b_1
XANTENNA__13679__B1 net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19259__RESET_B net1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14037_ net837 ag2.body\[497\] _04181_ net1039 vssd1 vssd1 vccd1 vccd1 _08198_ sky130_fd_sc_hd__o22a_1
X_11249_ ag2.body\[196\] net1138 vssd1 vssd1 vccd1 vccd1 _06222_ sky130_fd_sc_hd__nand2_1
X_18914_ clknet_leaf_142_clk img_gen.tracker.next_frame\[352\] net1253 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[352\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_129_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19894_ clknet_leaf_86_clk _00838_ net1462 vssd1 vssd1 vccd1 vccd1 ag2.body\[500\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_78_1603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18845_ clknet_leaf_4_clk img_gen.tracker.next_frame\[283\] net1277 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[283\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__16712__S0 net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17290__B1 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18776_ clknet_leaf_16_clk img_gen.tracker.next_frame\[214\] net1315 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[214\] sky130_fd_sc_hd__dfrtp_1
X_15988_ _01667_ _01671_ vssd1 vssd1 vccd1 vccd1 _01672_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_89_210 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12103__B1 net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17727_ net497 _03405_ _03404_ _01709_ vssd1 vssd1 vccd1 vccd1 _03406_ sky130_fd_sc_hd__a211o_1
X_14939_ net895 _04792_ net65 vssd1 vssd1 vccd1 vccd1 _01545_ sky130_fd_sc_hd__and3_2
Xclkbuf_4_11__f_clk clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_11__leaf_clk
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__16576__S net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14885__A net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17658_ ag2.body\[106\] net866 vssd1 vssd1 vccd1 vccd1 _03337_ sky130_fd_sc_hd__nand2_1
XANTENNA__09979__A net1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16609_ obsg2.obstacleArray\[94\] obsg2.obstacleArray\[95\] net445 vssd1 vssd1 vccd1
+ vccd1 _02288_ sky130_fd_sc_hd__mux2_1
XANTENNA__09698__B net1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17589_ ag2.body\[58\] net725 net705 ag2.body\[61\] vssd1 vssd1 vccd1 vccd1 _03268_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_4_1629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18823__RESET_B net1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_15_clk clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_15_clk
+ sky130_fd_sc_hd__clkbuf_8
X_19328_ clknet_leaf_104_clk net2185 net1431 vssd1 vssd1 vccd1 vccd1 control.body\[1070\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_324 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14159__A1 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19259_ clknet_leaf_74_clk _00203_ net1495 vssd1 vssd1 vccd1 vccd1 ag2.body\[122\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__15356__B1 _01592_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14159__B2 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16553__C1 net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17896__A2 _03531_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09012_ ag2.body\[138\] vssd1 vssd1 vccd1 vccd1 _04037_ sky130_fd_sc_hd__inv_2
XFILLER_0_116_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold100 img_gen.tracker.frame\[483\] vssd1 vssd1 vccd1 vccd1 net1662 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_130_4280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11749__A net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16305__C1 net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout201_A net204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold111 img_gen.tracker.frame\[523\] vssd1 vssd1 vccd1 vccd1 net1673 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_130_4291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14125__A net1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold122 img_gen.tracker.frame\[133\] vssd1 vssd1 vccd1 vccd1 net1684 sky130_fd_sc_hd__dlygate4sd3_1
Xhold133 img_gen.tracker.frame\[145\] vssd1 vssd1 vccd1 vccd1 net1695 sky130_fd_sc_hd__dlygate4sd3_1
Xhold144 img_gen.tracker.frame\[233\] vssd1 vssd1 vccd1 vccd1 net1706 sky130_fd_sc_hd__dlygate4sd3_1
Xhold155 img_gen.tracker.frame\[422\] vssd1 vssd1 vccd1 vccd1 net1717 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__16320__A2 net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold166 img_gen.tracker.frame\[217\] vssd1 vssd1 vccd1 vccd1 net1728 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold177 img_gen.tracker.frame\[302\] vssd1 vssd1 vccd1 vccd1 net1739 sky130_fd_sc_hd__dlygate4sd3_1
X_20103_ clknet_leaf_78_clk _01047_ net1489 vssd1 vssd1 vccd1 vccd1 ag2.body\[293\]
+ sky130_fd_sc_hd__dfrtp_4
Xhold188 img_gen.tracker.frame\[385\] vssd1 vssd1 vccd1 vccd1 net1750 sky130_fd_sc_hd__dlygate4sd3_1
X_09914_ ag2.body\[134\] net1090 vssd1 vssd1 vccd1 vccd1 _04887_ sky130_fd_sc_hd__xor2_1
XANTENNA__13964__A _05347_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout602 _06476_ vssd1 vssd1 vccd1 vccd1 net602 sky130_fd_sc_hd__clkbuf_4
Xhold199 img_gen.tracker.frame\[500\] vssd1 vssd1 vccd1 vccd1 net1761 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_1624 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout613 net615 vssd1 vssd1 vccd1 vccd1 net613 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_61_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1110_A net1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout624 net625 vssd1 vssd1 vccd1 vccd1 net624 sky130_fd_sc_hd__buf_2
XANTENNA_fanout1208_A net1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20034_ clknet_leaf_67_clk _00978_ net1494 vssd1 vssd1 vccd1 vccd1 ag2.body\[352\]
+ sky130_fd_sc_hd__dfrtp_4
Xfanout646 net654 vssd1 vssd1 vccd1 vccd1 net646 sky130_fd_sc_hd__buf_2
XFILLER_0_42_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input6_A gpio_in[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout657 net658 vssd1 vssd1 vccd1 vccd1 net657 sky130_fd_sc_hd__dlymetal6s2s_1
X_09845_ _04784_ _04786_ _04795_ _04817_ vssd1 vssd1 vccd1 vccd1 _04818_ sky130_fd_sc_hd__o31a_1
XANTENNA_fanout191_X net191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout668 net669 vssd1 vssd1 vccd1 vccd1 net668 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout570_A net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12893__A1 net246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout679 net681 vssd1 vssd1 vccd1 vccd1 net679 sky130_fd_sc_hd__clkbuf_2
XANTENNA__16084__A1 net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20516__RESET_B net1403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout668_A net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout289_X net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18624__CLK clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09776_ _04072_ net1159 net755 ag2.body\[237\] _04741_ vssd1 vssd1 vccd1 vccd1 _04749_
+ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_124_4095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16486__S net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout835_A net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout456_X net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1198_X net1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09889__A _04446_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17584__A1 ag2.body\[56\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14398__A1 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14398__B2 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18774__CLK clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout623_X net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10671__A3 _05632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11605__C1 _06485_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10620_ ag2.body\[52\] net1121 vssd1 vssd1 vccd1 vccd1 _05593_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_137_4489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13070__A1 net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_1088 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10547__B net1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_201 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10551_ ag2.body\[224\] net1231 vssd1 vssd1 vccd1 vccd1 _05524_ sky130_fd_sc_hd__xor2_1
XFILLER_0_52_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13270_ net236 _07821_ _07822_ net1745 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[405\]
+ sky130_fd_sc_hd__a22o_1
X_10482_ ag2.body\[584\] net1219 vssd1 vssd1 vccd1 vccd1 _05455_ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout992_X net992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12762__B _07584_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12221_ img_gen.updater.commands.count\[2\] _07189_ img_gen.updater.commands.count\[3\]
+ img_gen.updater.commands.count\[4\] vssd1 vssd1 vccd1 vccd1 _07191_ sky130_fd_sc_hd__a211o_1
XFILLER_0_126_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14035__A net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12481__C net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12152_ img_gen.tracker.frame\[435\] net597 net579 img_gen.tracker.frame\[441\] _07123_
+ vssd1 vssd1 vccd1 vccd1 _07124_ sky130_fd_sc_hd__o221a_1
XFILLER_0_62_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17457__A2_N net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11103_ ag2.body\[429\] net754 net1081 _04153_ _06070_ vssd1 vssd1 vccd1 vccd1 _06076_
+ sky130_fd_sc_hd__o221a_1
XANTENNA__13874__A _04903_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17346__A net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14322__B2 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16960_ ag2.body\[293\] net955 vssd1 vssd1 vccd1 vccd1 _02639_ sky130_fd_sc_hd__nand2_1
X_12083_ net576 _07054_ vssd1 vssd1 vccd1 vccd1 _07055_ sky130_fd_sc_hd__or2_1
XFILLER_0_124_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15911_ ag2.body\[184\] net131 _01652_ ag2.body\[176\] vssd1 vssd1 vccd1 vccd1 _01146_
+ sky130_fd_sc_hd__a22o_1
X_11034_ net786 control.body\[1040\] control.body\[1045\] net755 _06006_ vssd1 vssd1
+ vccd1 vccd1 _06007_ sky130_fd_sc_hd__o221a_1
XFILLER_0_60_1183 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17065__B net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16891_ ag2.body\[212\] net964 vssd1 vssd1 vccd1 vccd1 _02570_ sky130_fd_sc_hd__or2_1
XFILLER_0_102_1482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18630_ clknet_leaf_0_clk img_gen.tracker.next_frame\[68\] net1242 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[68\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__11394__A net1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15842_ ag2.body\[251\] net181 _01644_ ag2.body\[243\] vssd1 vssd1 vccd1 vccd1 _01085_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_107_3581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18561_ clknet_leaf_132_clk _00087_ net1304 vssd1 vssd1 vccd1 vccd1 ag2.x\[3\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_107_3592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15773_ ag2.body\[317\] net203 _01637_ ag2.body\[309\] vssd1 vssd1 vccd1 vccd1 _01023_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12636__A1 net241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12985_ net337 net333 _07508_ vssd1 vssd1 vccd1 vccd1 _07688_ sky130_fd_sc_hd__and3_1
XFILLER_0_73_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_3456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17512_ ag2.body\[589\] net946 vssd1 vssd1 vccd1 vccd1 _03191_ sky130_fd_sc_hd__xor2_1
X_14724_ net985 ag2.body\[114\] vssd1 vssd1 vccd1 vccd1 _08885_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_103_3467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11936_ img_gen.tracker.frame\[181\] net621 net603 img_gen.tracker.frame\[184\] _06907_
+ vssd1 vssd1 vccd1 vccd1 _06908_ sky130_fd_sc_hd__o221a_1
X_18492_ net1516 net1510 vssd1 vssd1 vccd1 vccd1 _00023_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_103_3478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17443_ _04134_ net862 net705 ag2.body\[381\] vssd1 vssd1 vccd1 vccd1 _03122_ sky130_fd_sc_hd__a22o_1
X_14655_ net1013 ag2.body\[151\] vssd1 vssd1 vccd1 vccd1 _08816_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10297__X _05270_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14389__B2 net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11867_ img_gen.tracker.frame\[265\] net622 vssd1 vssd1 vccd1 vccd1 _06839_ sky130_fd_sc_hd__or2_1
XFILLER_0_39_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13606_ control.divider.count\[0\] net220 vssd1 vssd1 vccd1 vccd1 control.divider.next_count\[0\]
+ sky130_fd_sc_hd__and2b_1
X_17374_ _03007_ _03047_ vssd1 vssd1 vccd1 vccd1 _03053_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_27_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10818_ _05788_ _05789_ _05790_ vssd1 vssd1 vccd1 vccd1 _05791_ sky130_fd_sc_hd__a21o_1
XANTENNA__13061__A1 net246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14586_ net977 _04013_ ag2.body\[86\] net802 _08746_ vssd1 vssd1 vccd1 vccd1 _08747_
+ sky130_fd_sc_hd__a221o_1
XANTENNA__10457__B net1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11798_ net472 _06761_ _06764_ _06769_ net466 vssd1 vssd1 vccd1 vccd1 _06770_ sky130_fd_sc_hd__o221a_1
X_19113_ clknet_leaf_0_clk img_gen.tracker.next_frame\[551\] net1245 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[551\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_28_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11072__B1 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16325_ net369 _02003_ _02000_ net368 vssd1 vssd1 vccd1 vccd1 _02004_ sky130_fd_sc_hd__o211a_1
XANTENNA__15338__B1 _01590_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13537_ img_gen.tracker.frame\[569\] net659 _07925_ vssd1 vssd1 vccd1 vccd1 _07926_
+ sky130_fd_sc_hd__and3_1
X_10749_ _05718_ _05719_ _05720_ _05721_ vssd1 vssd1 vccd1 vccd1 _05722_ sky130_fd_sc_hd__or4_1
XFILLER_0_40_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12953__A net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15889__A1 ag2.body\[213\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19044_ clknet_leaf_7_clk img_gen.tracker.next_frame\[482\] net1268 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[482\] sky130_fd_sc_hd__dfrtp_1
X_16256_ obsg2.obstacleArray\[56\] net407 vssd1 vssd1 vccd1 vccd1 _01935_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_11_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_1561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13468_ net256 _07898_ _07899_ net1899 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[526\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_125_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1640 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15207_ control.body\[822\] net92 _01574_ net2402 vssd1 vssd1 vccd1 vccd1 _00520_
+ sky130_fd_sc_hd__a22o_1
X_12419_ net767 _06477_ vssd1 vssd1 vccd1 vccd1 _07381_ sky130_fd_sc_hd__nand2_1
X_16187_ obsg2.obstacleArray\[50\] obsg2.obstacleArray\[51\] net422 vssd1 vssd1 vccd1
+ vccd1 _01866_ sky130_fd_sc_hd__mux2_1
XANTENNA__10473__A net1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13399_ net259 net312 _07551_ _07872_ net1688 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[484\]
+ sky130_fd_sc_hd__a32o_1
XANTENNA__16838__B1 net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15138_ control.body\[872\] net105 _01567_ net2411 vssd1 vssd1 vccd1 vccd1 _00458_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_65_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10192__B net1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19946_ clknet_leaf_45_clk _00890_ net1382 vssd1 vssd1 vccd1 vccd1 ag2.body\[440\]
+ sky130_fd_sc_hd__dfrtp_2
X_15069_ control.body\[938\] net149 _01560_ net2425 vssd1 vssd1 vccd1 vccd1 _00396_
+ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_4_clk clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_4_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_71_2478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_2489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_1411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19877_ clknet_leaf_91_clk _00821_ net1415 vssd1 vssd1 vccd1 vccd1 ag2.body\[515\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__10920__B net1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17263__B1 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09630_ net890 net900 net904 net896 vssd1 vssd1 vccd1 vccd1 _04603_ sky130_fd_sc_hd__or4bb_4
XFILLER_0_120_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18828_ clknet_leaf_4_clk img_gen.tracker.next_frame\[266\] net1262 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[266\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_88_2997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09561_ _04523_ _04524_ _04529_ _04533_ vssd1 vssd1 vccd1 vccd1 _04534_ sky130_fd_sc_hd__or4_2
XANTENNA__13008__B _07523_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18759_ clknet_leaf_15_clk img_gen.tracker.next_frame\[197\] net1313 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[197\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_136_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18087__A net44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09492_ ag2.body\[375\] net1056 vssd1 vssd1 vccd1 vccd1 _04465_ sky130_fd_sc_hd__xor2_1
XANTENNA__14608__A1_N net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12847__B _07624_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16319__B net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout151_A net154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16038__C net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13052__A1 net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_882 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20583_ clknet_leaf_107_clk _01440_ _00047_ vssd1 vssd1 vccd1 vccd1 sound_gen.osc1.count\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_132_4342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1060_A net1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout416_A net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_132_4353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1158_A net1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_132_4364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_41_1570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_552 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19422__CLK clknet_leaf_111_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout204_X net204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16829__B1 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout785_A net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14304__A1 net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09891__B net1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14304__B2 net1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10670__X _05643_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1113_X net1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11118__B2 _06090_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout410 net412 vssd1 vssd1 vccd1 vccd1 net410 sky130_fd_sc_hd__buf_2
XANTENNA__12315__B1 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1408 net1409 vssd1 vssd1 vccd1 vccd1 net1408 sky130_fd_sc_hd__clkbuf_2
Xfanout421 net423 vssd1 vssd1 vccd1 vccd1 net421 sky130_fd_sc_hd__clkbuf_4
Xfanout1419 net1435 vssd1 vssd1 vccd1 vccd1 net1419 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_54_1964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout432 _01705_ vssd1 vssd1 vccd1 vccd1 net432 sky130_fd_sc_hd__buf_2
XFILLER_0_100_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_54_1975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout443 _02214_ vssd1 vssd1 vccd1 vccd1 net443 sky130_fd_sc_hd__clkbuf_4
XANTENNA_input9_X net9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout454 net459 vssd1 vssd1 vccd1 vccd1 net454 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_126_4168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout952_A net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout573_X net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout465 _07180_ vssd1 vssd1 vccd1 vccd1 net465 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_35_1385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20017_ clknet_leaf_56_clk _00961_ net1467 vssd1 vssd1 vccd1 vccd1 ag2.body\[383\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_35_1396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17254__B1 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_122_Right_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout487 net489 vssd1 vssd1 vccd1 vccd1 net487 sky130_fd_sc_hd__clkbuf_4
X_09828_ net1133 control.body\[924\] vssd1 vssd1 vccd1 vccd1 _04801_ sky130_fd_sc_hd__or2_1
XFILLER_0_57_1506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout498 net499 vssd1 vssd1 vccd1 vccd1 net498 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout64_A _08131_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10341__A2 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout740_X net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09759_ ag2.body\[214\] net1089 vssd1 vssd1 vccd1 vccd1 _04732_ sky130_fd_sc_hd__or2_1
XANTENNA__12618__A1 net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17613__B net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_100_Left_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1482_X net1482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17006__B1 net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout838_X net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13291__A1 net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12770_ net235 _07588_ _07589_ net1932 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[138\]
+ sky130_fd_sc_hd__a22o_1
X_11721_ img_gen.tracker.frame\[227\] net590 net551 img_gen.tracker.frame\[224\] _06692_
+ vssd1 vssd1 vccd1 vccd1 _06693_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_48_1779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11841__A2 net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14440_ net840 ag2.body\[16\] _03983_ net1035 _08595_ vssd1 vssd1 vccd1 vccd1 _08601_
+ sky130_fd_sc_hd__o221a_1
X_11652_ net1118 net1070 vssd1 vssd1 vccd1 vccd1 _06625_ sky130_fd_sc_hd__nor2_1
XFILLER_0_132_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout50 _01548_ vssd1 vssd1 vccd1 vccd1 net50 sky130_fd_sc_hd__buf_2
Xfanout61 net62 vssd1 vssd1 vccd1 vccd1 net61 sky130_fd_sc_hd__buf_6
Xfanout72 net79 vssd1 vssd1 vccd1 vccd1 net72 sky130_fd_sc_hd__dlymetal6s2s_1
X_10603_ net1161 control.body\[987\] vssd1 vssd1 vccd1 vccd1 _05576_ sky130_fd_sc_hd__nand2_1
XANTENNA__13869__A net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14371_ net1037 ag2.body\[420\] vssd1 vssd1 vccd1 vccd1 _08532_ sky130_fd_sc_hd__xor2_1
Xfanout83 net91 vssd1 vssd1 vccd1 vccd1 net83 sky130_fd_sc_hd__buf_2
XFILLER_0_135_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16517__C1 net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout94 net100 vssd1 vssd1 vccd1 vccd1 net94 sky130_fd_sc_hd__buf_2
X_11583_ net1192 net1144 vssd1 vssd1 vccd1 vccd1 _06556_ sky130_fd_sc_hd__nand2_1
XANTENNA__12773__A net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_852 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16110_ net374 _01786_ _01788_ net348 vssd1 vssd1 vccd1 vccd1 _01789_ sky130_fd_sc_hd__a211o_1
X_13322_ _06823_ _07498_ vssd1 vssd1 vccd1 vccd1 _07842_ sky130_fd_sc_hd__nor2_1
XFILLER_0_52_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17090_ ag2.body\[303\] net933 vssd1 vssd1 vccd1 vccd1 _02769_ sky130_fd_sc_hd__xnor2_1
X_10534_ net1158 control.body\[915\] vssd1 vssd1 vccd1 vccd1 _05507_ sky130_fd_sc_hd__xor2_1
XFILLER_0_122_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_111_3703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_3179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_3714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16041_ net433 _01719_ vssd1 vssd1 vccd1 vccd1 _01720_ sky130_fd_sc_hd__nor2_2
XANTENNA__11389__A net1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10465_ net1109 control.body\[1013\] vssd1 vssd1 vccd1 vccd1 _05438_ sky130_fd_sc_hd__or2_1
X_13253_ _07443_ net303 vssd1 vssd1 vccd1 vccd1 _07815_ sky130_fd_sc_hd__nor2_1
X_12204_ _06825_ _07175_ vssd1 vssd1 vccd1 vccd1 _07176_ sky130_fd_sc_hd__nor2_1
XFILLER_0_62_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19915__CLK clknet_leaf_52_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13184_ net336 net277 net327 _07515_ _07782_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[359\]
+ sky130_fd_sc_hd__a41o_1
X_10396_ net1110 control.body\[1061\] vssd1 vssd1 vccd1 vccd1 _05369_ sky130_fd_sc_hd__nand2_1
X_19800_ clknet_leaf_127_clk _00744_ net1330 vssd1 vssd1 vccd1 vccd1 ag2.body\[598\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__17493__B1 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12135_ img_gen.tracker.frame\[483\] net602 net586 img_gen.tracker.frame\[489\] _07106_
+ vssd1 vssd1 vccd1 vccd1 _07107_ sky130_fd_sc_hd__o221a_1
X_17992_ net38 _03608_ vssd1 vssd1 vccd1 vccd1 _03609_ sky130_fd_sc_hd__and2_1
XFILLER_0_100_1419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19731_ clknet_leaf_129_clk _00675_ net1327 vssd1 vssd1 vccd1 vccd1 control.body\[657\]
+ sky130_fd_sc_hd__dfrtp_1
X_16943_ _02617_ _02619_ _02621_ vssd1 vssd1 vccd1 vccd1 _02622_ sky130_fd_sc_hd__or3_4
X_12066_ _06690_ _07036_ _07037_ net435 vssd1 vssd1 vccd1 vccd1 _07038_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_109_3643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10740__B net1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_3654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17245__B1 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11017_ _05986_ _05987_ _05988_ _05989_ vssd1 vssd1 vccd1 vccd1 _05990_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_105_3518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1032 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16874_ ag2.body\[466\] net723 net929 _04167_ _02552_ vssd1 vssd1 vccd1 vccd1 _02553_
+ sky130_fd_sc_hd__a221o_1
X_19662_ clknet_leaf_134_clk _00606_ net1391 vssd1 vssd1 vccd1 vccd1 control.body\[732\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_105_3529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20020__RESET_B net1464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15825_ ag2.body\[267\] net201 _01643_ ag2.body\[259\] vssd1 vssd1 vccd1 vccd1 _01069_
+ sky130_fd_sc_hd__a22o_1
X_18613_ clknet_leaf_145_clk img_gen.tracker.next_frame\[51\] net1241 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[51\] sky130_fd_sc_hd__dfrtp_1
X_19593_ clknet_leaf_117_clk _00537_ net1386 vssd1 vssd1 vccd1 vccd1 control.body\[807\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_95_1087 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10883__A3 _04471_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15756_ ag2.body\[334\] net216 _01635_ ag2.body\[326\] vssd1 vssd1 vccd1 vccd1 _01008_
+ sky130_fd_sc_hd__a22o_1
X_18544_ clknet_leaf_135_clk _00070_ net1298 vssd1 vssd1 vccd1 vccd1 img_gen.updater.commands.count\[13\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__20587__D ag2.goodColl vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_83_2850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12968_ net278 _07678_ _07679_ net1938 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[245\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__13282__A1 net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12085__A2 net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_83_2861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12667__B _06639_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_0_clk_A clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14707_ net975 ag2.body\[235\] vssd1 vssd1 vccd1 vccd1 _08868_ sky130_fd_sc_hd__xor2_1
X_11919_ net1225 net1199 img_gen.tracker.frame\[325\] vssd1 vssd1 vccd1 vccd1 _06891_
+ sky130_fd_sc_hd__or3_1
XFILLER_0_73_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18475_ net1514 net1508 vssd1 vssd1 vccd1 vccd1 _00006_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_64_2260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15687_ ag2.body\[385\] net136 _01616_ ag2.body\[377\] vssd1 vssd1 vccd1 vccd1 _00947_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11832__A2 net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10468__A net1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_2271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12899_ img_gen.tracker.frame\[208\] net661 vssd1 vssd1 vccd1 vccd1 _07649_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_64_2282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17426_ ag2.body\[114\] net728 net702 ag2.body\[118\] vssd1 vssd1 vccd1 vccd1 _03105_
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_136_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14638_ net840 ag2.body\[576\] ag2.body\[577\] net832 _08798_ vssd1 vssd1 vccd1 vccd1
+ _08799_ sky130_fd_sc_hd__o221ai_1
XFILLER_0_111_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_2146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16771__A2 net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_2157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18354__B _07181_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_2168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14594__A1_N net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17357_ _03013_ _03015_ _03021_ _03033_ vssd1 vssd1 vccd1 vccd1 _03036_ sky130_fd_sc_hd__or4_1
XFILLER_0_43_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14782__A1 net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14569_ net977 _04127_ _04128_ net1013 _08727_ vssd1 vssd1 vccd1 vccd1 _08730_ sky130_fd_sc_hd__a221o_1
XANTENNA__12683__A net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14782__B2 net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16308_ obsg2.obstacleArray\[104\] net405 vssd1 vssd1 vccd1 vccd1 _01987_ sky130_fd_sc_hd__or2_1
XFILLER_0_12_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_351 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17288_ ag2.body\[304\] net887 vssd1 vssd1 vccd1 vccd1 _02967_ sky130_fd_sc_hd__xor2_1
XANTENNA__10915__B net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload20 clknet_leaf_10_clk vssd1 vssd1 vccd1 vccd1 clkload20/Y sky130_fd_sc_hd__inv_6
XFILLER_0_125_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11299__A net1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19027_ clknet_leaf_1_clk img_gen.tracker.next_frame\[465\] net1246 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[465\] sky130_fd_sc_hd__dfrtp_1
X_16239_ _01892_ _01917_ vssd1 vssd1 vccd1 vccd1 _01918_ sky130_fd_sc_hd__or2_4
XTAP_TAPCELL_ROW_77_2665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload31 clknet_leaf_136_clk vssd1 vssd1 vccd1 vccd1 clkload31/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_63_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14534__A1 net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_2676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload42 clknet_leaf_129_clk vssd1 vssd1 vccd1 vccd1 clkload42/Y sky130_fd_sc_hd__inv_6
XFILLER_0_42_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14534__B2 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload53 clknet_leaf_35_clk vssd1 vssd1 vccd1 vccd1 clkload53/Y sky130_fd_sc_hd__clkinv_8
XFILLER_0_109_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload64 clknet_leaf_53_clk vssd1 vssd1 vccd1 vccd1 clkload64/Y sky130_fd_sc_hd__inv_4
XFILLER_0_3_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_58_2086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload75 clknet_leaf_116_clk vssd1 vssd1 vccd1 vccd1 clkload75/Y sky130_fd_sc_hd__bufinv_16
XFILLER_0_23_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload86 clknet_leaf_104_clk vssd1 vssd1 vccd1 vccd1 clkload86/Y sky130_fd_sc_hd__clkinv_8
XTAP_TAPCELL_ROW_58_2097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload97 clknet_leaf_95_clk vssd1 vssd1 vccd1 vccd1 clkload97/Y sky130_fd_sc_hd__inv_6
XFILLER_0_11_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14403__A net1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08992_ ag2.body\[89\] vssd1 vssd1 vccd1 vccd1 _04017_ sky130_fd_sc_hd__inv_2
XANTENNA__14298__B1 net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14837__A2 _08479_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19929_ clknet_leaf_51_clk _00873_ net1369 vssd1 vssd1 vccd1 vccd1 ag2.body\[471\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__15218__B net53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10650__B net1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17236__B1 net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout199_A net200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_3_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09713__A1 net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_121_4010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09613_ net891 net909 net913 vssd1 vssd1 vccd1 vccd1 _04586_ sky130_fd_sc_hd__or3_4
XFILLER_0_78_500 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout366_A _02067_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09544_ net761 control.body\[1028\] net895 vssd1 vssd1 vccd1 vccd1 _04517_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_78_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12076__A2 net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_4540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09475_ ag2.body\[469\] net1102 vssd1 vssd1 vccd1 vccd1 _04448_ sky130_fd_sc_hd__xor2_1
XFILLER_0_38_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11823__A2 net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_4551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout533_A net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout154_X net154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_4562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1275_A net1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_134_4404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_134_4415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13025__A1 net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_43_1621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_1632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20635_ net1552 vssd1 vssd1 vccd1 vccd1 gpio_out[30] sky130_fd_sc_hd__buf_2
XANTENNA_fanout700_A net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12593__A net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1442_A net1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout419_X net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload3 clknet_4_7__leaf_clk vssd1 vssd1 vccd1 vccd1 clkload3/X sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout1063_X net1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_24_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20566_ clknet_leaf_43_clk _01425_ net1379 vssd1 vssd1 vccd1 vccd1 obsg2.randCord\[2\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_11_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20497_ clknet_leaf_21_clk _01384_ net1361 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[133\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA_fanout1230_X net1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10250_ net890 _04979_ _04492_ vssd1 vssd1 vccd1 vccd1 _05223_ sky130_fd_sc_hd__o21a_1
XFILLER_0_132_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout690_X net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_4219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout788_X net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10181_ ag2.body\[423\] net1057 vssd1 vssd1 vccd1 vccd1 _05154_ sky130_fd_sc_hd__or2_1
XFILLER_0_121_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_37_1447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14313__A net996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1205 net1214 vssd1 vssd1 vccd1 vccd1 net1205 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10562__A2 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1628 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11656__B net1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1216 net1221 vssd1 vssd1 vccd1 vccd1 net1216 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12839__A1 net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1227 net1228 vssd1 vssd1 vccd1 vccd1 net1227 sky130_fd_sc_hd__clkbuf_4
XANTENNA__15128__B net58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout955_X net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1238 ag2.y\[0\] vssd1 vssd1 vccd1 vccd1 net1238 sky130_fd_sc_hd__clkbuf_8
Xfanout240 net242 vssd1 vssd1 vccd1 vccd1 net240 sky130_fd_sc_hd__clkbuf_4
Xfanout1249 net1250 vssd1 vssd1 vccd1 vccd1 net1249 sky130_fd_sc_hd__clkbuf_4
Xfanout251 net260 vssd1 vssd1 vccd1 vccd1 net251 sky130_fd_sc_hd__clkbuf_2
XANTENNA__17227__B1 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout262 net264 vssd1 vssd1 vccd1 vccd1 net262 sky130_fd_sc_hd__clkbuf_2
X_13940_ ag2.body\[82\] net197 _08154_ ag2.body\[74\] vssd1 vssd1 vccd1 vccd1 _00163_
+ sky130_fd_sc_hd__a22o_1
Xfanout273 _04306_ vssd1 vssd1 vccd1 vccd1 net273 sky130_fd_sc_hd__clkbuf_2
XANTENNA__19318__CLK clknet_leaf_105_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout284 net285 vssd1 vssd1 vccd1 vccd1 net284 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout67_X net67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout295 _07335_ vssd1 vssd1 vccd1 vccd1 net295 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_92_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17343__B net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13871_ _08139_ _08143_ vssd1 vssd1 vccd1 vccd1 _08145_ sky130_fd_sc_hd__or2_1
XFILLER_0_9_1101 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12768__A net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15610_ ag2.body\[459\] net123 _01620_ ag2.body\[451\] vssd1 vssd1 vccd1 vccd1 _00877_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_119_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12822_ net386 _07518_ vssd1 vssd1 vccd1 vccd1 _07612_ sky130_fd_sc_hd__nor2_1
XFILLER_0_119_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16590_ obsg2.obstacleArray\[68\] obsg2.obstacleArray\[69\] net446 vssd1 vssd1 vccd1
+ vccd1 _02269_ sky130_fd_sc_hd__mux2_1
XANTENNA__09468__B1 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1612 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_706 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15541_ ag2.body\[527\] net160 _01611_ ag2.body\[519\] vssd1 vssd1 vccd1 vccd1 _00817_
+ sky130_fd_sc_hd__a22o_1
X_12753_ net257 _07579_ _07580_ net2080 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[130\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_9_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16674__S net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11814__A2 net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18260_ _03699_ net37 obsg2.obstacleArray\[127\] vssd1 vssd1 vccd1 vccd1 _03769_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_96_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11704_ _06673_ _06674_ vssd1 vssd1 vccd1 vccd1 _06676_ sky130_fd_sc_hd__or2_1
XFILLER_0_56_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13016__A1 net240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15472_ ag2.body\[577\] net111 _01604_ ag2.body\[569\] vssd1 vssd1 vccd1 vccd1 _00755_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__19785__RESET_B net1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12684_ net245 _07547_ _07548_ net1824 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[93\]
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_117_3901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16753__A2 net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17950__A1 net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18174__B net35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17211_ ag2.body\[48\] net879 vssd1 vssd1 vccd1 vccd1 _02890_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_13_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14423_ _08580_ _08582_ _08583_ vssd1 vssd1 vccd1 vccd1 _08584_ sky130_fd_sc_hd__or3b_1
XFILLER_0_65_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18191_ net526 _03734_ vssd1 vssd1 vccd1 vccd1 _01343_ sky130_fd_sc_hd__and2_1
XFILLER_0_112_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11635_ net504 _06606_ _06607_ net759 vssd1 vssd1 vccd1 vccd1 _06608_ sky130_fd_sc_hd__a211o_1
XFILLER_0_0_1610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17142_ ag2.body\[268\] net965 vssd1 vssd1 vccd1 vccd1 _02821_ sky130_fd_sc_hd__xor2_1
X_14354_ net1037 ag2.body\[404\] vssd1 vssd1 vccd1 vccd1 _08515_ sky130_fd_sc_hd__xor2_1
X_11566_ net504 _06537_ _06538_ vssd1 vssd1 vccd1 vccd1 _06539_ sky130_fd_sc_hd__or3_1
XFILLER_0_107_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13319__A2 net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13305_ net235 _07835_ _07836_ net1718 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[426\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_64_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17073_ _02748_ _02749_ _02750_ _02751_ vssd1 vssd1 vccd1 vccd1 _02752_ sky130_fd_sc_hd__or4_1
X_10517_ _04023_ net1210 net757 ag2.body\[101\] _05485_ vssd1 vssd1 vccd1 vccd1 _05490_
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_52_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13111__B _07578_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14285_ _08439_ _08440_ _08441_ _08445_ vssd1 vssd1 vccd1 vccd1 _08446_ sky130_fd_sc_hd__or4b_1
XFILLER_0_126_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11497_ obsg2.obstacleArray\[114\] obsg2.obstacleArray\[118\] net512 vssd1 vssd1
+ vccd1 vccd1 _06470_ sky130_fd_sc_hd__mux2_1
X_16024_ _01695_ _01701_ vssd1 vssd1 vccd1 vccd1 _01703_ sky130_fd_sc_hd__or2_2
X_13236_ net382 net314 vssd1 vssd1 vccd1 vccd1 _07807_ sky130_fd_sc_hd__nand2_4
X_10448_ ag2.body\[453\] net1103 vssd1 vssd1 vccd1 vccd1 _05421_ sky130_fd_sc_hd__or2_1
XANTENNA__17518__B net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1616 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10173__D _05145_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15319__A _05036_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13167_ net278 _07773_ _07774_ net1994 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[350\]
+ sky130_fd_sc_hd__a22o_1
X_10379_ _05348_ _05349_ _05350_ _05351_ vssd1 vssd1 vccd1 vccd1 _05352_ sky130_fd_sc_hd__or4_1
XFILLER_0_0_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12118_ _07085_ _07087_ _07089_ net574 vssd1 vssd1 vccd1 vccd1 _07090_ sky130_fd_sc_hd__o22a_1
XFILLER_0_137_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17975_ net539 net380 net462 net486 vssd1 vssd1 vccd1 vccd1 _03597_ sky130_fd_sc_hd__and4_1
XANTENNA__12014__Y _06986_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13098_ net290 _07740_ _07741_ net2029 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[314\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_100_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19714_ clknet_leaf_133_clk _00658_ net1308 vssd1 vssd1 vccd1 vccd1 control.body\[672\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__15606__X _01620_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16926_ ag2.body\[372\] net963 vssd1 vssd1 vccd1 vccd1 _02605_ sky130_fd_sc_hd__xor2_1
X_12049_ img_gen.tracker.frame\[276\] net627 net554 img_gen.tracker.frame\[282\] _07020_
+ vssd1 vssd1 vccd1 vccd1 _07021_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_85_2901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19645_ clknet_leaf_128_clk _00589_ net1329 vssd1 vssd1 vccd1 vccd1 control.body\[747\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__17253__B net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16857_ ag2.body\[204\] net962 vssd1 vssd1 vccd1 vccd1 _02536_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_66_2322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_2333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16441__B2 net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_2344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15808_ ag2.body\[284\] net206 _01641_ ag2.body\[276\] vssd1 vssd1 vccd1 vccd1 _01054_
+ sky130_fd_sc_hd__a22o_1
X_16788_ net460 _02464_ _02465_ _02466_ net350 vssd1 vssd1 vccd1 vccd1 _02467_ sky130_fd_sc_hd__o311a_1
XFILLER_0_88_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19576_ clknet_leaf_116_clk _00520_ net1385 vssd1 vssd1 vccd1 vccd1 control.body\[822\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12058__A2 net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13255__A1 net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09459__B1 net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12397__B net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_2208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_62_2219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15739_ ag2.body\[351\] net211 _01633_ ag2.body\[343\] vssd1 vssd1 vccd1 vccd1 _00993_
+ sky130_fd_sc_hd__a22o_1
X_18527_ clknet_leaf_137_clk _00053_ net1298 vssd1 vssd1 vccd1 vccd1 img_gen.updater.commands.cmd_num\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__16729__C1 net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16584__S net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11805__A2 net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18365__A net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09260_ sound_gen.osc1.keepCounting sound_gen.posDetector1.N\[1\] vssd1 vssd1 vccd1
+ vccd1 _04285_ sky130_fd_sc_hd__and2b_2
XANTENNA__13007__A1 net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18835__CLK clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18458_ _05075_ _06173_ _03844_ _03946_ vssd1 vssd1 vccd1 vccd1 _03947_ sky130_fd_sc_hd__o31a_1
XANTENNA__16744__A2 net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09191_ ag2.body\[589\] vssd1 vssd1 vccd1 vccd1 _04216_ sky130_fd_sc_hd__inv_2
X_17409_ _03080_ _03081_ _03083_ _03085_ vssd1 vssd1 vccd1 vccd1 _03088_ sky130_fd_sc_hd__or4_1
XFILLER_0_117_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18389_ _03876_ _03877_ _03878_ vssd1 vssd1 vccd1 vccd1 _03879_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_79_2727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_79_2738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_794 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20420_ clknet_leaf_37_clk _01307_ net1349 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[56\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_15_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkload120 clknet_leaf_77_clk vssd1 vssd1 vccd1 vccd1 clkload120/X sky130_fd_sc_hd__clkbuf_8
X_20351_ clknet_leaf_139_clk _01242_ net1288 vssd1 vssd1 vccd1 vccd1 img_gen.updater.commands.rR1.rainbowRNG\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload131 clknet_leaf_72_clk vssd1 vssd1 vccd1 vccd1 clkload131/Y sky130_fd_sc_hd__bufinv_16
XANTENNA__15704__B1 _01629_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout114_A net219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20282_ clknet_leaf_36_clk control.divider.next_count\[3\] net1348 vssd1 vssd1 vccd1
+ vccd1 control.divider.count\[3\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_105_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17457__B1 net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14133__A net1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1023_A net1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11476__B net1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08975_ ag2.body\[66\] vssd1 vssd1 vccd1 vccd1 _04000_ sky130_fd_sc_hd__inv_2
XFILLER_0_122_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout483_A _02373_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold15 ag2.body\[6\] vssd1 vssd1 vccd1 vccd1 net1577 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10380__B net1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold26 img_gen.tracker.frame\[504\] vssd1 vssd1 vccd1 vccd1 net1588 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__16680__A1 net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold37 img_gen.tracker.frame\[448\] vssd1 vssd1 vccd1 vccd1 net1599 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13494__A1 net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold48 img_gen.tracker.frame\[424\] vssd1 vssd1 vccd1 vccd1 net1610 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold59 img_gen.tracker.frame\[0\] vssd1 vssd1 vccd1 vccd1 net1621 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__17163__B net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout369_X net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout748_A _04233_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1392_A net1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12049__A2 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09527_ net1226 control.body\[832\] vssd1 vssd1 vccd1 vccd1 _04500_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_45_1705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16494__S net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1180_X net1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout915_A net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_26_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09458_ net917 _04421_ vssd1 vssd1 vccd1 vccd1 _04431_ sky130_fd_sc_hd__nand2_1
XANTENNA__16507__B net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11009__B1 net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19196__RESET_B net1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout703_X net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09389_ _04363_ _04378_ vssd1 vssd1 vccd1 vccd1 _01408_ sky130_fd_sc_hd__nor2_1
XANTENNA__14308__A net1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_3230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11420_ net1171 control.body\[850\] vssd1 vssd1 vccd1 vccd1 _06393_ sky130_fd_sc_hd__xor2_1
X_20618_ net1561 vssd1 vssd1 vccd1 vccd1 gpio_oeb[30] sky130_fd_sc_hd__buf_2
XFILLER_0_46_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_75_clk_X clknet_leaf_75_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_3105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17696__B1 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11351_ ag2.body\[445\] net1103 vssd1 vssd1 vccd1 vccd1 _06324_ sky130_fd_sc_hd__nand2_1
XFILLER_0_62_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20549_ clknet_leaf_105_clk _01414_ _00023_ vssd1 vssd1 vccd1 vccd1 sound_gen.osc1.stayCount\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_39_1509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10302_ net1170 control.body\[698\] vssd1 vssd1 vccd1 vccd1 _05275_ sky130_fd_sc_hd__xor2_1
X_14070_ net814 ag2.body\[212\] ag2.body\[213\] net808 vssd1 vssd1 vccd1 vccd1 _08231_
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_120_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11282_ net1206 control.body\[1105\] vssd1 vssd1 vccd1 vccd1 _06255_ sky130_fd_sc_hd__xor2_1
XFILLER_0_120_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17448__B1 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13021_ net668 _07705_ vssd1 vssd1 vccd1 vccd1 _07706_ sky130_fd_sc_hd__nor2_1
XANTENNA__11667__A net1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10233_ _05178_ _05191_ _05192_ _05205_ vssd1 vssd1 vccd1 vccd1 _05206_ sky130_fd_sc_hd__o22a_1
XFILLER_0_105_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_89_3023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11732__A1 net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_3034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1002 net1005 vssd1 vssd1 vccd1 vccd1 net1002 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_7_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10164_ ag2.body\[582\] net1077 vssd1 vssd1 vccd1 vccd1 _05137_ sky130_fd_sc_hd__xor2_1
Xfanout1013 net1014 vssd1 vssd1 vccd1 vccd1 net1013 sky130_fd_sc_hd__buf_4
XANTENNA__16120__B1 net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_3045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10290__B net1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1024 ag2.randCord\[6\] vssd1 vssd1 vccd1 vccd1 net1024 sky130_fd_sc_hd__buf_4
XANTENNA__16669__S net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18708__CLK clknet_leaf_144_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1035 net1042 vssd1 vssd1 vccd1 vccd1 net1035 sky130_fd_sc_hd__buf_4
Xfanout1046 net1053 vssd1 vssd1 vccd1 vccd1 net1046 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_101_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17760_ net381 _03406_ _03410_ _03438_ vssd1 vssd1 vccd1 vccd1 _03439_ sky130_fd_sc_hd__and4_1
Xfanout1057 net1069 vssd1 vssd1 vccd1 vccd1 net1057 sky130_fd_sc_hd__buf_4
XFILLER_0_76_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10095_ net1229 control.body\[936\] vssd1 vssd1 vccd1 vccd1 _05068_ sky130_fd_sc_hd__xor2_1
XFILLER_0_41_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14972_ net2554 net159 net51 control.body\[1022\] vssd1 vssd1 vccd1 vccd1 _00312_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__08976__A ag2.body\[70\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1068 net1069 vssd1 vssd1 vccd1 vccd1 net1068 sky130_fd_sc_hd__buf_4
XANTENNA_clkbuf_leaf_13_clk_X clknet_leaf_13_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1079 net1082 vssd1 vssd1 vccd1 vccd1 net1079 sky130_fd_sc_hd__buf_4
X_16711_ obsg2.obstacleArray\[92\] obsg2.obstacleArray\[93\] obsg2.obstacleArray\[94\]
+ obsg2.obstacleArray\[95\] net957 net537 vssd1 vssd1 vccd1 vccd1 _02390_ sky130_fd_sc_hd__mux4_1
XFILLER_0_89_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13923_ ag2.body\[67\] net134 _08152_ ag2.body\[59\] vssd1 vssd1 vccd1 vccd1 _00148_
+ sky130_fd_sc_hd__a22o_1
X_17691_ ag2.body\[157\] net953 vssd1 vssd1 vccd1 vccd1 _03370_ sky130_fd_sc_hd__xor2_1
XFILLER_0_107_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12498__A _06724_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19290__CLK clknet_leaf_98_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16423__A1 net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16642_ net395 _02318_ _02320_ net359 vssd1 vssd1 vccd1 vccd1 _02321_ sky130_fd_sc_hd__a211o_1
X_19430_ clknet_leaf_111_clk _00374_ net1422 vssd1 vssd1 vccd1 vccd1 control.body\[964\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_138_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13854_ ag2.body\[17\] net116 _08134_ ag2.body\[9\] vssd1 vssd1 vccd1 vccd1 _00097_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_57_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_650 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12805_ net286 _07603_ _07604_ net2071 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[158\]
+ sky130_fd_sc_hd__a22o_1
X_16573_ net359 _02251_ _02248_ _02228_ vssd1 vssd1 vccd1 vccd1 _02252_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_18_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19361_ clknet_leaf_102_clk _00305_ net1439 vssd1 vssd1 vccd1 vccd1 control.body\[1039\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17801__B net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13785_ _08070_ _08092_ _08093_ vssd1 vssd1 vccd1 vccd1 _00069_ sky130_fd_sc_hd__and3_1
XFILLER_0_134_1378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10997_ _04118_ net1235 net752 ag2.body\[342\] _05969_ vssd1 vssd1 vccd1 vccd1 _05970_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_29_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11799__A1 _06661_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18312_ _03793_ _03807_ _03794_ vssd1 vssd1 vccd1 vccd1 _03808_ sky130_fd_sc_hd__a21o_1
X_15524_ _05304_ net65 vssd1 vssd1 vccd1 vccd1 _01610_ sky130_fd_sc_hd__and2_2
XFILLER_0_112_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12736_ net284 _07570_ _07571_ net1793 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[122\]
+ sky130_fd_sc_hd__a22o_1
X_19292_ clknet_leaf_98_clk _00236_ net1447 vssd1 vssd1 vccd1 vccd1 control.body\[1098\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_127_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16726__A2 net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18243_ obsg2.obstacleArray\[118\] _03760_ net527 vssd1 vssd1 vccd1 vccd1 _01369_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_112_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09600__A net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15455_ ag2.body\[594\] net86 _01602_ ag2.body\[586\] vssd1 vssd1 vccd1 vccd1 _00740_
+ sky130_fd_sc_hd__a22o_1
X_12667_ net603 _06639_ net435 net563 vssd1 vssd1 vccd1 vccd1 _07538_ sky130_fd_sc_hd__or4_1
XFILLER_0_127_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14406_ net825 ag2.body\[2\] net812 net927 _08566_ vssd1 vssd1 vccd1 vccd1 _08567_
+ sky130_fd_sc_hd__a221o_1
XANTENNA__13122__A net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18174_ _03611_ net35 vssd1 vssd1 vccd1 vccd1 _03726_ sky130_fd_sc_hd__nor2_1
X_11618_ net504 _06589_ _06590_ net1125 vssd1 vssd1 vccd1 vccd1 _06591_ sky130_fd_sc_hd__a211o_1
XFILLER_0_108_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15386_ control.body\[660\] net82 _01595_ net2419 vssd1 vssd1 vccd1 vccd1 _00678_
+ sky130_fd_sc_hd__a22o_1
X_12598_ net252 _07499_ _07500_ net1903 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[55\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_83_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18333__D1 net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17125_ ag2.body\[516\] net964 vssd1 vssd1 vccd1 vccd1 _02804_ sky130_fd_sc_hd__nand2_1
X_14337_ _08490_ _08493_ _08496_ _08497_ vssd1 vssd1 vccd1 vccd1 _08498_ sky130_fd_sc_hd__or4b_1
XFILLER_0_107_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11549_ net1174 _06491_ vssd1 vssd1 vccd1 vccd1 _06522_ sky130_fd_sc_hd__nor2_1
XFILLER_0_53_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1284 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold507 img_gen.tracker.frame\[575\] vssd1 vssd1 vccd1 vccd1 net2069 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_55_2001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold518 img_gen.tracker.frame\[130\] vssd1 vssd1 vccd1 vccd1 net2080 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_55_2012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_814 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17056_ _04007_ net968 net708 ag2.body\[77\] vssd1 vssd1 vccd1 vccd1 _02735_ sky130_fd_sc_hd__o22a_1
Xhold529 img_gen.tracker.frame\[562\] vssd1 vssd1 vccd1 vccd1 net2091 sky130_fd_sc_hd__dlygate4sd3_1
X_14268_ net1016 ag2.body\[14\] vssd1 vssd1 vccd1 vccd1 _08429_ sky130_fd_sc_hd__or2_1
XFILLER_0_64_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12680__B _06639_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17439__B1 net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16007_ _01684_ _01685_ vssd1 vssd1 vccd1 vccd1 _01686_ sky130_fd_sc_hd__nor2_1
XFILLER_0_0_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13219_ net383 _07630_ vssd1 vssd1 vccd1 vccd1 _07799_ sky130_fd_sc_hd__nor2_1
X_14199_ net1028 ag2.body\[365\] vssd1 vssd1 vccd1 vccd1 _08360_ sky130_fd_sc_hd__xor2_1
XANTENNA__13495__C _07813_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16662__B2 net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17958_ net318 _03583_ obsg2.obstacleArray\[10\] vssd1 vssd1 vccd1 vccd1 _03584_
+ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_68_2406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16909_ _02581_ _02582_ _02584_ _02587_ vssd1 vssd1 vccd1 vccd1 _02588_ sky130_fd_sc_hd__a211o_1
XFILLER_0_79_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17889_ _08141_ _03519_ _03528_ _03518_ vssd1 vssd1 vccd1 vccd1 _03529_ sky130_fd_sc_hd__o211ai_4
XANTENNA__17551__X _03230_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19628_ clknet_leaf_123_clk _00572_ net1409 vssd1 vssd1 vccd1 vccd1 control.body\[762\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__19783__CLK clknet_leaf_127_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19559_ clknet_leaf_115_clk _00503_ net1397 vssd1 vssd1 vccd1 vccd1 control.body\[837\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__18095__A net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1598 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09312_ sound_gen.osc1.count\[4\] sound_gen.osc1.count\[3\] _04321_ sound_gen.osc1.count\[5\]
+ vssd1 vssd1 vccd1 vccd1 _04330_ sky130_fd_sc_hd__a31o_1
XFILLER_0_87_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16717__A2 net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17914__A1 _01691_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09243_ net939 vssd1 vssd1 vccd1 vccd1 _04268_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout231_A net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11104__X _06077_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13032__A net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09174_ ag2.body\[543\] vssd1 vssd1 vccd1 vccd1 _04199_ sky130_fd_sc_hd__inv_2
XANTENNA__13400__A1 net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10375__B net1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17678__B1 net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20403_ clknet_leaf_25_clk _01290_ net1340 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[39\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__13951__A2 net191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1140_A net1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12871__A net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19163__CLK clknet_leaf_52_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1238_A ag2.y\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20334_ clknet_leaf_21_clk _01225_ net1364 vssd1 vssd1 vccd1 vccd1 ag2.apple_cord\[2\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_4_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout698_A _04268_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput16 net16 vssd1 vssd1 vccd1 vccd1 gpio_out[15] sky130_fd_sc_hd__buf_2
XANTENNA__11487__A net1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput27 net27 vssd1 vssd1 vccd1 vccd1 gpio_out[2] sky130_fd_sc_hd__buf_2
X_20265_ clknet_leaf_42_clk net1565 net1372 vssd1 vssd1 vccd1 vccd1 control.detect3.Q\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_102_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1026_X net1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10517__A2 net1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16997__B net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20196_ clknet_leaf_88_clk _01140_ net1454 vssd1 vssd1 vccd1 vccd1 ag2.body\[194\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__14798__A net1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout865_A net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout486_X net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16653__A1 net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08958_ ag2.body\[20\] vssd1 vssd1 vccd1 vccd1 _03983_ sky130_fd_sc_hd__inv_2
XANTENNA__13467__A1 net235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1008 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1395_X net1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17461__X _03140_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10920_ ag2.body\[456\] net1224 vssd1 vssd1 vccd1 vccd1 _05893_ sky130_fd_sc_hd__xor2_1
XANTENNA__17902__A net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16956__A2 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20101__Q ag2.body\[291\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout820_X net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17621__B net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10851_ _05820_ _05821_ _05823_ _05815_ vssd1 vssd1 vccd1 vccd1 _05824_ sky130_fd_sc_hd__a211o_1
XFILLER_0_6_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13570_ _04282_ _07940_ vssd1 vssd1 vccd1 vccd1 _07947_ sky130_fd_sc_hd__nand2_1
XFILLER_0_17_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10782_ net1073 control.body\[630\] vssd1 vssd1 vccd1 vccd1 _05755_ sky130_fd_sc_hd__xor2_1
XANTENNA__16708__A2 net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14719__A1 net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09420__A ag2.goodColl vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12521_ net315 _07457_ vssd1 vssd1 vccd1 vccd1 _07458_ sky130_fd_sc_hd__or2_1
XFILLER_0_52_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14719__B2 net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15916__B1 _01652_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_40_clk_A clknet_4_7__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15240_ control.body\[787\] net99 _01578_ control.body\[779\] vssd1 vssd1 vccd1 vccd1
+ _00549_ sky130_fd_sc_hd__a22o_1
X_12452_ _06658_ _06659_ _07299_ vssd1 vssd1 vccd1 vccd1 _07412_ sky130_fd_sc_hd__o21a_1
XANTENNA__10285__B net1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10205__A1 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11403_ ag2.body\[571\] net1150 vssd1 vssd1 vccd1 vccd1 _06376_ sky130_fd_sc_hd__or2_1
X_15171_ control.body\[854\] net94 _01570_ control.body\[846\] vssd1 vssd1 vccd1 vccd1
+ _00488_ sky130_fd_sc_hd__a22o_1
XFILLER_0_65_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13942__A2 net191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12383_ _07270_ _07279_ vssd1 vssd1 vccd1 vccd1 _07348_ sky130_fd_sc_hd__nor2_1
XFILLER_0_50_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10077__A1_N _05036_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14122_ net1037 ag2.body\[372\] vssd1 vssd1 vccd1 vccd1 _08283_ sky130_fd_sc_hd__xor2_1
X_11334_ net1146 control.body\[659\] vssd1 vssd1 vccd1 vccd1 _06307_ sky130_fd_sc_hd__xor2_1
XANTENNA__16341__B1 net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_55_clk_A clknet_4_12__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14053_ _08213_ _08206_ _08212_ vssd1 vssd1 vccd1 vccd1 _08214_ sky130_fd_sc_hd__or3b_1
X_18930_ clknet_leaf_140_clk img_gen.tracker.next_frame\[368\] net1290 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[368\] sky130_fd_sc_hd__dfrtp_1
X_11265_ _05543_ _06226_ _06232_ _06237_ vssd1 vssd1 vccd1 vccd1 _06238_ sky130_fd_sc_hd__o22a_1
XFILLER_0_120_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13004_ net669 _07697_ vssd1 vssd1 vccd1 vccd1 _07698_ sky130_fd_sc_hd__nor2_1
X_10216_ net1204 control.body\[993\] vssd1 vssd1 vccd1 vccd1 _05189_ sky130_fd_sc_hd__xnor2_1
XANTENNA__14301__A1_N net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18861_ clknet_leaf_18_clk img_gen.tracker.next_frame\[299\] net1323 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[299\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__16399__S net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11196_ net785 control.body\[872\] control.body\[877\] net754 vssd1 vssd1 vccd1 vccd1
+ _06169_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_118_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17812_ _03477_ _03478_ net927 vssd1 vssd1 vccd1 vccd1 _03480_ sky130_fd_sc_hd__a21o_1
X_10147_ _04640_ net634 vssd1 vssd1 vccd1 vccd1 _05120_ sky130_fd_sc_hd__nor2_1
XANTENNA__13458__A1 net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18792_ clknet_leaf_17_clk img_gen.tracker.next_frame\[230\] net1319 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[230\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__12499__Y _07445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_113_clk_A clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17743_ _02773_ _02779_ _02589_ vssd1 vssd1 vccd1 vccd1 _03422_ sky130_fd_sc_hd__o21a_1
X_14955_ net2513 net174 _01546_ control.body\[1038\] vssd1 vssd1 vccd1 vccd1 _00296_
+ sky130_fd_sc_hd__a22o_1
X_10078_ net890 net904 net900 net896 vssd1 vssd1 vccd1 vccd1 _05051_ sky130_fd_sc_hd__or4bb_4
XFILLER_0_136_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13117__A net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13906_ ag2.body\[52\] net119 _08150_ ag2.body\[44\] vssd1 vssd1 vccd1 vccd1 _00133_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__14407__B1 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17674_ ag2.body\[449\] net733 net690 ag2.body\[455\] _03350_ vssd1 vssd1 vccd1 vccd1
+ _03353_ sky130_fd_sc_hd__a221o_1
XFILLER_0_89_458 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14886_ control.body\[1096\] net180 _01539_ net2181 vssd1 vssd1 vccd1 vccd1 _00234_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__16947__A2 net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19413_ clknet_leaf_103_clk _00357_ net1432 vssd1 vssd1 vccd1 vccd1 control.body\[979\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_98_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16625_ obsg2.obstacleArray\[34\] net441 vssd1 vssd1 vccd1 vccd1 _02304_ sky130_fd_sc_hd__or2_1
X_13837_ _06636_ _08103_ _08129_ net1094 vssd1 vssd1 vccd1 vccd1 _00085_ sky130_fd_sc_hd__a22o_1
XANTENNA__17531__B net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_128_clk_A clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16556_ obsg2.obstacleArray\[108\] obsg2.obstacleArray\[109\] net442 vssd1 vssd1
+ vccd1 vccd1 _02235_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19344_ clknet_leaf_100_clk _00288_ net1443 vssd1 vssd1 vccd1 vccd1 control.body\[1054\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09601__Y _04574_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13768_ img_gen.updater.commands.count\[7\] _08081_ vssd1 vssd1 vccd1 vccd1 _08082_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_58_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12675__B net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12719_ net284 _07562_ _07563_ net1723 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[113\]
+ sky130_fd_sc_hd__a22o_1
X_15507_ ag2.body\[544\] net155 _01608_ ag2.body\[536\] vssd1 vssd1 vccd1 vccd1 _00786_
+ sky130_fd_sc_hd__a22o_1
X_16487_ net364 _02165_ _02164_ net363 vssd1 vssd1 vccd1 vccd1 _02166_ sky130_fd_sc_hd__o211a_1
XFILLER_0_57_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19275_ clknet_leaf_97_clk _00219_ net1450 vssd1 vssd1 vccd1 vccd1 control.body\[1113\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_0_clk clk vssd1 vssd1 vccd1 vccd1 clknet_0_clk sky130_fd_sc_hd__clkbuf_16
X_13699_ net923 track.highScore\[0\] track.highScore\[1\] vssd1 vssd1 vccd1 vccd1
+ _08040_ sky130_fd_sc_hd__a21o_1
XANTENNA__19186__CLK clknet_leaf_53_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18226_ _03668_ net40 vssd1 vssd1 vccd1 vccd1 _03752_ sky130_fd_sc_hd__nor2_1
X_15438_ ag2.body\[611\] net85 _01600_ ag2.body\[603\] vssd1 vssd1 vccd1 vccd1 _00725_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__10195__B net1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18157_ net523 _03717_ vssd1 vssd1 vccd1 vccd1 _01326_ sky130_fd_sc_hd__and2_1
X_15369_ net2521 net68 _01593_ control.body\[669\] vssd1 vssd1 vccd1 vccd1 _00663_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_87_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18081__C net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17108_ _03975_ net870 net960 _03978_ _02786_ vssd1 vssd1 vccd1 vccd1 _02787_ sky130_fd_sc_hd__a221o_1
Xhold304 img_gen.tracker.frame\[357\] vssd1 vssd1 vccd1 vccd1 net1866 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11035__A_N net1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18088_ obsg2.obstacleArray\[49\] _03674_ net527 vssd1 vssd1 vccd1 vccd1 _01300_
+ sky130_fd_sc_hd__o21a_1
Xhold315 img_gen.tracker.frame\[80\] vssd1 vssd1 vccd1 vccd1 net1877 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_48_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold326 sound_gen.dac1.dacCount\[1\] vssd1 vssd1 vccd1 vccd1 net1888 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold337 img_gen.tracker.frame\[526\] vssd1 vssd1 vccd1 vccd1 net1899 sky130_fd_sc_hd__dlygate4sd3_1
Xhold348 img_gen.tracker.frame\[240\] vssd1 vssd1 vccd1 vccd1 net1910 sky130_fd_sc_hd__dlygate4sd3_1
X_17039_ _04029_ net878 net713 ag2.body\[124\] vssd1 vssd1 vccd1 vccd1 _02718_ sky130_fd_sc_hd__a22o_1
XFILLER_0_110_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09930_ net890 _04792_ vssd1 vssd1 vccd1 vccd1 _04903_ sky130_fd_sc_hd__nor2_4
XFILLER_0_1_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold359 img_gen.tracker.frame\[275\] vssd1 vssd1 vccd1 vccd1 net1921 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_15_Right_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13697__A1 _04425_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20050_ clknet_leaf_72_clk _00994_ net1503 vssd1 vssd1 vccd1 vccd1 ag2.body\[336\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_110_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout806 net807 vssd1 vssd1 vccd1 vccd1 net806 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_1_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09861_ ag2.body\[154\] net1185 vssd1 vssd1 vccd1 vccd1 _04834_ sky130_fd_sc_hd__xor2_1
Xfanout817 net819 vssd1 vssd1 vccd1 vccd1 net817 sky130_fd_sc_hd__buf_4
XFILLER_0_106_1299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout828 net830 vssd1 vssd1 vccd1 vccd1 net828 sky130_fd_sc_hd__buf_4
Xfanout839 _03965_ vssd1 vssd1 vccd1 vccd1 net839 sky130_fd_sc_hd__buf_4
XANTENNA__16096__C1 net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17832__A0 net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13449__A1 net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09792_ _04756_ _04757_ _04762_ _04764_ vssd1 vssd1 vccd1 vccd1 _04765_ sky130_fd_sc_hd__or4_1
Xhold1004 control.body\[805\] vssd1 vssd1 vccd1 vccd1 net2566 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_84_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1015 control.body\[1082\] vssd1 vssd1 vccd1 vccd1 net2577 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1026 control.body\[844\] vssd1 vssd1 vccd1 vccd1 net2588 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1037 control.body\[770\] vssd1 vssd1 vccd1 vccd1 net2599 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1048 control.body\[842\] vssd1 vssd1 vccd1 vccd1 net2610 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_84_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1059 control.body\[774\] vssd1 vssd1 vccd1 vccd1 net2621 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout181_A net182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12121__A1 net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout279_A _07335_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13027__A net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1528 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16938__A2 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11880__B1 net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1090_A net1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_992 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12866__A net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_24_Right_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout446_A net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1188_A net1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09240__A net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16057__B net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout613_A net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout234_X net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1355_A net1356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_1435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__20304__RESET_B net1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09226_ control.body\[1017\] vssd1 vssd1 vccd1 vccd1 _04251_ sky130_fd_sc_hd__inv_2
XFILLER_0_90_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18553__CLK clknet_leaf_37_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11769__X _06741_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout401_X net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09894__B net1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09157_ ag2.body\[501\] vssd1 vssd1 vccd1 vccd1 _04182_ sky130_fd_sc_hd__inv_2
XFILLER_0_90_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13924__A2 net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1143_X net1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09088_ ag2.body\[328\] vssd1 vssd1 vccd1 vccd1 _04113_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout982_A ag2.randCord\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10833__B net1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_33_Right_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_1018 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20317_ clknet_leaf_44_clk obsrand1.next_randY\[3\] net1381 vssd1 vssd1 vccd1 vccd1
+ ag2.randCord\[3\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_13_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1310_X net1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold860 control.body\[756\] vssd1 vssd1 vccd1 vccd1 net2422 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout94_A net100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold871 control.body\[867\] vssd1 vssd1 vccd1 vccd1 net2433 sky130_fd_sc_hd__dlygate4sd3_1
Xhold882 control.body\[647\] vssd1 vssd1 vccd1 vccd1 net2444 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11050_ ag2.body\[384\] net784 net1080 _04141_ _06022_ vssd1 vssd1 vccd1 vccd1 _06023_
+ sky130_fd_sc_hd__o221a_1
Xhold893 _00633_ vssd1 vssd1 vccd1 vccd1 net2455 sky130_fd_sc_hd__dlygate4sd3_1
X_20248_ clknet_leaf_68_clk _01192_ net1496 vssd1 vssd1 vccd1 vccd1 ag2.body\[150\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA_fanout770_X net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout868_X net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10001_ net1170 control.body\[730\] vssd1 vssd1 vccd1 vccd1 _04974_ sky130_fd_sc_hd__or2_1
XFILLER_0_102_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1387 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11360__A1_N net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20179_ clknet_leaf_87_clk _01123_ net1460 vssd1 vssd1 vccd1 vccd1 ag2.body\[209\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_137_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11664__B net1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12112__A1 net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14740_ net978 ag2.body\[331\] vssd1 vssd1 vccd1 vccd1 _08901_ sky130_fd_sc_hd__xor2_1
XFILLER_0_93_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11952_ img_gen.tracker.frame\[112\] net601 net586 img_gen.tracker.frame\[118\] vssd1
+ vssd1 vccd1 vccd1 _06924_ sky130_fd_sc_hd__o22a_1
XFILLER_0_58_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16929__A2 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_42_Right_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14975__B net59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10903_ net1118 control.body\[676\] vssd1 vssd1 vccd1 vccd1 _05876_ sky130_fd_sc_hd__xor2_1
X_14671_ net990 _04139_ ag2.body\[386\] net826 _08831_ vssd1 vssd1 vccd1 vccd1 _08832_
+ sky130_fd_sc_hd__a221o_1
X_11883_ net576 _06854_ vssd1 vssd1 vccd1 vccd1 _06855_ sky130_fd_sc_hd__nand2_1
XANTENNA__12776__A net225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_3974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16410_ obsg2.obstacleArray\[96\] obsg2.obstacleArray\[97\] net452 vssd1 vssd1 vccd1
+ vccd1 _02089_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13622_ net2083 _07987_ _07989_ vssd1 vssd1 vccd1 vccd1 control.divider.next_count\[7\]
+ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_120_3985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_3996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10834_ ag2.body\[309\] net1115 vssd1 vssd1 vccd1 vccd1 _05807_ sky130_fd_sc_hd__nand2_1
X_17390_ _03066_ _03067_ _03068_ vssd1 vssd1 vccd1 vccd1 _03069_ sky130_fd_sc_hd__or3b_1
XFILLER_0_13_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_3395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16341_ net370 _02019_ net368 vssd1 vssd1 vccd1 vccd1 _02020_ sky130_fd_sc_hd__o21a_1
XANTENNA__10426__A1 net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13553_ ssdec1.in\[2\] _07931_ _07934_ _04282_ vssd1 vssd1 vccd1 vccd1 _07935_ sky130_fd_sc_hd__o211a_1
X_10765_ net751 control.body\[894\] _05735_ _05736_ _05737_ vssd1 vssd1 vccd1 vccd1
+ _05738_ sky130_fd_sc_hd__a2111o_1
XANTENNA__20045__RESET_B net1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20186__CLK clknet_leaf_88_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12504_ net227 _07446_ _07447_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[14\]
+ sky130_fd_sc_hd__o21bai_1
X_19060_ clknet_leaf_9_clk img_gen.tracker.next_frame\[498\] net1271 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[498\] sky130_fd_sc_hd__dfrtp_1
X_16272_ obsg2.obstacleArray\[26\] net411 vssd1 vssd1 vccd1 vccd1 _01951_ sky130_fd_sc_hd__or2_1
X_13484_ net1700 _07905_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[536\]
+ sky130_fd_sc_hd__and2_1
XFILLER_0_70_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10696_ _05656_ _05657_ _05664_ _05668_ vssd1 vssd1 vccd1 vccd1 _05669_ sky130_fd_sc_hd__o22a_2
XANTENNA__18182__B net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18011_ net45 _03622_ vssd1 vssd1 vccd1 vccd1 _03623_ sky130_fd_sc_hd__nor2_1
XFILLER_0_129_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15223_ net2642 net93 _01576_ control.body\[796\] vssd1 vssd1 vccd1 vccd1 _00534_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11679__X _06651_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12435_ _07222_ _07279_ _07277_ vssd1 vssd1 vccd1 vccd1 _07396_ sky130_fd_sc_hd__o21bai_1
XANTENNA__17106__A2 net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_51_Right_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10729__A2 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15154_ control.body\[871\] net106 _01568_ control.body\[863\] vssd1 vssd1 vccd1
+ vccd1 _00473_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_114_3789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12366_ net241 vssd1 vssd1 vccd1 vccd1 _07332_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_136_Right_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10743__B net1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14105_ net970 ag2.body\[587\] vssd1 vssd1 vccd1 vccd1 _08266_ sky130_fd_sc_hd__xnor2_1
XANTENNA__17366__X _03045_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12661__D net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11317_ net904 _04601_ _05074_ _05192_ vssd1 vssd1 vccd1 vccd1 _06290_ sky130_fd_sc_hd__o31a_1
X_19962_ clknet_leaf_62_clk _00906_ net1470 vssd1 vssd1 vccd1 vccd1 ag2.body\[424\]
+ sky130_fd_sc_hd__dfrtp_4
X_15085_ net2581 net148 _01562_ net2264 vssd1 vssd1 vccd1 vccd1 _00410_ sky130_fd_sc_hd__a22o_1
X_12297_ _07218_ _07221_ vssd1 vssd1 vccd1 vccd1 _07264_ sky130_fd_sc_hd__and2_1
X_14036_ net1004 ag2.body\[496\] vssd1 vssd1 vccd1 vccd1 _08197_ sky130_fd_sc_hd__nand2_1
X_18913_ clknet_leaf_3_clk img_gen.tracker.next_frame\[351\] net1258 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[351\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_103_1439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11248_ ag2.body\[196\] net1138 vssd1 vssd1 vccd1 vccd1 _06221_ sky130_fd_sc_hd__or2_1
X_19893_ clknet_leaf_85_clk _00837_ net1462 vssd1 vssd1 vccd1 vccd1 ag2.body\[499\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_129_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16617__A1 net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18844_ clknet_leaf_4_clk img_gen.tracker.next_frame\[282\] net1277 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[282\] sky130_fd_sc_hd__dfrtp_1
X_11179_ _05451_ _06135_ _06137_ _06138_ _06151_ vssd1 vssd1 vccd1 vccd1 _06152_ sky130_fd_sc_hd__o32a_1
XANTENNA__10362__B1 _05323_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18775_ clknet_leaf_16_clk img_gen.tracker.next_frame\[213\] net1321 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[213\] sky130_fd_sc_hd__dfrtp_1
X_15987_ _01668_ _01670_ vssd1 vssd1 vccd1 vccd1 _01671_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_60_Right_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19228__RESET_B net1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17726_ obsg2.obstacleArray\[132\] obsg2.obstacleArray\[133\] obsg2.obstacleArray\[134\]
+ obsg2.obstacleArray\[135\] net958 net538 vssd1 vssd1 vccd1 vccd1 _03405_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_19_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14938_ control.body\[1063\] net168 _01544_ net2179 vssd1 vssd1 vccd1 vccd1 _00281_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_72_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14885__B _04861_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09612__X _04585_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17261__B net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17657_ ag2.body\[107\] net856 vssd1 vssd1 vccd1 vccd1 _03336_ sky130_fd_sc_hd__xor2_1
XANTENNA__16896__A2_N net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11862__B1 net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14869_ net2123 net181 _01537_ control.body\[1105\] vssd1 vssd1 vccd1 vccd1 _00219_
+ sky130_fd_sc_hd__a22o_1
X_16608_ obsg2.obstacleArray\[92\] obsg2.obstacleArray\[93\] net445 vssd1 vssd1 vccd1
+ vccd1 _02287_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17588_ _03263_ _03264_ _03266_ vssd1 vssd1 vccd1 vccd1 _03267_ sky130_fd_sc_hd__and3b_1
XANTENNA__10918__B net1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15997__A net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19327_ clknet_leaf_104_clk _00271_ net1432 vssd1 vssd1 vccd1 vccd1 control.body\[1069\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16592__S net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16539_ obsg2.obstacleArray\[98\] obsg2.obstacleArray\[99\] net441 vssd1 vssd1 vccd1
+ vccd1 _02218_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_1529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19821__CLK clknet_leaf_124_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19258_ clknet_leaf_73_clk _00202_ net1500 vssd1 vssd1 vccd1 vccd1 ag2.body\[121\]
+ sky130_fd_sc_hd__dfrtp_4
X_09011_ ag2.body\[136\] vssd1 vssd1 vccd1 vccd1 _04036_ sky130_fd_sc_hd__inv_2
XFILLER_0_14_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18209_ net523 _03743_ vssd1 vssd1 vccd1 vccd1 _01352_ sky130_fd_sc_hd__and2_1
XFILLER_0_6_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19189_ clknet_leaf_20_clk _00133_ net1366 vssd1 vssd1 vccd1 vccd1 ag2.body\[52\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_115_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11917__A1 net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold101 img_gen.tracker.frame\[45\] vssd1 vssd1 vccd1 vccd1 net1663 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_130_4281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold112 img_gen.tracker.frame\[291\] vssd1 vssd1 vccd1 vccd1 net1674 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_130_4292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10653__B net1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold123 img_gen.tracker.frame\[553\] vssd1 vssd1 vccd1 vccd1 net1685 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_48_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12590__A1 net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_103_Right_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold134 img_gen.tracker.frame\[345\] vssd1 vssd1 vccd1 vccd1 net1696 sky130_fd_sc_hd__dlygate4sd3_1
Xhold145 img_gen.tracker.frame\[534\] vssd1 vssd1 vccd1 vccd1 net1707 sky130_fd_sc_hd__dlygate4sd3_1
Xhold156 img_gen.tracker.frame\[426\] vssd1 vssd1 vccd1 vccd1 net1718 sky130_fd_sc_hd__dlygate4sd3_1
Xhold167 img_gen.tracker.frame\[94\] vssd1 vssd1 vccd1 vccd1 net1729 sky130_fd_sc_hd__dlygate4sd3_1
X_09913_ ag2.body\[135\] net1067 vssd1 vssd1 vccd1 vccd1 _04886_ sky130_fd_sc_hd__xor2_1
X_20102_ clknet_leaf_78_clk _01046_ net1486 vssd1 vssd1 vccd1 vccd1 ag2.body\[292\]
+ sky130_fd_sc_hd__dfrtp_4
Xhold178 img_gen.tracker.frame\[453\] vssd1 vssd1 vccd1 vccd1 net1740 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1528 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13964__B net67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold189 img_gen.tracker.frame\[441\] vssd1 vssd1 vccd1 vccd1 net1751 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout603 net605 vssd1 vssd1 vccd1 vccd1 net603 sky130_fd_sc_hd__clkbuf_4
Xfanout614 net615 vssd1 vssd1 vccd1 vccd1 net614 sky130_fd_sc_hd__clkbuf_2
XANTENNA__11145__A2 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_1636 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12946__A_N _07483_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout625 net626 vssd1 vssd1 vccd1 vccd1 net625 sky130_fd_sc_hd__clkbuf_4
X_20033_ clknet_leaf_67_clk _00977_ net1473 vssd1 vssd1 vccd1 vccd1 ag2.body\[367\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_0_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout636 _04492_ vssd1 vssd1 vccd1 vccd1 net636 sky130_fd_sc_hd__buf_4
XANTENNA__17805__B1 net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09844_ _04800_ _04805_ _04815_ _04816_ vssd1 vssd1 vccd1 vccd1 _04817_ sky130_fd_sc_hd__or4_2
Xfanout647 net648 vssd1 vssd1 vccd1 vccd1 net647 sky130_fd_sc_hd__buf_2
XANTENNA__14141__A net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout658 net659 vssd1 vssd1 vccd1 vccd1 net658 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__14619__B1 ag2.body\[62\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_13_Left_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1103_A net1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout669 net674 vssd1 vssd1 vccd1 vccd1 net669 sky130_fd_sc_hd__clkbuf_2
X_09775_ ag2.body\[234\] net1182 vssd1 vssd1 vccd1 vccd1 _04748_ sky130_fd_sc_hd__xor2_1
XANTENNA__16767__S net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout563_A net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_4096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15831__A2 net204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_1_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09510__A2 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17171__B net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout351_X net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09889__B net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12596__A net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout730_A net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout828_A net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1093_X net1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout449_X net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17584__A2 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15595__A1 ag2.body\[478\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10828__B net1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_22_Left_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout616_X net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13070__A2 _07726_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_10__f_clk_X clknet_4_10__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10550_ ag2.body\[227\] net1159 vssd1 vssd1 vccd1 vccd1 _05523_ sky130_fd_sc_hd__nand2_1
XFILLER_0_106_213 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15898__A2 net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09209_ net1047 vssd1 vssd1 vccd1 vccd1 _04234_ sky130_fd_sc_hd__inv_2
XFILLER_0_51_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10481_ ag2.body\[590\] net1074 vssd1 vssd1 vccd1 vccd1 _05454_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_66_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12220_ img_gen.updater.commands.count\[4\] img_gen.updater.commands.count\[3\] _07189_
+ vssd1 vssd1 vccd1 vccd1 _07190_ sky130_fd_sc_hd__or3_1
XANTENNA__13220__A net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12030__B1 net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout985_X net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12151_ img_gen.tracker.frame\[432\] net613 net541 img_gen.tracker.frame\[438\] vssd1
+ vssd1 vccd1 vccd1 _07123_ sky130_fd_sc_hd__o22a_1
XANTENNA__12481__D _07312_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14858__B1 _08413_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11102_ _04152_ net1104 net749 ag2.body\[430\] _06071_ vssd1 vssd1 vccd1 vccd1 _06075_
+ sky130_fd_sc_hd__o221a_1
XANTENNA__13874__B net56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12082_ img_gen.tracker.frame\[315\] net611 net594 img_gen.tracker.frame\[321\] _07053_
+ vssd1 vssd1 vccd1 vccd1 _07054_ sky130_fd_sc_hd__a221o_1
Xhold690 control.body\[1049\] vssd1 vssd1 vccd1 vccd1 net2252 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_31_Left_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11675__A _06638_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11033_ net1207 control.body\[1041\] vssd1 vssd1 vccd1 vccd1 _06006_ sky130_fd_sc_hd__nand2b_1
X_15910_ _05544_ net54 vssd1 vssd1 vccd1 vccd1 _01652_ sky130_fd_sc_hd__nor2_4
X_16890_ ag2.body\[212\] net964 vssd1 vssd1 vccd1 vccd1 _02569_ sky130_fd_sc_hd__nand2_1
XFILLER_0_60_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16075__A2 net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15841_ ag2.body\[250\] net181 _01644_ ag2.body\[242\] vssd1 vssd1 vccd1 vccd1 _01084_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_137_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_107_3582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12097__B1 net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18560_ clknet_leaf_132_clk _00086_ net1304 vssd1 vssd1 vccd1 vccd1 ag2.x\[2\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_38_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_107_3593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15772_ ag2.body\[316\] net208 _01637_ ag2.body\[308\] vssd1 vssd1 vccd1 vccd1 _01022_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_77_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12984_ net278 _07686_ _07687_ net1774 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[254\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__18221__B1 net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17511_ ag2.body\[584\] net879 vssd1 vssd1 vccd1 vccd1 _03190_ sky130_fd_sc_hd__xor2_1
XFILLER_0_115_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_3457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17081__B net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11935_ img_gen.tracker.frame\[190\] net587 vssd1 vssd1 vccd1 vccd1 _06907_ sky130_fd_sc_hd__or2_1
XFILLER_0_38_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14723_ _08866_ _08867_ _08871_ _08883_ vssd1 vssd1 vccd1 vccd1 _08884_ sky130_fd_sc_hd__o31a_1
XANTENNA__11844__B1 net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_103_3468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18491_ net1516 net1510 vssd1 vssd1 vccd1 vccd1 _00022_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_103_3479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14654_ net839 ag2.body\[145\] _04042_ net1040 _08814_ vssd1 vssd1 vccd1 vccd1 _08815_
+ sky130_fd_sc_hd__a221o_1
X_17442_ ag2.body\[377\] net872 vssd1 vssd1 vccd1 vccd1 _03121_ sky130_fd_sc_hd__xor2_1
X_11866_ img_gen.tracker.frame\[271\] net548 vssd1 vssd1 vccd1 vccd1 _06838_ sky130_fd_sc_hd__or2_1
XANTENNA__15586__B2 ag2.body\[478\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10738__B net1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13605_ control.divider.count\[20\] _07949_ _07979_ control.divider.count\[21\] control.divider.count\[22\]
+ vssd1 vssd1 vccd1 vccd1 _07980_ sky130_fd_sc_hd__a2111oi_1
XFILLER_0_129_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10817_ net1136 control.body\[1092\] vssd1 vssd1 vccd1 vccd1 _05790_ sky130_fd_sc_hd__xor2_1
X_17373_ _03014_ _03015_ _03026_ _03974_ _03016_ vssd1 vssd1 vccd1 vccd1 _03052_ sky130_fd_sc_hd__o221a_1
X_14585_ net1032 ag2.body\[85\] vssd1 vssd1 vccd1 vccd1 _08746_ sky130_fd_sc_hd__xor2_1
XFILLER_0_89_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11797_ net563 _06766_ net467 vssd1 vssd1 vccd1 vccd1 _06769_ sky130_fd_sc_hd__a21o_1
XANTENNA__13061__A2 _07723_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19112_ clknet_leaf_0_clk img_gen.tracker.next_frame\[550\] net1244 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[550\] sky130_fd_sc_hd__dfrtp_1
X_16324_ _02001_ _02002_ net416 vssd1 vssd1 vccd1 vccd1 _02003_ sky130_fd_sc_hd__mux2_1
X_13536_ net2086 net655 _07925_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[568\]
+ sky130_fd_sc_hd__and3_1
X_10748_ ag2.body\[497\] net1213 vssd1 vssd1 vccd1 vccd1 _05721_ sky130_fd_sc_hd__xor2_1
XFILLER_0_137_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16255_ obsg2.obstacleArray\[58\] obsg2.obstacleArray\[59\] net407 vssd1 vssd1 vccd1
+ vccd1 _01934_ sky130_fd_sc_hd__mux2_1
X_19043_ clknet_leaf_7_clk img_gen.tracker.next_frame\[481\] net1268 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[481\] sky130_fd_sc_hd__dfrtp_1
X_13467_ net235 _07898_ _07899_ net1882 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[525\]
+ sky130_fd_sc_hd__a22o_1
X_10679_ ag2.body\[349\] net1113 vssd1 vssd1 vccd1 vccd1 _05652_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_11_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_1573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_11_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15206_ net2632 net92 _01574_ net2176 vssd1 vssd1 vccd1 vccd1 _00519_ sky130_fd_sc_hd__a22o_1
XFILLER_0_35_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12418_ _06525_ _07379_ vssd1 vssd1 vccd1 vccd1 _07380_ sky130_fd_sc_hd__nor2_1
X_16186_ _01863_ _01864_ net373 vssd1 vssd1 vccd1 vccd1 _01865_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13398_ net238 net312 _07551_ _07872_ net1662 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[483\]
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_45_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19224__CLK clknet_leaf_75_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12572__A1 net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_290 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15137_ _05051_ _06173_ net50 vssd1 vssd1 vccd1 vccd1 _01567_ sky130_fd_sc_hd__o21a_2
X_12349_ net317 _07315_ vssd1 vssd1 vccd1 vccd1 _07316_ sky130_fd_sc_hd__and2_1
XFILLER_0_49_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_1372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19945_ clknet_leaf_46_clk _00889_ net1376 vssd1 vssd1 vccd1 vccd1 ag2.body\[455\]
+ sky130_fd_sc_hd__dfrtp_4
X_15068_ net2245 net149 _01560_ control.body\[929\] vssd1 vssd1 vccd1 vccd1 _00395_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_71_2479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14019_ net999 _04161_ ag2.body\[458\] net825 _08173_ vssd1 vssd1 vccd1 vccd1 _08180_
+ sky130_fd_sc_hd__o221a_1
XANTENNA__11585__A net1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19876_ clknet_leaf_87_clk _00820_ net1479 vssd1 vssd1 vccd1 vccd1 ag2.body\[514\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__19374__CLK clknet_leaf_102_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16066__A2 net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18460__B1 net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18827_ clknet_leaf_4_clk img_gen.tracker.next_frame\[265\] net1262 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[265\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__16471__C1 net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09560_ _04525_ _04530_ _04531_ _04532_ vssd1 vssd1 vccd1 vccd1 _04533_ sky130_fd_sc_hd__or4_1
XANTENNA__12088__B1 net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18758_ clknet_leaf_15_clk img_gen.tracker.next_frame\[196\] net1313 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[196\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_88_2998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17709_ obsg2.obstacleArray\[128\] obsg2.obstacleArray\[129\] net448 vssd1 vssd1
+ vccd1 vccd1 _03388_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09491_ ag2.body\[370\] net1176 vssd1 vssd1 vccd1 vccd1 _04464_ sky130_fd_sc_hd__xor2_1
XANTENNA__11835__B1 net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18689_ clknet_leaf_28_clk img_gen.tracker.next_frame\[127\] net1335 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[127\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__15026__B1 _01555_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17566__A2 net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09502__B net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16774__B1 net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10648__B net1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkload83_A clknet_leaf_124_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16038__D net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13052__A2 _07718_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout144_A net219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20582_ clknet_leaf_107_clk _01439_ _00046_ vssd1 vssd1 vccd1 vccd1 sound_gen.osc1.count\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_132_4343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_132_4354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14001__A1 net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10664__A net1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_1571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14136__A net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14001__B2 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1053_A net1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout409_A net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_1582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11479__B net1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10383__B net1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1220_A net1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17166__B net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout400 _02064_ vssd1 vssd1 vccd1 vccd1 net400 sky130_fd_sc_hd__buf_2
XFILLER_0_26_1580 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout680_A net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout411 net412 vssd1 vssd1 vccd1 vccd1 net411 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11118__A2 _06075_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1409 net1415 vssd1 vssd1 vccd1 vccd1 net1409 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_121_1347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout399_X net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout422 net423 vssd1 vssd1 vccd1 vccd1 net422 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout778_A net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17734__X _03413_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout433 _01705_ vssd1 vssd1 vccd1 vccd1 net433 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_1444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_54_1976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout444 net445 vssd1 vssd1 vccd1 vccd1 net444 sky130_fd_sc_hd__clkbuf_4
Xfanout455 net459 vssd1 vssd1 vccd1 vccd1 net455 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout1106_X net1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout466 _06660_ vssd1 vssd1 vccd1 vccd1 net466 sky130_fd_sc_hd__clkbuf_4
X_20016_ clknet_leaf_59_clk _00960_ net1467 vssd1 vssd1 vccd1 vccd1 ag2.body\[382\]
+ sky130_fd_sc_hd__dfrtp_4
X_09827_ _04796_ _04797_ _04798_ _04799_ vssd1 vssd1 vccd1 vccd1 _04800_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_35_1386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_1397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout488 net489 vssd1 vssd1 vccd1 vccd1 net488 sky130_fd_sc_hd__buf_4
XANTENNA_fanout945_A obsg2.randCord\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout499 _01711_ vssd1 vssd1 vccd1 vccd1 net499 sky130_fd_sc_hd__buf_4
XANTENNA__18741__CLK clknet_leaf_141_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout566_X net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09758_ ag2.body\[214\] net1089 vssd1 vssd1 vccd1 vccd1 _04731_ sky130_fd_sc_hd__nand2_1
XANTENNA__12079__B1 _06660_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20390__RESET_B net1374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout57_A net62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18203__B1 net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11826__B1 net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout733_X net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09689_ ag2.body\[64\] net1233 vssd1 vssd1 vccd1 vccd1 _04662_ sky130_fd_sc_hd__xor2_1
XFILLER_0_119_1298 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15017__B1 _01553_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11720_ img_gen.tracker.frame\[218\] net623 net607 img_gen.tracker.frame\[221\] vssd1
+ vssd1 vccd1 vccd1 _06692_ sky130_fd_sc_hd__o22a_1
XANTENNA__11921__S0 net1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16765__B1 net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11661__C _06623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10558__B net1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11651_ net1167 _06557_ vssd1 vssd1 vccd1 vccd1 _06624_ sky130_fd_sc_hd__nor2_1
XFILLER_0_138_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_1562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14240__A1 net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout40 _03702_ vssd1 vssd1 vccd1 vccd1 net40 sky130_fd_sc_hd__clkbuf_4
XANTENNA__14240__B2 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout51 _01536_ vssd1 vssd1 vccd1 vccd1 net51 sky130_fd_sc_hd__clkbuf_4
Xfanout62 _08132_ vssd1 vssd1 vccd1 vccd1 net62 sky130_fd_sc_hd__buf_6
X_10602_ net1134 control.body\[988\] vssd1 vssd1 vccd1 vccd1 _05575_ sky130_fd_sc_hd__xor2_1
XFILLER_0_25_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14370_ _08528_ _08529_ _08530_ vssd1 vssd1 vccd1 vccd1 _08531_ sky130_fd_sc_hd__nand3b_4
X_11582_ _06511_ _06541_ _06554_ _06528_ vssd1 vssd1 vccd1 vccd1 _06555_ sky130_fd_sc_hd__a31o_1
XFILLER_0_80_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout73 net74 vssd1 vssd1 vccd1 vccd1 net73 sky130_fd_sc_hd__buf_2
Xfanout84 net85 vssd1 vssd1 vccd1 vccd1 net84 sky130_fd_sc_hd__buf_2
Xfanout95 net100 vssd1 vssd1 vccd1 vccd1 net95 sky130_fd_sc_hd__clkbuf_2
XANTENNA__12773__B net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19247__CLK clknet_leaf_83_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13321_ net275 net316 _07495_ _07841_ net1839 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[437\]
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_36_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10533_ _05502_ _05503_ _05504_ _05505_ vssd1 vssd1 vccd1 vccd1 _05506_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_115_3840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14046__A net1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_1046 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17190__B1 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_9__f_clk_X clknet_4_9__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16040_ net502 net463 net498 _01718_ vssd1 vssd1 vccd1 vccd1 _01719_ sky130_fd_sc_hd__a31o_1
XFILLER_0_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_111_3704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13252_ _06724_ net341 vssd1 vssd1 vccd1 vccd1 _07814_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_111_3715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10464_ net1231 control.body\[1008\] vssd1 vssd1 vccd1 vccd1 _05437_ sky130_fd_sc_hd__xor2_1
XANTENNA__10293__B net1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16532__Y _02211_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12203_ _06986_ _07149_ _07174_ _06634_ vssd1 vssd1 vccd1 vccd1 _07175_ sky130_fd_sc_hd__o211a_1
XANTENNA__11957__X _06929_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13183_ img_gen.tracker.frame\[359\] net644 _07781_ vssd1 vssd1 vccd1 vccd1 _07782_
+ sky130_fd_sc_hd__and3_1
X_10395_ _05366_ _05367_ _05365_ vssd1 vssd1 vccd1 vccd1 _05368_ sky130_fd_sc_hd__a21o_1
XANTENNA__19397__CLK clknet_leaf_111_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16296__A2 net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11676__Y _06648_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12134_ img_gen.tracker.frame\[480\] net618 net546 img_gen.tracker.frame\[486\] vssd1
+ vssd1 vccd1 vccd1 _07106_ sky130_fd_sc_hd__o22a_1
X_17991_ net345 net299 _03557_ vssd1 vssd1 vccd1 vccd1 _03608_ sky130_fd_sc_hd__and3_1
XFILLER_0_27_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19730_ clknet_leaf_128_clk _00674_ net1329 vssd1 vssd1 vccd1 vccd1 control.body\[656\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_104_1578 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12065_ net575 _07030_ _07028_ net468 vssd1 vssd1 vccd1 vccd1 _07037_ sky130_fd_sc_hd__a211o_1
X_16942_ _02612_ _02613_ _02615_ _02620_ vssd1 vssd1 vccd1 vccd1 _02621_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_109_3633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11514__C1 net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_3644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_3655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11016_ ag2.body\[598\] net1073 vssd1 vssd1 vccd1 vccd1 _05989_ sky130_fd_sc_hd__xor2_1
X_19661_ clknet_leaf_134_clk _00605_ net1307 vssd1 vssd1 vccd1 vccd1 control.body\[731\]
+ sky130_fd_sc_hd__dfrtp_1
X_16873_ ag2.body\[468\] net959 vssd1 vssd1 vccd1 vccd1 _02552_ sky130_fd_sc_hd__xor2_1
XANTENNA__14059__A1 net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_105_3519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14059__B2 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15256__B1 net50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_1044 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18612_ clknet_leaf_146_clk img_gen.tracker.next_frame\[50\] net1241 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[50\] sky130_fd_sc_hd__dfrtp_1
X_15824_ ag2.body\[266\] net205 _01643_ ag2.body\[258\] vssd1 vssd1 vccd1 vccd1 _01068_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_5_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19592_ clknet_leaf_117_clk _00536_ net1404 vssd1 vssd1 vccd1 vccd1 control.body\[806\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_99_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18543_ clknet_leaf_135_clk _00069_ net1298 vssd1 vssd1 vccd1 vccd1 img_gen.updater.commands.count\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09603__A net1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11817__B1 net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15755_ ag2.body\[333\] net211 _01635_ ag2.body\[325\] vssd1 vssd1 vccd1 vccd1 _01007_
+ sky130_fd_sc_hd__a22o_1
X_12967_ _07680_ net254 _07678_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[244\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_83_2840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15008__B1 _01552_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13282__A2 _07825_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17548__A2 net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16205__C1 _01728_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_83_2851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_2862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14706_ net983 ag2.body\[234\] vssd1 vssd1 vccd1 vccd1 _08867_ sky130_fd_sc_hd__xor2_1
X_11918_ img_gen.tracker.frame\[334\] net590 net577 vssd1 vssd1 vccd1 vccd1 _06890_
+ sky130_fd_sc_hd__o21a_1
X_18474_ net1514 net1508 vssd1 vssd1 vccd1 vccd1 _00005_ sky130_fd_sc_hd__or2_1
XANTENNA__10101__X _05074_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15686_ ag2.body\[384\] net136 _01616_ ag2.body\[376\] vssd1 vssd1 vccd1 vccd1 _00946_
+ sky130_fd_sc_hd__a22o_1
X_12898_ net245 _07647_ _07648_ net2004 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[207\]
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_64_2261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_2272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_2283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17425_ _03101_ _03102_ _03103_ _03100_ vssd1 vssd1 vccd1 vccd1 _03104_ sky130_fd_sc_hd__a211o_1
X_11849_ _06691_ _06720_ vssd1 vssd1 vccd1 vccd1 _06821_ sky130_fd_sc_hd__and2_2
X_14637_ net979 _04210_ ag2.body\[581\] net806 vssd1 vssd1 vccd1 vccd1 _08798_ sky130_fd_sc_hd__o22a_1
XANTENNA__14231__A1 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12964__A net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_2147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14231__B2 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_60_2158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14568_ _03965_ ag2.body\[353\] ag2.body\[354\] net829 _08728_ vssd1 vssd1 vccd1
+ vccd1 _08729_ sky130_fd_sc_hd__a221o_1
X_17356_ _03034_ vssd1 vssd1 vccd1 vccd1 _03035_ sky130_fd_sc_hd__inv_2
XANTENNA__16508__B1 net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12793__A1 net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16307_ net415 _01985_ _01984_ net371 vssd1 vssd1 vccd1 vccd1 _01986_ sky130_fd_sc_hd__a211o_1
X_13519_ _06821_ net309 _07618_ vssd1 vssd1 vccd1 vccd1 _07919_ sky130_fd_sc_hd__or3_1
X_17287_ ag2.body\[306\] net729 net934 _04102_ _02965_ vssd1 vssd1 vccd1 vccd1 _02966_
+ sky130_fd_sc_hd__a221o_1
X_14499_ net838 ag2.body\[257\] ag2.body\[258\] net828 _08657_ vssd1 vssd1 vccd1 vccd1
+ _08660_ sky130_fd_sc_hd__a221o_1
XFILLER_0_113_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload10 clknet_leaf_3_clk vssd1 vssd1 vccd1 vccd1 clkload10/Y sky130_fd_sc_hd__inv_6
XFILLER_0_24_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19026_ clknet_leaf_6_clk img_gen.tracker.next_frame\[464\] net1264 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[464\] sky130_fd_sc_hd__dfrtp_1
Xclkload21 clknet_leaf_11_clk vssd1 vssd1 vccd1 vccd1 clkload21/Y sky130_fd_sc_hd__clkinv_8
X_16238_ net432 _01891_ vssd1 vssd1 vccd1 vccd1 _01917_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_77_2666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload32 clknet_leaf_137_clk vssd1 vssd1 vccd1 vccd1 clkload32/Y sky130_fd_sc_hd__inv_16
XFILLER_0_67_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_2677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkload43 clknet_leaf_130_clk vssd1 vssd1 vccd1 vccd1 clkload43/Y sky130_fd_sc_hd__inv_8
Xclkload54 clknet_leaf_36_clk vssd1 vssd1 vccd1 vccd1 clkload54/Y sky130_fd_sc_hd__inv_6
XFILLER_0_80_1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload65 clknet_leaf_40_clk vssd1 vssd1 vccd1 vccd1 clkload65/Y sky130_fd_sc_hd__clkinv_8
Xclkload76 clknet_leaf_117_clk vssd1 vssd1 vccd1 vccd1 clkload76/Y sky130_fd_sc_hd__inv_12
XTAP_TAPCELL_ROW_58_2087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16169_ obsg2.obstacleArray\[14\] obsg2.obstacleArray\[15\] net426 vssd1 vssd1 vccd1
+ vccd1 _01848_ sky130_fd_sc_hd__mux2_1
Xclkload87 clknet_leaf_105_clk vssd1 vssd1 vccd1 vccd1 clkload87/Y sky130_fd_sc_hd__clkinvlp_4
XTAP_TAPCELL_ROW_58_2098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload98 clknet_leaf_96_clk vssd1 vssd1 vccd1 vccd1 clkload98/Y sky130_fd_sc_hd__clkinv_4
XANTENNA__10020__A2 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08991_ ag2.body\[88\] vssd1 vssd1 vccd1 vccd1 _04016_ sky130_fd_sc_hd__inv_2
XFILLER_0_122_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18764__CLK clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10571__A3 _05238_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19928_ clknet_leaf_51_clk _00872_ net1368 vssd1 vssd1 vccd1 vccd1 ag2.body\[470\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_76_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19243__RESET_B net1482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12204__A _06825_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09713__A2 _04427_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_4000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19859_ clknet_leaf_94_clk _00803_ net1436 vssd1 vssd1 vccd1 vccd1 ag2.body\[529\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_3_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09612_ _04574_ _04583_ _04584_ vssd1 vssd1 vccd1 vccd1 _04585_ sky130_fd_sc_hd__or3_2
XANTENNA__15515__A _05303_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15798__A1 ag2.body\[291\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12858__B net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09513__A net1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09543_ net1108 control.body\[1029\] vssd1 vssd1 vccd1 vccd1 _04516_ sky130_fd_sc_hd__or2_1
XANTENNA__11808__B1 net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout261_A net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14470__A1 net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout359_A net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14470__B2 net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_4530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09474_ _04427_ _04446_ net642 vssd1 vssd1 vccd1 vccd1 _04447_ sky130_fd_sc_hd__a21oi_2
XANTENNA__16747__B1 net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_4541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10378__B net1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10763__A_N net1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_4552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_4563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_4405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_4416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10946__X _05919_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout526_A net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1170_A net1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_1622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_1633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20634_ net1551 vssd1 vssd1 vccd1 vccd1 gpio_out[29] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_28_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16065__B net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_1371 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_24_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload4 clknet_4_9__leaf_clk vssd1 vssd1 vccd1 vccd1 clkload4/Y sky130_fd_sc_hd__clkinv_4
XTAP_TAPCELL_ROW_24_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20565_ clknet_leaf_43_clk _01424_ net1378 vssd1 vssd1 vccd1 vccd1 obsg2.randCord\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__16780__S net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17172__B1 net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10394__A net1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1056_X net1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1435_A net1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_823 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_514 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20496_ clknet_leaf_23_clk _01383_ net1360 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[132\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA_fanout895_A control.body_update.curr_length\[7\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_30_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_372 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1223_X net1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16278__A2 net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10180_ ag2.body\[423\] net1057 vssd1 vssd1 vccd1 vccd1 _05153_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_37_1448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout683_X net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15486__B1 _01605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10841__B net1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1206 net1214 vssd1 vssd1 vccd1 vccd1 net1206 sky130_fd_sc_hd__clkbuf_4
XANTENNA__17905__A _03533_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1217 net1221 vssd1 vssd1 vccd1 vccd1 net1217 sky130_fd_sc_hd__buf_4
Xfanout230 net233 vssd1 vssd1 vccd1 vccd1 net230 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12114__A net1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1228 net1238 vssd1 vssd1 vccd1 vccd1 net1228 sky130_fd_sc_hd__buf_4
Xfanout241 net242 vssd1 vssd1 vccd1 vccd1 net241 sky130_fd_sc_hd__clkbuf_4
Xfanout1239 net1243 vssd1 vssd1 vccd1 vccd1 net1239 sky130_fd_sc_hd__clkbuf_4
XANTENNA__20104__Q ag2.body\[294\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout252 net254 vssd1 vssd1 vccd1 vccd1 net252 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout850_X net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout263 net264 vssd1 vssd1 vccd1 vccd1 net263 sky130_fd_sc_hd__buf_2
XANTENNA__17624__B net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout274 net279 vssd1 vssd1 vccd1 vccd1 net274 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout948_X net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15238__B1 _01578_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout285 _07335_ vssd1 vssd1 vccd1 vccd1 net285 sky130_fd_sc_hd__clkbuf_2
XANTENNA__16435__C1 net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout296 _03552_ vssd1 vssd1 vccd1 vccd1 net296 sky130_fd_sc_hd__clkbuf_2
XANTENNA__15425__A _05686_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13870_ _08139_ _08143_ vssd1 vssd1 vccd1 vccd1 _08144_ sky130_fd_sc_hd__nor2_1
XFILLER_0_96_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15789__B2 ag2.body\[291\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16986__B1 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1040 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12147__S0 net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12768__B _07587_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12821_ net278 _07610_ _07611_ net1916 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[167\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_9_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_1359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14461__A1 net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14461__B2 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12752_ net236 _07579_ _07580_ net2089 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[129\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_55_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15540_ ag2.body\[526\] net160 _01611_ ag2.body\[518\] vssd1 vssd1 vccd1 vccd1 _00816_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__16738__B1 net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12472__B1 _06724_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10288__B net1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11703_ _06673_ _06674_ vssd1 vssd1 vccd1 vccd1 _06675_ sky130_fd_sc_hd__nor2_1
XFILLER_0_35_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15471_ ag2.body\[576\] net111 _01604_ ag2.body\[568\] vssd1 vssd1 vccd1 vccd1 _00754_
+ sky130_fd_sc_hd__a22o_1
X_12683_ net680 _07547_ vssd1 vssd1 vccd1 vccd1 _07548_ sky130_fd_sc_hd__nor2_1
XFILLER_0_127_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_3902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17210_ ag2.body\[53\] net947 vssd1 vssd1 vccd1 vccd1 _02889_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_13_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14422_ net976 _04195_ ag2.body\[532\] net814 _08575_ vssd1 vssd1 vccd1 vccd1 _08583_
+ sky130_fd_sc_hd__o221a_1
X_11634_ obsg2.obstacleArray\[39\] net631 net510 obsg2.obstacleArray\[35\] net506
+ vssd1 vssd1 vccd1 vccd1 _06607_ sky130_fd_sc_hd__o221a_1
XANTENNA__18637__CLK clknet_leaf_131_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18190_ _01703_ _03633_ _03705_ obsg2.obstacleArray\[92\] vssd1 vssd1 vccd1 vccd1
+ _03734_ sky130_fd_sc_hd__a31o_1
XFILLER_0_21_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09625__D1 _04585_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_1622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14353_ net1028 ag2.body\[405\] vssd1 vssd1 vccd1 vccd1 _08514_ sky130_fd_sc_hd__or2_1
X_17141_ ag2.body\[266\] net864 vssd1 vssd1 vccd1 vccd1 _02820_ sky130_fd_sc_hd__xor2_1
X_11565_ obsg2.obstacleArray\[79\] net631 net515 obsg2.obstacleArray\[75\] net1123
+ vssd1 vssd1 vccd1 vccd1 _06538_ sky130_fd_sc_hd__o221a_1
XANTENNA__16543__X _02222_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13304_ net671 net297 vssd1 vssd1 vccd1 vccd1 _07836_ sky130_fd_sc_hd__nor2_1
X_17072_ ag2.body\[27\] net848 vssd1 vssd1 vccd1 vccd1 _02751_ sky130_fd_sc_hd__xor2_1
X_10516_ ag2.body\[99\] net772 net1115 _04025_ _05488_ vssd1 vssd1 vccd1 vccd1 _05489_
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_0_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14284_ net821 ag2.body\[139\] ag2.body\[142\] net803 vssd1 vssd1 vccd1 vccd1 _08445_
+ sky130_fd_sc_hd__o22a_1
X_11496_ obsg2.obstacleArray\[112\] obsg2.obstacleArray\[116\] net512 vssd1 vssd1
+ vccd1 vccd1 _06469_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18787__CLK clknet_leaf_13_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16023_ _01695_ _01701_ vssd1 vssd1 vccd1 vccd1 _01702_ sky130_fd_sc_hd__nor2_1
X_13235_ _06821_ net309 vssd1 vssd1 vccd1 vccd1 _07806_ sky130_fd_sc_hd__nor2_1
XFILLER_0_123_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10447_ ag2.body\[453\] net1103 vssd1 vssd1 vccd1 vccd1 _05420_ sky130_fd_sc_hd__nand2_1
XFILLER_0_27_1130 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18258__A3 net37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14504__A net999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_2530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_1152 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13166_ net252 _07773_ _07774_ net1991 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[349\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_42_1628 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10378_ ag2.body\[110\] net1091 vssd1 vssd1 vccd1 vccd1 _05351_ sky130_fd_sc_hd__xor2_1
XANTENNA__15319__B net63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12117_ img_gen.tracker.frame\[147\] net609 net554 img_gen.tracker.frame\[150\] _07088_
+ vssd1 vssd1 vccd1 vccd1 _07089_ sky130_fd_sc_hd__a221o_1
X_17974_ obsg2.obstacleArray\[13\] _03596_ net529 vssd1 vssd1 vccd1 vccd1 _01264_
+ sky130_fd_sc_hd__o21a_1
XANTENNA__12024__A net1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13097_ net266 _07740_ _07741_ net1958 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[313\]
+ sky130_fd_sc_hd__a22o_1
X_19713_ clknet_leaf_134_clk _00657_ net1306 vssd1 vssd1 vccd1 vccd1 control.body\[687\]
+ sky130_fd_sc_hd__dfrtp_1
X_16925_ ag2.body\[373\] net949 vssd1 vssd1 vccd1 vccd1 _02604_ sky130_fd_sc_hd__xor2_1
X_12048_ img_gen.tracker.frame\[279\] net609 net593 img_gen.tracker.frame\[285\] vssd1
+ vssd1 vccd1 vccd1 _07020_ sky130_fd_sc_hd__a22o_1
XANTENNA__12959__A net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_2902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_1584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19644_ clknet_leaf_133_clk _00588_ net1309 vssd1 vssd1 vccd1 vccd1 control.body\[746\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_85_2924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16856_ ag2.body\[201\] net874 vssd1 vssd1 vccd1 vccd1 _02535_ sky130_fd_sc_hd__xor2_1
XFILLER_0_75_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_66_2323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15807_ ag2.body\[283\] net206 _01641_ ag2.body\[275\] vssd1 vssd1 vccd1 vccd1 _01053_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_66_2334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19575_ clknet_leaf_116_clk _00519_ net1385 vssd1 vssd1 vccd1 vccd1 control.body\[821\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09459__A1 net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_2345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16787_ net463 _02447_ vssd1 vssd1 vccd1 vccd1 _02466_ sky130_fd_sc_hd__or2_1
XANTENNA__19412__CLK clknet_leaf_103_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10479__A net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13999_ ag2.body\[135\] net212 _08160_ ag2.body\[127\] vssd1 vssd1 vccd1 vccd1 _00216_
+ sky130_fd_sc_hd__a22o_1
X_18526_ clknet_leaf_138_clk _00052_ net1293 vssd1 vssd1 vccd1 vccd1 img_gen.updater.commands.cmd_num\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_62_2209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15738_ ag2.body\[350\] net198 _01633_ ag2.body\[342\] vssd1 vssd1 vccd1 vccd1 _00992_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_1_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10198__B net1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18457_ _08145_ _03943_ _03944_ _03945_ vssd1 vssd1 vccd1 vccd1 _03946_ sky130_fd_sc_hd__a31o_1
X_15669_ ag2.body\[400\] net143 _01626_ ag2.body\[392\] vssd1 vssd1 vccd1 vccd1 _00930_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__10766__X _05739_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15401__B1 _01581_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17408_ ag2.body\[41\] net730 net848 _03989_ _03086_ vssd1 vssd1 vccd1 vccd1 _03087_
+ sky130_fd_sc_hd__a221o_1
X_09190_ ag2.body\[587\] vssd1 vssd1 vccd1 vccd1 _04215_ sky130_fd_sc_hd__inv_2
X_18388_ net326 _03808_ _03795_ vssd1 vssd1 vccd1 vccd1 _03878_ sky130_fd_sc_hd__o21a_1
XFILLER_0_111_1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_79_2728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_2739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12766__A1 net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17339_ _03013_ _03017_ vssd1 vssd1 vccd1 vccd1 _03018_ sky130_fd_sc_hd__nor2_1
XFILLER_0_16_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09631__A1 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_1577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkload110 clknet_leaf_88_clk vssd1 vssd1 vccd1 vccd1 clkload110/X sky130_fd_sc_hd__clkbuf_8
X_20350_ clknet_leaf_139_clk _01241_ net1289 vssd1 vssd1 vccd1 vccd1 img_gen.updater.commands.rR1.rainbowRNG\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_47_1528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload121 clknet_leaf_78_clk vssd1 vssd1 vccd1 vccd1 clkload121/Y sky130_fd_sc_hd__inv_4
XFILLER_0_15_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16901__B1 net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload132 clknet_leaf_73_clk vssd1 vssd1 vccd1 vccd1 clkload132/Y sky130_fd_sc_hd__clkinv_2
XFILLER_0_102_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_1242 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19009_ clknet_leaf_1_clk img_gen.tracker.next_frame\[447\] net1244 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[447\] sky130_fd_sc_hd__dfrtp_1
X_20281_ clknet_leaf_35_clk control.divider.next_count\[2\] net1348 vssd1 vssd1 vccd1
+ vccd1 control.divider.count\[2\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__14414__A net1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout107_A net114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15468__B1 _01603_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11741__A2 net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17725__A net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08974_ ag2.body\[65\] vssd1 vssd1 vccd1 vccd1 _03999_ sky130_fd_sc_hd__inv_2
XANTENNA__14701__X _08862_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1016_A net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_32_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold16 control.detect4.Q\[0\] vssd1 vssd1 vccd1 vccd1 net1578 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_89_Right_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_32_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold27 sound_gen.dac1.dacCount\[0\] vssd1 vssd1 vccd1 vccd1 net1589 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__17444__B net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold38 img_gen.tracker.frame\[136\] vssd1 vssd1 vccd1 vccd1 net1600 sky130_fd_sc_hd__dlygate4sd3_1
Xhold49 img_gen.tracker.frame\[369\] vssd1 vssd1 vccd1 vccd1 net1611 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_1619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09243__A net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10389__A net1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_1224 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout264_X net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_1831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1385_A net1386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09526_ net1226 control.body\[832\] vssd1 vssd1 vccd1 vccd1 _04499_ sky130_fd_sc_hd__nand2_1
XFILLER_0_52_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12875__Y _07638_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_26_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09457_ net901 _04238_ net640 _04429_ vssd1 vssd1 vccd1 vccd1 _04430_ sky130_fd_sc_hd__a31o_1
XANTENNA_fanout431_X net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1173_X net1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_98_Right_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11009__A1 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15943__A1 ag2.body\[165\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09388_ sound_gen.osc1.stayCount\[9\] _04354_ net270 vssd1 vssd1 vccd1 vccd1 _04378_
+ sky130_fd_sc_hd__o21ai_1
XANTENNA__10480__A2 _05254_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_464 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10836__B net1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_3220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_3231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20617_ net1560 vssd1 vssd1 vccd1 vccd1 gpio_oeb[29] sky130_fd_sc_hd__buf_2
XFILLER_0_30_1576 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12109__A net1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16804__A ag2.body\[68\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_683 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_3106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11350_ ag2.body\[441\] net1198 vssd1 vssd1 vccd1 vccd1 _06323_ sky130_fd_sc_hd__or2_1
X_20548_ clknet_leaf_105_clk _01413_ _00022_ vssd1 vssd1 vccd1 vccd1 sound_gen.osc1.stayCount\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_50_927 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10301_ net1046 control.body\[703\] vssd1 vssd1 vccd1 vccd1 _05274_ sky130_fd_sc_hd__xor2_1
XANTENNA_fanout898_X net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11980__A2 net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11281_ net1182 control.body\[1106\] vssd1 vssd1 vccd1 vccd1 _06254_ sky130_fd_sc_hd__xor2_1
X_20479_ clknet_leaf_39_clk _01366_ net1352 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[115\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_104_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10852__A net1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13020_ net342 _07532_ vssd1 vssd1 vccd1 vccd1 _07705_ sky130_fd_sc_hd__nor2_1
X_10232_ _05197_ _05198_ _05199_ _05204_ vssd1 vssd1 vccd1 vccd1 _05205_ sky130_fd_sc_hd__or4_1
XPHY_EDGE_ROW_5_Left_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09951__A_N net1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15459__B1 _01602_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_3024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1003 net1004 vssd1 vssd1 vccd1 vccd1 net1003 sky130_fd_sc_hd__buf_4
XANTENNA__17635__A ag2.body\[162\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_1504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_89_3035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10163_ ag2.body\[581\] net1101 vssd1 vssd1 vccd1 vccd1 _05136_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_89_3046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1014 ag2.randCord\[7\] vssd1 vssd1 vccd1 vccd1 net1014 sky130_fd_sc_hd__buf_6
XFILLER_0_101_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1025 net1026 vssd1 vssd1 vccd1 vccd1 net1025 sky130_fd_sc_hd__buf_4
XFILLER_0_41_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1036 net1037 vssd1 vssd1 vccd1 vccd1 net1036 sky130_fd_sc_hd__clkbuf_4
Xfanout1047 net1053 vssd1 vssd1 vccd1 vccd1 net1047 sky130_fd_sc_hd__buf_4
X_10094_ _05061_ _05062_ _05063_ _05066_ vssd1 vssd1 vccd1 vccd1 _05067_ sky130_fd_sc_hd__or4_1
X_14971_ control.body\[1029\] net157 net51 net2223 vssd1 vssd1 vccd1 vccd1 _00311_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12779__A net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1058 net1063 vssd1 vssd1 vccd1 vccd1 net1058 sky130_fd_sc_hd__clkbuf_4
Xfanout1069 ag2.x\[3\] vssd1 vssd1 vccd1 vccd1 net1069 sky130_fd_sc_hd__clkbuf_8
XANTENNA__12142__C1 net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16710_ _02386_ _02388_ net499 vssd1 vssd1 vccd1 vccd1 _02389_ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13922_ ag2.body\[66\] net184 _08152_ ag2.body\[58\] vssd1 vssd1 vccd1 vccd1 _00147_
+ sky130_fd_sc_hd__a22o_1
X_17690_ ag2.body\[158\] net701 net694 ag2.body\[159\] vssd1 vssd1 vccd1 vccd1 _03369_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12693__B1 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12498__B net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16641_ obsg2.obstacleArray\[55\] net450 net391 _02319_ vssd1 vssd1 vccd1 vccd1 _02320_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_18_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13853_ ag2.body\[16\] net116 _08134_ ag2.body\[8\] vssd1 vssd1 vccd1 vccd1 _00096_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_88_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10299__A _05177_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15631__B1 _01621_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12804_ net261 _07603_ _07604_ net1984 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[157\]
+ sky130_fd_sc_hd__a22o_1
X_19360_ clknet_leaf_94_clk _00304_ net1439 vssd1 vssd1 vccd1 vccd1 control.body\[1038\]
+ sky130_fd_sc_hd__dfrtp_1
X_16572_ _02249_ _02250_ net391 vssd1 vssd1 vccd1 vccd1 _02251_ sky130_fd_sc_hd__mux2_1
XANTENNA__17801__C net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10996_ ag2.body\[341\] net1115 vssd1 vssd1 vccd1 vccd1 _05969_ sky130_fd_sc_hd__xor2_1
X_13784_ img_gen.updater.commands.count\[11\] _08088_ img_gen.updater.commands.count\[12\]
+ vssd1 vssd1 vccd1 vccd1 _08093_ sky130_fd_sc_hd__a21o_1
X_18311_ net325 _03798_ vssd1 vssd1 vccd1 vccd1 _03807_ sky130_fd_sc_hd__or2_1
XANTENNA__12996__A1 net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15523_ ag2.body\[543\] net156 _01609_ ag2.body\[535\] vssd1 vssd1 vccd1 vccd1 _00801_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_123_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12735_ net258 _07570_ _07571_ net1770 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[121\]
+ sky130_fd_sc_hd__a22o_1
X_19291_ clknet_leaf_98_clk _00235_ net1446 vssd1 vssd1 vccd1 vccd1 control.body\[1097\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_112_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1070 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18242_ _03683_ net35 vssd1 vssd1 vccd1 vccd1 _03760_ sky130_fd_sc_hd__nor2_1
X_12666_ net292 _07536_ _07537_ net1967 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[86\]
+ sky130_fd_sc_hd__a22o_1
X_15454_ ag2.body\[593\] net88 _01602_ ag2.body\[585\] vssd1 vssd1 vccd1 vccd1 _00739_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__15934__B2 ag2.body\[164\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10746__B net1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_710 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12748__A1 net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14405_ net972 ag2.body\[3\] vssd1 vssd1 vccd1 vccd1 _08566_ sky130_fd_sc_hd__xor2_1
X_11617_ obsg2.obstacleArray\[54\] net631 net511 obsg2.obstacleArray\[50\] net508
+ vssd1 vssd1 vccd1 vccd1 _06590_ sky130_fd_sc_hd__o221a_1
X_18173_ net519 _03725_ vssd1 vssd1 vccd1 vccd1 _01334_ sky130_fd_sc_hd__nor2_1
X_12597_ net231 _07499_ _07500_ net2097 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[54\]
+ sky130_fd_sc_hd__a22o_1
X_15385_ net2595 net82 _01595_ net2229 vssd1 vssd1 vccd1 vccd1 _00677_ sky130_fd_sc_hd__a22o_1
XFILLER_0_37_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11956__C1 net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17124_ ag2.body\[516\] net964 vssd1 vssd1 vccd1 vccd1 _02803_ sky130_fd_sc_hd__or2_1
X_14336_ net812 ag2.body\[428\] ag2.body\[431\] net792 _08492_ vssd1 vssd1 vccd1 vccd1
+ _08497_ sky130_fd_sc_hd__o221a_1
X_11548_ _06511_ _06520_ _06503_ vssd1 vssd1 vccd1 vccd1 _06521_ sky130_fd_sc_hd__and3b_1
XANTENNA__17529__B net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_55_2002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_1296 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold508 img_gen.tracker.frame\[36\] vssd1 vssd1 vccd1 vccd1 net2070 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17055_ ag2.body\[77\] net706 net701 ag2.body\[78\] vssd1 vssd1 vccd1 vccd1 _02734_
+ sky130_fd_sc_hd__a22o_1
X_14267_ net1016 ag2.body\[14\] vssd1 vssd1 vccd1 vccd1 _08428_ sky130_fd_sc_hd__nand2_1
Xhold519 img_gen.tracker.frame\[28\] vssd1 vssd1 vccd1 vccd1 net2081 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_55_2013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11479_ ag2.body\[489\] net1208 vssd1 vssd1 vccd1 vccd1 _06452_ sky130_fd_sc_hd__xor2_1
XFILLER_0_64_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14234__A net1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13173__A1 net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16006_ net882 net850 vssd1 vssd1 vccd1 vccd1 _01685_ sky130_fd_sc_hd__and2b_1
X_13218_ net287 _07796_ _07797_ net1597 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[377\]
+ sky130_fd_sc_hd__a22o_1
X_14198_ net1042 ag2.body\[364\] vssd1 vssd1 vccd1 vccd1 _08359_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_106_1459 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10481__B net1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11723__A2 net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13149_ _07766_ net252 _07764_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[340\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17957_ net47 net296 _03582_ vssd1 vssd1 vccd1 vccd1 _03583_ sky130_fd_sc_hd__and3_1
XANTENNA__15336__Y _01590_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_68_2407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16908_ _04077_ net951 net692 ag2.body\[247\] _02583_ vssd1 vssd1 vccd1 vccd1 _02587_
+ sky130_fd_sc_hd__a221o_1
X_17888_ _08141_ _03519_ _03521_ _03522_ _03527_ vssd1 vssd1 vccd1 vccd1 _03528_ sky130_fd_sc_hd__a221o_1
XFILLER_0_79_1392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19928__CLK clknet_leaf_51_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19627_ clknet_leaf_119_clk _00571_ net1391 vssd1 vssd1 vccd1 vccd1 control.body\[761\]
+ sky130_fd_sc_hd__dfrtp_1
X_16839_ ag2.body\[97\] net735 net699 ag2.body\[102\] _02511_ vssd1 vssd1 vccd1 vccd1
+ _02518_ sky130_fd_sc_hd__o221a_1
XFILLER_0_75_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09998__A net1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19558_ clknet_leaf_115_clk _00502_ net1389 vssd1 vssd1 vccd1 vccd1 control.body\[836\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_94_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10002__A net1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09311_ _04319_ _04327_ _04329_ net272 sound_gen.osc1.count\[6\] vssd1 vssd1 vccd1
+ vccd1 _01441_ sky130_fd_sc_hd__a32o_1
XFILLER_0_48_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18509_ net1517 net1511 vssd1 vssd1 vccd1 vccd1 _00040_ sky130_fd_sc_hd__or2_1
XANTENNA__12987__A1 net233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19489_ clknet_leaf_114_clk _00433_ net1400 vssd1 vssd1 vccd1 vccd1 control.body\[911\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__18952__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10998__B1 net1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14409__A net1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10937__A ag2.body\[303\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09242_ net947 vssd1 vssd1 vccd1 vccd1 _04267_ sky130_fd_sc_hd__inv_2
XANTENNA__13313__A _07490_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10656__B net1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09173_ ag2.body\[542\] vssd1 vssd1 vccd1 vccd1 _04198_ sky130_fd_sc_hd__inv_2
XANTENNA__17127__B1 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20402_ clknet_leaf_25_clk _01289_ net1341 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[38\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_82_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11962__A2 net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20333_ clknet_leaf_21_clk _01224_ net1364 vssd1 vssd1 vccd1 vccd1 ag2.apple_cord\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__16350__A1 _01919_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1133_A net1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput17 net17 vssd1 vssd1 vccd1 vccd1 gpio_out[16] sky130_fd_sc_hd__buf_2
XANTENNA__09238__A net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput28 net28 vssd1 vssd1 vccd1 vccd1 gpio_out[3] sky130_fd_sc_hd__buf_2
XFILLER_0_25_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20264_ clknet_leaf_43_clk _01208_ net1372 vssd1 vssd1 vccd1 vccd1 control.body_update.direction\[2\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__11487__B net1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout593_A net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16638__C1 _02228_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11714__A2 net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20163__RESET_B net1480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20195_ clknet_leaf_88_clk _01139_ net1454 vssd1 vssd1 vccd1 vccd1 ag2.body\[193\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__10922__B1 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1019_X net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17174__B net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout381_X net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08957_ ag2.body\[18\] vssd1 vssd1 vccd1 vccd1 _03982_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout760_A net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout858_A net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout646_X net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14416__A1 net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15613__B1 _01620_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1378 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14416__B2 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11008__A net1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10850_ _03987_ net1196 net1147 _03989_ _05822_ vssd1 vssd1 vccd1 vccd1 _05823_ sky130_fd_sc_hd__a221o_1
XFILLER_0_6_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09509_ _04144_ net1162 _04473_ _04474_ _04481_ vssd1 vssd1 vccd1 vccd1 _04482_ sky130_fd_sc_hd__a221o_1
XFILLER_0_78_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout813_X net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10781_ net1047 control.body\[631\] vssd1 vssd1 vccd1 vccd1 _05754_ sky130_fd_sc_hd__nand2_1
X_12520_ net339 _07314_ vssd1 vssd1 vccd1 vccd1 _07457_ sky130_fd_sc_hd__or2_1
XANTENNA__09420__B net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_117_Right_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12451_ _07322_ _07354_ _07410_ vssd1 vssd1 vccd1 vccd1 _07411_ sky130_fd_sc_hd__and3_1
XFILLER_0_129_1415 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11402_ ag2.body\[571\] net1150 vssd1 vssd1 vccd1 vccd1 _06375_ sky130_fd_sc_hd__nand2_1
X_15170_ control.body\[853\] net95 _01570_ control.body\[845\] vssd1 vssd1 vccd1 vccd1
+ _00487_ sky130_fd_sc_hd__a22o_1
XFILLER_0_30_1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10205__A2 _04599_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12382_ _07218_ _07221_ _07346_ vssd1 vssd1 vccd1 vccd1 _07347_ sky130_fd_sc_hd__and3_1
XFILLER_0_34_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14121_ net1018 ag2.body\[374\] vssd1 vssd1 vccd1 vccd1 _08282_ sky130_fd_sc_hd__or2_1
XFILLER_0_104_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11333_ net1118 control.body\[660\] vssd1 vssd1 vccd1 vccd1 _06306_ sky130_fd_sc_hd__xor2_1
XANTENNA__11953__A2 net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1150 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16341__A1 net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15144__A2 net107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14054__A net1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13155__A1 net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14052_ net824 ag2.body\[186\] ag2.body\[190\] net799 vssd1 vssd1 vccd1 vccd1 _08213_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_120_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11264_ _06233_ _06234_ _06235_ _06236_ vssd1 vssd1 vccd1 vccd1 _06237_ sky130_fd_sc_hd__or4_1
XANTENNA__16629__C1 net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13003_ _07519_ _07639_ vssd1 vssd1 vccd1 vccd1 _07697_ sky130_fd_sc_hd__nor2_1
XANTENNA__11705__A2 net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10215_ _05186_ _05187_ vssd1 vssd1 vccd1 vccd1 _05188_ sky130_fd_sc_hd__nand2_1
X_18860_ clknet_leaf_18_clk img_gen.tracker.next_frame\[298\] net1320 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[298\] sky130_fd_sc_hd__dfrtp_1
X_11195_ _06164_ _06165_ _06166_ _06167_ net637 vssd1 vssd1 vccd1 vccd1 _06168_ sky130_fd_sc_hd__a221o_1
XFILLER_0_105_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17811_ net927 _03477_ _03478_ vssd1 vssd1 vccd1 vccd1 _03479_ sky130_fd_sc_hd__nand3_1
XANTENNA__16644__A2 net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10146_ _04520_ _05098_ _05103_ _05118_ vssd1 vssd1 vccd1 vccd1 _05119_ sky130_fd_sc_hd__o31a_1
XFILLER_0_118_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18791_ clknet_leaf_17_clk img_gen.tracker.next_frame\[229\] net1319 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[229\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_98_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17742_ _03075_ _03079_ _03273_ _02800_ _02692_ vssd1 vssd1 vccd1 vccd1 _03421_ sky130_fd_sc_hd__o2111a_1
X_10077_ _05036_ net479 _05026_ _05035_ vssd1 vssd1 vccd1 vccd1 _05050_ sky130_fd_sc_hd__o2bb2a_1
X_14954_ control.body\[1045\] net174 _01546_ net2437 vssd1 vssd1 vccd1 vccd1 _00295_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_76_1554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12130__A2 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13905_ ag2.body\[51\] net90 _08150_ ag2.body\[43\] vssd1 vssd1 vccd1 vccd1 _00132_
+ sky130_fd_sc_hd__a22o_1
X_17673_ ag2.body\[449\] net732 net690 ag2.body\[455\] _03351_ vssd1 vssd1 vccd1 vccd1
+ _03352_ sky130_fd_sc_hd__o221a_1
XANTENNA__14407__A1 net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16268__X _01947_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14885_ net895 _04861_ net66 vssd1 vssd1 vccd1 vccd1 _01539_ sky130_fd_sc_hd__and3_2
XANTENNA__18975__CLK clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15604__B1 _01619_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkload2_A clknet_4_4__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19412_ clknet_leaf_103_clk _00356_ net1432 vssd1 vssd1 vccd1 vccd1 control.body\[978\]
+ sky130_fd_sc_hd__dfrtp_1
X_16624_ _02301_ _02302_ net394 vssd1 vssd1 vccd1 vccd1 _02303_ sky130_fd_sc_hd__mux2_1
XANTENNA__10692__A2 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13836_ _08103_ _08129_ net1119 vssd1 vssd1 vccd1 vccd1 _00084_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19343_ clknet_leaf_100_clk net2304 net1444 vssd1 vssd1 vccd1 vccd1 control.body\[1053\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_130_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16555_ obsg2.obstacleArray\[111\] net449 net390 _02233_ vssd1 vssd1 vccd1 vccd1
+ _02234_ sky130_fd_sc_hd__o211a_1
XANTENNA__10757__A net1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13767_ net320 _08079_ vssd1 vssd1 vccd1 vccd1 _08081_ sky130_fd_sc_hd__nor2_1
X_10979_ net1119 control.body\[756\] vssd1 vssd1 vccd1 vccd1 _05952_ sky130_fd_sc_hd__xor2_1
XANTENNA__14229__A net997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12675__C _07542_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15506_ _05302_ net65 vssd1 vssd1 vccd1 vccd1 _01608_ sky130_fd_sc_hd__and2_2
XFILLER_0_84_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12718_ net258 _07562_ _07563_ net2006 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[112\]
+ sky130_fd_sc_hd__a22o_1
X_19274_ clknet_leaf_97_clk net2158 net1450 vssd1 vssd1 vccd1 vccd1 control.body\[1112\]
+ sky130_fd_sc_hd__dfrtp_1
X_16486_ _02156_ _02157_ net401 vssd1 vssd1 vccd1 vccd1 _02165_ sky130_fd_sc_hd__mux2_1
X_13698_ net923 track.highScore\[0\] track.highScore\[1\] vssd1 vssd1 vccd1 vccd1
+ _08039_ sky130_fd_sc_hd__and3_1
XFILLER_0_72_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18225_ obsg2.obstacleArray\[109\] _03751_ net520 vssd1 vssd1 vccd1 vccd1 _01360_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_116_929 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15437_ ag2.body\[610\] net83 _01600_ ag2.body\[602\] vssd1 vssd1 vccd1 vccd1 _00724_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__17109__B1 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12649_ net311 _07528_ vssd1 vssd1 vccd1 vccd1 _07529_ sky130_fd_sc_hd__and2_1
XFILLER_0_109_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13394__A1 net238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18156_ net47 _03586_ _03704_ obsg2.obstacleArray\[75\] vssd1 vssd1 vccd1 vccd1 _03717_
+ sky130_fd_sc_hd__a31o_1
X_15368_ net2563 net69 _01593_ net2244 vssd1 vssd1 vccd1 vccd1 _00662_ sky130_fd_sc_hd__a22o_1
XFILLER_0_13_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_68_Left_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17107_ ag2.body\[9\] net732 net690 ag2.body\[15\] vssd1 vssd1 vccd1 vccd1 _02786_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11944__A2 net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14319_ net825 ag2.body\[450\] ag2.body\[453\] net807 vssd1 vssd1 vccd1 vccd1 _08480_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_68_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold305 img_gen.tracker.frame\[115\] vssd1 vssd1 vccd1 vccd1 net1867 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18087_ net44 _03673_ vssd1 vssd1 vccd1 vccd1 _03674_ sky130_fd_sc_hd__nor2_1
XANTENNA__15135__A2 net107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold316 img_gen.tracker.frame\[490\] vssd1 vssd1 vccd1 vccd1 net1878 sky130_fd_sc_hd__dlygate4sd3_1
X_15299_ control.body\[743\] net76 _01585_ control.body\[735\] vssd1 vssd1 vccd1 vccd1
+ _00601_ sky130_fd_sc_hd__a22o_1
XFILLER_0_48_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold327 _04341_ vssd1 vssd1 vccd1 vccd1 net1889 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold338 img_gen.tracker.frame\[134\] vssd1 vssd1 vccd1 vccd1 net1900 sky130_fd_sc_hd__dlygate4sd3_1
X_17038_ ag2.body\[120\] net740 net734 ag2.body\[121\] vssd1 vssd1 vccd1 vccd1 _02717_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__16883__A2 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold349 img_gen.tracker.frame\[446\] vssd1 vssd1 vccd1 vccd1 net1911 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11100__B net1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09860_ ag2.body\[155\] net1163 vssd1 vssd1 vccd1 vccd1 _04833_ sky130_fd_sc_hd__xor2_1
Xfanout807 net810 vssd1 vssd1 vccd1 vccd1 net807 sky130_fd_sc_hd__buf_4
XFILLER_0_106_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout818 net819 vssd1 vssd1 vccd1 vccd1 net818 sky130_fd_sc_hd__buf_4
XFILLER_0_110_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout829 net830 vssd1 vssd1 vccd1 vccd1 net829 sky130_fd_sc_hd__buf_4
XFILLER_0_123_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16635__A2 net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09791_ net1229 control.body\[944\] vssd1 vssd1 vccd1 vccd1 _04764_ sky130_fd_sc_hd__xor2_1
X_18989_ clknet_leaf_8_clk img_gen.tracker.next_frame\[427\] net1270 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[427\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__12106__C1 _06661_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1005 control.body\[795\] vssd1 vssd1 vccd1 vccd1 net2567 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14646__A1 net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1016 control.body\[811\] vssd1 vssd1 vccd1 vccd1 net2578 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__15843__B1 _01644_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14646__B2 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1027 control.body\[638\] vssd1 vssd1 vccd1 vccd1 net2589 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13308__A net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09505__B net1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1606 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1038 control.body\[788\] vssd1 vssd1 vccd1 vccd1 net2600 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1049 control.body\[818\] vssd1 vssd1 vccd1 vccd1 net2611 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_1575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10354__A_N ag2.body\[294\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_77_Left_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_960 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17060__A2 net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout341_A net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1083_A net1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout439_A net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13043__A net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_602 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11632__A1 net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19130__CLK clknet_leaf_141_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_132_clk_X clknet_leaf_132_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09225_ control.body\[973\] vssd1 vssd1 vccd1 vccd1 _04250_ sky130_fd_sc_hd__inv_2
XFILLER_0_106_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout606_A net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1250_A net1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12882__A net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout227_X net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1348_A net1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_86_Left_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13385__A1 net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09156_ ag2.body\[500\] vssd1 vssd1 vccd1 vccd1 _04181_ sky130_fd_sc_hd__inv_2
XFILLER_0_115_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20344__RESET_B net1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_910 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09087_ ag2.body\[327\] vssd1 vssd1 vccd1 vccd1 _04112_ sky130_fd_sc_hd__inv_2
XANTENNA__09239__Y _04264_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15126__A2 net107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_110_clk clknet_4_10__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_110_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_62_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1136_X net1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18848__CLK clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20316_ clknet_leaf_44_clk obsrand1.next_randY\[2\] net1381 vssd1 vssd1 vccd1 vccd1
+ ag2.randCord\[2\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_101_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16874__A2 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11148__B1 _06109_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold850 control.body\[724\] vssd1 vssd1 vccd1 vccd1 net2412 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout975_A net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout596_X net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold861 control.body\[656\] vssd1 vssd1 vccd1 vccd1 net2423 sky130_fd_sc_hd__dlygate4sd3_1
Xhold872 _00469_ vssd1 vssd1 vccd1 vccd1 net2434 sky130_fd_sc_hd__dlygate4sd3_1
X_20247_ clknet_leaf_69_clk _01191_ net1497 vssd1 vssd1 vccd1 vccd1 ag2.body\[149\]
+ sky130_fd_sc_hd__dfrtp_2
Xhold883 _00697_ vssd1 vssd1 vccd1 vccd1 net2445 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold894 control.body\[942\] vssd1 vssd1 vccd1 vccd1 net2456 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10000_ _04969_ _04970_ _04971_ _04972_ vssd1 vssd1 vccd1 vccd1 _04973_ sky130_fd_sc_hd__a22o_1
XANTENNA__16626__A2 net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20178_ clknet_leaf_88_clk _01122_ net1461 vssd1 vssd1 vccd1 vccd1 ag2.body\[208\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_60_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout763_X net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10371__A1 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09989_ net742 _04947_ _04961_ _04937_ _04943_ vssd1 vssd1 vccd1 vccd1 _04962_ sky130_fd_sc_hd__o32a_2
XANTENNA__14637__A1 net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_95_Left_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10371__B2 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14637__B2 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17913__A _01818_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout930_X net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11951_ img_gen.tracker.frame\[97\] net619 _06921_ _06922_ vssd1 vssd1 vccd1 vccd1
+ _06923_ sky130_fd_sc_hd__o211a_1
XANTENNA__17587__B1 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16529__A _01700_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17051__A2 net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10902_ _05872_ _05873_ _05874_ vssd1 vssd1 vccd1 vccd1 _05875_ sky130_fd_sc_hd__a21o_1
X_14670_ net1009 ag2.body\[391\] vssd1 vssd1 vccd1 vccd1 _08831_ sky130_fd_sc_hd__xor2_1
X_11882_ img_gen.tracker.frame\[13\] img_gen.tracker.frame\[16\] img_gen.tracker.frame\[19\]
+ img_gen.tracker.frame\[22\] net1216 net1191 vssd1 vssd1 vccd1 vccd1 _06854_ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout42_X net42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09431__A net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13621_ control.divider.count\[7\] _07987_ net220 vssd1 vssd1 vccd1 vccd1 _07989_
+ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_120_3975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10833_ ag2.body\[309\] net1115 vssd1 vssd1 vccd1 vccd1 _05806_ sky130_fd_sc_hd__or2_1
XANTENNA__11680__B net1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_3986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_120_3997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_101_3396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16340_ _02017_ _02018_ net417 vssd1 vssd1 vccd1 vccd1 _02019_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10764_ control.body\[888\] net1227 vssd1 vssd1 vccd1 vccd1 _05737_ sky130_fd_sc_hd__and2b_1
X_13552_ ssdec1.in\[2\] _07932_ vssd1 vssd1 vccd1 vccd1 _07934_ sky130_fd_sc_hd__nand2_1
XFILLER_0_32_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16535__Y _02214_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12503_ img_gen.tracker.frame\[14\] net649 _07446_ vssd1 vssd1 vccd1 vccd1 _07447_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_66_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16271_ _01948_ _01949_ net419 vssd1 vssd1 vccd1 vccd1 _01950_ sky130_fd_sc_hd__mux2_1
X_13483_ net250 _07904_ _07905_ net1810 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[535\]
+ sky130_fd_sc_hd__a22o_1
X_10695_ _05660_ _05661_ _05665_ _05667_ vssd1 vssd1 vccd1 vccd1 _05668_ sky130_fd_sc_hd__or4b_1
XANTENNA__12792__A net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10864__X _05837_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18010_ net351 _03621_ vssd1 vssd1 vccd1 vccd1 _03622_ sky130_fd_sc_hd__nand2_1
XANTENNA__13376__A1 net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15222_ control.body\[803\] net93 _01576_ net2440 vssd1 vssd1 vccd1 vccd1 _00533_
+ sky130_fd_sc_hd__a22o_1
X_12434_ net687 _07276_ _07300_ _07395_ _07366_ vssd1 vssd1 vccd1 vccd1 net30 sky130_fd_sc_hd__a221o_1
XFILLER_0_129_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17079__B net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15153_ control.body\[870\] net106 _01568_ net2201 vssd1 vssd1 vccd1 vccd1 _00472_
+ sky130_fd_sc_hd__a22o_1
X_12365_ _07172_ _07302_ vssd1 vssd1 vccd1 vccd1 _07331_ sky130_fd_sc_hd__and2_1
XFILLER_0_129_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_101_clk clknet_4_11__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_101_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_80_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11316_ _05870_ _06276_ _06277_ _06288_ vssd1 vssd1 vccd1 vccd1 _06289_ sky130_fd_sc_hd__o31a_1
X_14104_ net840 ag2.body\[584\] ag2.body\[591\] net790 _08264_ vssd1 vssd1 vccd1 vccd1
+ _08265_ sky130_fd_sc_hd__a221o_1
X_19961_ clknet_leaf_44_clk _00905_ net1381 vssd1 vssd1 vccd1 vccd1 ag2.body\[439\]
+ sky130_fd_sc_hd__dfrtp_4
X_15084_ _04816_ net58 vssd1 vssd1 vccd1 vccd1 _01562_ sky130_fd_sc_hd__nor2_2
XANTENNA__17807__B net56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12296_ _07202_ _07228_ vssd1 vssd1 vccd1 vccd1 _07263_ sky130_fd_sc_hd__and2_1
XFILLER_0_129_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14035_ net1004 ag2.body\[496\] vssd1 vssd1 vccd1 vccd1 _08196_ sky130_fd_sc_hd__or2_1
X_18912_ clknet_leaf_142_clk img_gen.tracker.next_frame\[350\] net1258 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[350\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_120_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11247_ ag2.body\[195\] net1155 vssd1 vssd1 vccd1 vccd1 _06220_ sky130_fd_sc_hd__or2_1
X_19892_ clknet_leaf_85_clk _00836_ net1463 vssd1 vssd1 vccd1 vccd1 ag2.body\[498\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__09606__A net1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18843_ clknet_leaf_5_clk img_gen.tracker.next_frame\[281\] net1276 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[281\] sky130_fd_sc_hd__dfrtp_1
X_11178_ _06143_ _06144_ _06148_ _06150_ vssd1 vssd1 vccd1 vccd1 _06151_ sky130_fd_sc_hd__or4_1
XANTENNA__14628__A1 net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14628__B2 net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15825__B1 _01643_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10362__B2 _05334_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13128__A net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10129_ net1218 control.body\[704\] vssd1 vssd1 vccd1 vccd1 _05102_ sky130_fd_sc_hd__xor2_1
XANTENNA__17290__A2 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18774_ clknet_leaf_16_clk img_gen.tracker.next_frame\[212\] net1321 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[212\] sky130_fd_sc_hd__dfrtp_1
X_15986_ ag2.body\[2\] _08119_ vssd1 vssd1 vccd1 vccd1 _01670_ sky130_fd_sc_hd__nand2_1
XANTENNA__09504__B1 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12103__A2 net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13300__A1 net235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17725_ net496 _03403_ vssd1 vssd1 vccd1 vccd1 _03404_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_19_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17542__B net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14937_ control.body\[1062\] net173 _01544_ net2298 vssd1 vssd1 vccd1 vccd1 _00280_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_19_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14885__C net66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17656_ ag2.body\[111\] net934 vssd1 vssd1 vccd1 vccd1 _03335_ sky130_fd_sc_hd__xnor2_1
XANTENNA__19153__CLK clknet_leaf_52_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14868_ net2157 net181 _01537_ control.body\[1104\] vssd1 vssd1 vccd1 vccd1 _00218_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_72_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16607_ net396 _02285_ _02284_ net362 vssd1 vssd1 vccd1 vccd1 _02286_ sky130_fd_sc_hd__a211o_1
X_13819_ control.body_update.direction\[0\] _08110_ _08115_ vssd1 vssd1 vccd1 vccd1
+ _08116_ sky130_fd_sc_hd__o21ba_1
XANTENNA__19268__RESET_B net1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17587_ ag2.body\[58\] net725 net689 ag2.body\[63\] _03265_ vssd1 vssd1 vccd1 vccd1
+ _03266_ sky130_fd_sc_hd__o221a_1
XFILLER_0_15_1622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_1502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14799_ net1020 ag2.body\[294\] vssd1 vssd1 vccd1 vccd1 _01470_ sky130_fd_sc_hd__nand2_1
XFILLER_0_85_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19326_ clknet_leaf_103_clk net2352 net1432 vssd1 vssd1 vccd1 vccd1 control.body\[1068\]
+ sky130_fd_sc_hd__dfrtp_1
X_16538_ _01737_ _02203_ _02215_ vssd1 vssd1 vccd1 vccd1 _02217_ sky130_fd_sc_hd__o21ai_1
XANTENNA__15997__B net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19257_ clknet_leaf_74_clk _00201_ net1500 vssd1 vssd1 vccd1 vccd1 ag2.body\[120\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_72_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16469_ _02145_ _02146_ _02147_ net364 _02076_ vssd1 vssd1 vccd1 vccd1 _02148_ sky130_fd_sc_hd__a221o_1
XANTENNA__16553__A1 net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09995__B _04695_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11090__A2 net1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09010_ ag2.body\[135\] vssd1 vssd1 vccd1 vccd1 _04035_ sky130_fd_sc_hd__inv_2
X_18208_ net301 _03566_ _03703_ obsg2.obstacleArray\[101\] vssd1 vssd1 vccd1 vccd1
+ _03743_ sky130_fd_sc_hd__a31o_1
XFILLER_0_66_1008 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19188_ clknet_leaf_126_clk _00132_ net1332 vssd1 vssd1 vccd1 vccd1 ag2.body\[51\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__11378__B1 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18139_ net529 _03708_ vssd1 vssd1 vccd1 vccd1 _01317_ sky130_fd_sc_hd__and2_1
XFILLER_0_13_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold102 img_gen.tracker.frame\[486\] vssd1 vssd1 vccd1 vccd1 net1664 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_130_4282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_1355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13119__A1 net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold113 img_gen.tracker.frame\[488\] vssd1 vssd1 vccd1 vccd1 net1675 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_130_4293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold124 img_gen.tracker.frame\[327\] vssd1 vssd1 vccd1 vccd1 net1686 sky130_fd_sc_hd__dlygate4sd3_1
Xhold135 img_gen.tracker.frame\[329\] vssd1 vssd1 vccd1 vccd1 net1697 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12590__A2 net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold146 img_gen.tracker.frame\[300\] vssd1 vssd1 vccd1 vccd1 net1708 sky130_fd_sc_hd__dlygate4sd3_1
Xhold157 img_gen.tracker.frame\[255\] vssd1 vssd1 vccd1 vccd1 net1719 sky130_fd_sc_hd__dlygate4sd3_1
X_20101_ clknet_leaf_79_clk _01045_ net1489 vssd1 vssd1 vccd1 vccd1 ag2.body\[291\]
+ sky130_fd_sc_hd__dfrtp_4
Xhold168 img_gen.tracker.frame\[183\] vssd1 vssd1 vccd1 vccd1 net1730 sky130_fd_sc_hd__dlygate4sd3_1
X_09912_ ag2.body\[133\] net1116 vssd1 vssd1 vccd1 vccd1 _04885_ sky130_fd_sc_hd__xor2_1
Xhold179 img_gen.tracker.frame\[420\] vssd1 vssd1 vccd1 vccd1 net1741 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16113__S net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout604 net605 vssd1 vssd1 vccd1 vccd1 net604 sky130_fd_sc_hd__clkbuf_2
Xfanout615 net626 vssd1 vssd1 vccd1 vccd1 net615 sky130_fd_sc_hd__buf_4
Xfanout626 _06474_ vssd1 vssd1 vccd1 vccd1 net626 sky130_fd_sc_hd__clkbuf_4
XANTENNA__17805__A1 net223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20032_ clknet_leaf_66_clk _00976_ net1472 vssd1 vssd1 vccd1 vccd1 ag2.body\[366\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__09743__B1 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09516__A net1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09843_ _04550_ _04791_ net892 vssd1 vssd1 vccd1 vccd1 _04816_ sky130_fd_sc_hd__a21oi_2
Xfanout637 _04491_ vssd1 vssd1 vccd1 vccd1 net637 sky130_fd_sc_hd__clkbuf_4
Xfanout648 net654 vssd1 vssd1 vccd1 vccd1 net648 sky130_fd_sc_hd__clkbuf_2
XANTENNA__14619__A1 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout659 _04394_ vssd1 vssd1 vccd1 vccd1 net659 sky130_fd_sc_hd__buf_1
XANTENNA_fanout291_A net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14619__B2 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13038__A net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09774_ ag2.body\[232\] net1231 vssd1 vssd1 vccd1 vccd1 _04747_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_124_4097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10949__X _05922_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17569__B1 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout556_A _06651_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1298_A net1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11853__A1 net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_54_clk_A clknet_4_12__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10397__A net1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout723_A net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout344_X net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1465_A net1478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1086_X net1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11605__A1 net1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_69_clk_A clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout609_X net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13501__A net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09208_ net1071 vssd1 vssd1 vccd1 vccd1 _04233_ sky130_fd_sc_hd__inv_2
X_10480_ _04601_ _05254_ _05450_ net637 vssd1 vssd1 vccd1 vccd1 _05453_ sky130_fd_sc_hd__o211ai_1
XANTENNA__19796__CLK clknet_leaf_127_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_112_clk_A clknet_4_10__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11369__B1 _06327_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09139_ ag2.body\[463\] vssd1 vssd1 vccd1 vccd1 _04164_ sky130_fd_sc_hd__inv_2
XFILLER_0_126_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17908__A net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_1406 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12150_ img_gen.tracker.frame\[450\] net540 _07120_ _07121_ vssd1 vssd1 vccd1 vccd1
+ _07122_ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout880_X net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11101_ _06068_ _06069_ _06072_ vssd1 vssd1 vccd1 vccd1 _06074_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_102_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12081_ img_gen.tracker.frame\[312\] net629 net556 img_gen.tracker.frame\[318\] vssd1
+ vssd1 vccd1 vccd1 _07053_ sky130_fd_sc_hd__a22o_1
XANTENNA__10860__A net1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold680 control.body\[923\] vssd1 vssd1 vccd1 vccd1 net2242 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_127_clk_A clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold691 control.body\[1085\] vssd1 vssd1 vccd1 vccd1 net2253 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09734__B1 net1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11032_ _06001_ _06002_ _06003_ _06004_ _06000_ vssd1 vssd1 vccd1 vccd1 _06005_ sky130_fd_sc_hd__a221o_1
XFILLER_0_95_1204 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15807__B1 _01641_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15840_ ag2.body\[249\] net181 _01644_ ag2.body\[241\] vssd1 vssd1 vccd1 vccd1 _01083_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__19176__CLK clknet_leaf_52_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16480__B1 net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_107_3572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15771_ ag2.body\[315\] net210 _01637_ ag2.body\[307\] vssd1 vssd1 vccd1 vccd1 _01021_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_107_3583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12983_ net254 _07686_ _07687_ net1763 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[253\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__13833__A2 net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_3594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17510_ ag2.body\[590\] net937 vssd1 vssd1 vccd1 vccd1 _03189_ sky130_fd_sc_hd__xor2_1
XFILLER_0_137_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14722_ _08880_ _08881_ _08882_ vssd1 vssd1 vccd1 vccd1 _08883_ sky130_fd_sc_hd__or3_2
XANTENNA__17930__X _03562_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_103_3458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_587 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11934_ img_gen.tracker.frame\[169\] net621 net587 img_gen.tracker.frame\[178\] _06905_
+ vssd1 vssd1 vccd1 vccd1 _06906_ sky130_fd_sc_hd__o221a_1
XFILLER_0_19_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18490_ net1516 net1510 vssd1 vssd1 vccd1 vccd1 _00021_ sky130_fd_sc_hd__or2_1
XFILLER_0_24_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_3469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17441_ _03112_ _03113_ _03114_ _03119_ vssd1 vssd1 vccd1 vccd1 _03120_ sky130_fd_sc_hd__or4b_1
XFILLER_0_129_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14653_ net1032 ag2.body\[149\] vssd1 vssd1 vccd1 vccd1 _08814_ sky130_fd_sc_hd__xor2_1
XFILLER_0_86_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16783__A1 net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11865_ net577 _06833_ _06834_ _06836_ vssd1 vssd1 vccd1 vccd1 _06837_ sky130_fd_sc_hd__a22o_1
X_13604_ control.divider.count\[20\] _07949_ _07952_ _07978_ vssd1 vssd1 vccd1 vccd1
+ _07979_ sky130_fd_sc_hd__o22a_1
XFILLER_0_55_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17372_ net927 net926 _03048_ vssd1 vssd1 vccd1 vccd1 _03051_ sky130_fd_sc_hd__and3_1
X_10816_ net1061 control.body\[1095\] vssd1 vssd1 vccd1 vccd1 _05789_ sky130_fd_sc_hd__nand2_1
X_14584_ net1023 _04014_ _04015_ net1013 vssd1 vssd1 vccd1 vccd1 _08745_ sky130_fd_sc_hd__a22o_1
X_11796_ net563 _06748_ _06750_ _06751_ net472 vssd1 vssd1 vccd1 vccd1 _06768_ sky130_fd_sc_hd__a221o_1
XFILLER_0_55_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_2790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19111_ clknet_leaf_0_clk img_gen.tracker.next_frame\[549\] net1240 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[549\] sky130_fd_sc_hd__dfrtp_1
X_16323_ obsg2.obstacleArray\[66\] obsg2.obstacleArray\[67\] net410 vssd1 vssd1 vccd1
+ vccd1 _02002_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13535_ net2131 net659 _07925_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[567\]
+ sky130_fd_sc_hd__and3_1
X_10747_ ag2.body\[500\] net1138 vssd1 vssd1 vccd1 vccd1 _05720_ sky130_fd_sc_hd__xor2_1
XANTENNA__17732__B1 _03355_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14507__A net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10280__B1 _04419_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19042_ clknet_leaf_5_clk img_gen.tracker.next_frame\[480\] net1268 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[480\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__13411__A net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16254_ _01931_ _01932_ net419 vssd1 vssd1 vccd1 vccd1 _01933_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10678_ _05646_ _05648_ _05649_ _05650_ vssd1 vssd1 vccd1 vccd1 _05651_ sky130_fd_sc_hd__or4_1
X_13466_ net671 _07898_ vssd1 vssd1 vccd1 vccd1 _07899_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_11_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15205_ control.body\[820\] net95 _01574_ net2413 vssd1 vssd1 vccd1 vccd1 _00518_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_10_1585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13130__B net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12417_ net773 net1144 vssd1 vssd1 vccd1 vccd1 _07379_ sky130_fd_sc_hd__nor2_1
XANTENNA__12021__A1 net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16185_ obsg2.obstacleArray\[32\] obsg2.obstacleArray\[33\] net421 vssd1 vssd1 vccd1
+ vccd1 _01864_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13397_ net312 _07551_ net671 vssd1 vssd1 vccd1 vccd1 _07872_ sky130_fd_sc_hd__a21oi_1
XANTENNA__16299__B1 net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16838__A2 net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15136_ control.body\[887\] net107 _01566_ net2370 vssd1 vssd1 vccd1 vccd1 _00457_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_45_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12348_ net343 _07314_ vssd1 vssd1 vccd1 vccd1 _07315_ sky130_fd_sc_hd__or2_2
XANTENNA__17537__B net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16394__S0 net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11780__B1 net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19944_ clknet_leaf_46_clk _00888_ net1375 vssd1 vssd1 vccd1 vccd1 ag2.body\[454\]
+ sky130_fd_sc_hd__dfrtp_4
X_15067_ net2291 net149 _01560_ net2479 vssd1 vssd1 vccd1 vccd1 _00394_ sky130_fd_sc_hd__a22o_1
X_12279_ img_gen.updater.commands.cmd_num\[2\] _07225_ img_gen.updater.commands.cmd_num\[1\]
+ _04273_ vssd1 vssd1 vccd1 vccd1 _07249_ sky130_fd_sc_hd__a211o_1
XFILLER_0_10_259 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14018_ _08177_ _08178_ vssd1 vssd1 vccd1 vccd1 _08179_ sky130_fd_sc_hd__nand2_1
XANTENNA__11585__B net1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15057__B _01554_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19875_ clknet_leaf_95_clk _00819_ net1440 vssd1 vssd1 vccd1 vccd1 ag2.body\[513\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__17799__B1 net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18826_ clknet_leaf_4_clk img_gen.tracker.next_frame\[264\] net1262 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[264\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__17263__A2 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18757_ clknet_leaf_16_clk img_gen.tracker.next_frame\[195\] net1313 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[195\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__17272__B net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15969_ ag2.body\[140\] net212 _01658_ ag2.body\[132\] vssd1 vssd1 vccd1 vccd1 _01198_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_88_2999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19669__CLK clknet_leaf_118_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12697__A net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17708_ obsg2.obstacleArray\[131\] net451 net392 _03386_ vssd1 vssd1 vccd1 vccd1
+ _03387_ sky130_fd_sc_hd__o211a_1
X_09490_ _04459_ _04460_ _04461_ _04462_ vssd1 vssd1 vccd1 vccd1 _04463_ sky130_fd_sc_hd__or4_1
X_18688_ clknet_leaf_29_clk img_gen.tracker.next_frame\[126\] net1335 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[126\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_118_1480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17639_ ag2.body\[163\] net852 vssd1 vssd1 vccd1 vccd1 _03318_ sky130_fd_sc_hd__or2_1
XFILLER_0_91_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15577__A2 net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11518__A_N net1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19309_ clknet_leaf_99_clk _00253_ net1445 vssd1 vssd1 vccd1 vccd1 control.body\[1083\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_15_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_136_4480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20581_ clknet_leaf_107_clk _01438_ _00045_ vssd1 vssd1 vccd1 vccd1 sound_gen.osc1.count\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__17723__B1 _01743_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout137_A net139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_132_4344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_4355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_1561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_638 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13040__B net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10009__X _04982_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1046_A net1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16829__A2 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17447__B net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11771__B1 net550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15501__A2 net113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1213_A net1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout401 net403 vssd1 vssd1 vccd1 vccd1 net401 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11118__A3 _06077_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout412 _01902_ vssd1 vssd1 vccd1 vccd1 net412 sky130_fd_sc_hd__buf_2
XFILLER_0_26_1592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_54_1955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09716__B1 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout423 net425 vssd1 vssd1 vccd1 vccd1 net423 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_100_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout434 _08023_ vssd1 vssd1 vccd1 vccd1 net434 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_54_1966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_126_4159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout445 _02214_ vssd1 vssd1 vccd1 vccd1 net445 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout673_A net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout294_X net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13991__A _04697_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20015_ clknet_leaf_59_clk _00959_ net1467 vssd1 vssd1 vccd1 vccd1 ag2.body\[381\]
+ sky130_fd_sc_hd__dfrtp_4
Xfanout456 net458 vssd1 vssd1 vccd1 vccd1 net456 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_35_1376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09826_ net1180 control.body\[922\] vssd1 vssd1 vccd1 vccd1 _04799_ sky130_fd_sc_hd__nand2_1
Xfanout467 net468 vssd1 vssd1 vccd1 vccd1 net467 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_35_1387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17254__A2 net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1001_X net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout489 _02372_ vssd1 vssd1 vccd1 vccd1 net489 sky130_fd_sc_hd__buf_2
X_09757_ ag2.body\[212\] net1140 vssd1 vssd1 vccd1 vccd1 _04730_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout840_A net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout559_X net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout938_A net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17006__A2 net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1266 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09688_ _04647_ _04655_ _04660_ _04631_ _04606_ vssd1 vssd1 vccd1 vccd1 _04661_ sky130_fd_sc_hd__o32a_1
XFILLER_0_96_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11921__S1 net1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_708 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1370_X net1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout726_X net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16765__B2 obsg2.obstacleArray\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11650_ _06497_ _06562_ _06622_ _06621_ vssd1 vssd1 vccd1 vccd1 _06623_ sky130_fd_sc_hd__or4b_1
XFILLER_0_49_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout41 _03702_ vssd1 vssd1 vccd1 vccd1 net41 sky130_fd_sc_hd__buf_4
XFILLER_0_64_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10601_ net1230 control.body\[984\] vssd1 vssd1 vccd1 vccd1 _05574_ sky130_fd_sc_hd__xor2_1
Xfanout52 net55 vssd1 vssd1 vccd1 vccd1 net52 sky130_fd_sc_hd__clkbuf_8
X_11581_ _06545_ _06553_ _06497_ vssd1 vssd1 vccd1 vccd1 _06554_ sky130_fd_sc_hd__or3b_2
XANTENNA__16517__A1 net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout63 _08131_ vssd1 vssd1 vccd1 vccd1 net63 sky130_fd_sc_hd__buf_4
XFILLER_0_135_821 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10855__A net1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout74 net79 vssd1 vssd1 vccd1 vccd1 net74 sky130_fd_sc_hd__buf_2
XFILLER_0_119_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout85 net91 vssd1 vssd1 vccd1 vccd1 net85 sky130_fd_sc_hd__buf_2
XANTENNA__11303__X _06276_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13231__A net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10532_ net1133 control.body\[916\] vssd1 vssd1 vccd1 vccd1 _05505_ sky130_fd_sc_hd__or2_1
X_13320_ net249 net316 _07495_ _07841_ net1957 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[436\]
+ sky130_fd_sc_hd__a32o_1
Xfanout96 net100 vssd1 vssd1 vccd1 vccd1 net96 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_115_3830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_3841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10574__B net1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17638__A ag2.body\[163\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_3705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10463_ net1158 control.body\[1011\] vssd1 vssd1 vccd1 vccd1 _05436_ sky130_fd_sc_hd__xor2_1
X_13251_ net384 net338 vssd1 vssd1 vccd1 vccd1 _07813_ sky130_fd_sc_hd__nor2_2
XFILLER_0_134_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16542__A net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_3716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13751__A1 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12202_ _07147_ _07172_ _07173_ _06987_ _07150_ vssd1 vssd1 vccd1 vccd1 _07174_ sky130_fd_sc_hd__o221a_1
XFILLER_0_62_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13182_ net2148 net646 _07781_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[358\]
+ sky130_fd_sc_hd__and3_1
XFILLER_0_66_1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10394_ net1135 control.body\[1060\] vssd1 vssd1 vccd1 vccd1 _05367_ sky130_fd_sc_hd__or2_1
XANTENNA__11762__B1 net550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10009__C_N _04980_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11686__A net1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12133_ _07101_ _07102_ _07104_ net564 vssd1 vssd1 vccd1 vccd1 _07105_ sky130_fd_sc_hd__a22o_1
XFILLER_0_62_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17925__X _03558_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17990_ obsg2.obstacleArray\[18\] _03607_ net531 vssd1 vssd1 vccd1 vccd1 _01269_
+ sky130_fd_sc_hd__o21a_1
XANTENNA__10590__A net1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13503__A1 net250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12064_ net569 _07032_ _07035_ vssd1 vssd1 vccd1 vccd1 _07036_ sky130_fd_sc_hd__o21ai_2
X_16941_ ag2.body\[520\] net740 net692 ag2.body\[527\] _02614_ vssd1 vssd1 vccd1 vccd1
+ _02620_ sky130_fd_sc_hd__a221o_1
XFILLER_0_79_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11514__B1 net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_3634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_3645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11015_ ag2.body\[599\] net1047 vssd1 vssd1 vccd1 vccd1 _05988_ sky130_fd_sc_hd__xor2_1
XANTENNA__11973__X _06945_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_3656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19660_ clknet_leaf_134_clk _00604_ net1307 vssd1 vssd1 vccd1 vccd1 control.body\[730\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__17245__A2 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16872_ ag2.body\[469\] net946 vssd1 vssd1 vccd1 vccd1 _02551_ sky130_fd_sc_hd__xor2_1
XFILLER_0_102_1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout990 net995 vssd1 vssd1 vccd1 vccd1 net990 sky130_fd_sc_hd__buf_4
XANTENNA__18188__B net41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18611_ clknet_leaf_146_clk img_gen.tracker.next_frame\[49\] net1239 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[49\] sky130_fd_sc_hd__dfrtp_1
X_15823_ ag2.body\[265\] net205 _01643_ ag2.body\[257\] vssd1 vssd1 vccd1 vccd1 _01067_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_126_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17092__B net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19591_ clknet_leaf_117_clk _00535_ net1384 vssd1 vssd1 vccd1 vccd1 control.body\[805\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_5_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18542_ clknet_leaf_135_clk _00068_ net1298 vssd1 vssd1 vccd1 vccd1 img_gen.updater.commands.count\[11\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__13406__A net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15754_ ag2.body\[332\] net215 _01635_ ag2.body\[324\] vssd1 vssd1 vccd1 vccd1 _01006_
+ sky130_fd_sc_hd__a22o_1
X_12966_ img_gen.tracker.frame\[244\] net645 vssd1 vssd1 vccd1 vccd1 _07680_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_83_2841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_2852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14705_ net991 ag2.body\[233\] vssd1 vssd1 vccd1 vccd1 _08866_ sky130_fd_sc_hd__xor2_1
X_18473_ _04261_ net851 _03950_ _03957_ vssd1 vssd1 vccd1 vccd1 _01426_ sky130_fd_sc_hd__a22o_1
XFILLER_0_87_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_83_2863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11917_ net559 _06884_ _06887_ net471 vssd1 vssd1 vccd1 vccd1 _06889_ sky130_fd_sc_hd__a211o_1
XANTENNA__12667__D net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15685_ ag2.body\[399\] net141 _01627_ ag2.body\[391\] vssd1 vssd1 vccd1 vccd1 _00945_
+ sky130_fd_sc_hd__a22o_1
X_12897_ net680 _07647_ vssd1 vssd1 vccd1 vccd1 _07648_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_64_2262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_2273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17424_ ag2.body\[112\] net740 net934 _04027_ vssd1 vssd1 vccd1 vccd1 _03103_ sky130_fd_sc_hd__a22o_1
XFILLER_0_74_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14636_ net970 _04211_ ag2.body\[582\] net798 _08795_ vssd1 vssd1 vccd1 vccd1 _08797_
+ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_64_2284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11848_ _06810_ _06819_ net437 vssd1 vssd1 vccd1 vccd1 _06820_ sky130_fd_sc_hd__mux2_1
XANTENNA__10565__A_N net1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_60_2148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_60_2159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17355_ net927 net925 _03030_ _03031_ _03033_ vssd1 vssd1 vccd1 vccd1 _03034_ sky130_fd_sc_hd__o311a_1
XTAP_TAPCELL_ROW_16_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14567_ net839 ag2.body\[353\] ag2.body\[355\] net822 vssd1 vssd1 vccd1 vccd1 _08728_
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_126_832 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11779_ img_gen.tracker.frame\[167\] net580 net574 vssd1 vssd1 vccd1 vccd1 _06751_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_82_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16306_ obsg2.obstacleArray\[102\] obsg2.obstacleArray\[103\] net404 vssd1 vssd1
+ vccd1 vccd1 _01985_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13141__A net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13518_ net226 _07917_ _07918_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[557\]
+ sky130_fd_sc_hd__o21bai_1
XFILLER_0_42_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17286_ ag2.body\[309\] net954 vssd1 vssd1 vccd1 vccd1 _02965_ sky130_fd_sc_hd__xor2_1
X_14498_ net1030 ag2.body\[261\] vssd1 vssd1 vccd1 vccd1 _08659_ sky130_fd_sc_hd__xor2_1
X_19025_ clknet_leaf_6_clk img_gen.tracker.next_frame\[463\] net1264 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[463\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16237_ net369 _01915_ net368 _01910_ vssd1 vssd1 vccd1 vccd1 _01916_ sky130_fd_sc_hd__o211a_1
XANTENNA__15192__B1 _01573_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload11 clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 clkload11/Y sky130_fd_sc_hd__clkinvlp_4
X_13449_ net282 _07890_ _07891_ net1821 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[515\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_2_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload22 clknet_leaf_12_clk vssd1 vssd1 vccd1 vccd1 clkload22/Y sky130_fd_sc_hd__clkinv_4
XANTENNA_max_cap357_X net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_2667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkload33 clknet_leaf_138_clk vssd1 vssd1 vccd1 vccd1 clkload33/Y sky130_fd_sc_hd__inv_16
XANTENNA__12980__A net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload44 clknet_leaf_25_clk vssd1 vssd1 vccd1 vccd1 clkload44/Y sky130_fd_sc_hd__inv_6
XTAP_TAPCELL_ROW_77_2678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload55 clknet_leaf_38_clk vssd1 vssd1 vccd1 vccd1 clkload55/Y sky130_fd_sc_hd__inv_6
XFILLER_0_109_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_58_2077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload66 clknet_leaf_41_clk vssd1 vssd1 vccd1 vccd1 clkload66/Y sky130_fd_sc_hd__inv_12
X_16168_ obsg2.obstacleArray\[12\] net423 net373 _01846_ vssd1 vssd1 vccd1 vccd1 _01847_
+ sky130_fd_sc_hd__o211a_1
XANTENNA__18130__B1 net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload77 clknet_leaf_119_clk vssd1 vssd1 vccd1 vccd1 clkload77/Y sky130_fd_sc_hd__inv_6
XTAP_TAPCELL_ROW_58_2088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10556__A1 _04553_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload88 clknet_leaf_106_clk vssd1 vssd1 vccd1 vccd1 clkload88/Y sky130_fd_sc_hd__clkinv_8
XANTENNA__11753__B1 net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_2099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11596__A net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18909__CLK clknet_leaf_144_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload99 clknet_leaf_97_clk vssd1 vssd1 vccd1 vccd1 clkload99/Y sky130_fd_sc_hd__clkinvlp_4
X_15119_ _05633_ net58 vssd1 vssd1 vccd1 vccd1 _01565_ sky130_fd_sc_hd__nor2_2
X_16099_ obsg2.obstacleArray\[82\] obsg2.obstacleArray\[83\] net428 vssd1 vssd1 vccd1
+ vccd1 _01778_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08990_ ag2.body\[87\] vssd1 vssd1 vccd1 vccd1 _04015_ sky130_fd_sc_hd__inv_2
X_19927_ clknet_leaf_51_clk _00871_ net1369 vssd1 vssd1 vccd1 vccd1 ag2.body\[469\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_76_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19491__CLK clknet_leaf_113_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17236__A2 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19858_ clknet_leaf_93_clk _00802_ net1437 vssd1 vssd1 vccd1 vccd1 ag2.body\[528\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_121_4001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_1243 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09611_ _04577_ _04580_ _04581_ _04582_ vssd1 vssd1 vccd1 vccd1 _04584_ sky130_fd_sc_hd__or4_1
X_18809_ clknet_leaf_3_clk img_gen.tracker.next_frame\[247\] net1259 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[247\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__15515__B net65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19789_ clknet_leaf_128_clk _00733_ net1328 vssd1 vssd1 vccd1 vccd1 ag2.body\[603\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_78_1298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_30_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_50_Left_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09542_ net1108 control.body\[1029\] vssd1 vssd1 vccd1 vccd1 _04515_ sky130_fd_sc_hd__nand2_1
XANTENNA__19212__RESET_B net1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_4520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09473_ net917 net913 net909 vssd1 vssd1 vccd1 vccd1 _04446_ sky130_fd_sc_hd__o21a_4
XTAP_TAPCELL_ROW_138_4531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10011__Y _04984_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_4542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout254_A net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_4553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_138_4564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_4406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_4417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11490__A_N net1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_1623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20633_ net1550 vssd1 vssd1 vccd1 vccd1 gpio_out[28] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_28_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_9__f_clk clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_9__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_135_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_28_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout421_A net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14147__A net1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1163_A net1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12593__C net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_24_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload5 clknet_4_11__leaf_clk vssd1 vssd1 vccd1 vccd1 clkload5/X sky130_fd_sc_hd__clkbuf_8
X_20564_ clknet_leaf_43_clk _01423_ net1378 vssd1 vssd1 vccd1 vccd1 obsg2.randCord\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10962__X _05935_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20495_ clknet_leaf_21_clk _01382_ net1360 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[131\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_6_595 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1330_A net1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout307_X net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_3170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1049_X net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout790_A net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18589__CLK clknet_leaf_13_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout888_A net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11744__B1 net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1216_X net1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1207 net1214 vssd1 vssd1 vccd1 vccd1 net1207 sky130_fd_sc_hd__buf_2
Xfanout220 net222 vssd1 vssd1 vccd1 vccd1 net220 sky130_fd_sc_hd__clkbuf_2
Xfanout1218 net1221 vssd1 vssd1 vccd1 vccd1 net1218 sky130_fd_sc_hd__clkbuf_4
Xfanout1229 net1230 vssd1 vssd1 vccd1 vccd1 net1229 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12114__B net1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout231 net232 vssd1 vssd1 vccd1 vccd1 net231 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout676_X net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout242 net247 vssd1 vssd1 vccd1 vccd1 net242 sky130_fd_sc_hd__clkbuf_2
XANTENNA__17227__A2 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout253 net254 vssd1 vssd1 vccd1 vccd1 net253 sky130_fd_sc_hd__clkbuf_2
Xfanout264 net269 vssd1 vssd1 vccd1 vccd1 net264 sky130_fd_sc_hd__buf_2
Xfanout275 net276 vssd1 vssd1 vccd1 vccd1 net275 sky130_fd_sc_hd__clkbuf_2
Xfanout286 net288 vssd1 vssd1 vccd1 vccd1 net286 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_57_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09809_ _04740_ _04750_ _04752_ _04781_ _04739_ vssd1 vssd1 vccd1 vccd1 _04782_ sky130_fd_sc_hd__o311a_1
XANTENNA__15425__B net52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout843_X net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17921__A net48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13226__A net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12820_ net253 _07610_ _07611_ net2062 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[166\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12147__S1 net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09468__A2 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16199__C1 _01742_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12751_ net682 _07579_ vssd1 vssd1 vccd1 vccd1 _07580_ sky130_fd_sc_hd__nor2_1
XANTENNA__12472__A1 net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_81_clk clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_81_clk
+ sky130_fd_sc_hd__clkbuf_8
X_11702_ _06641_ _06644_ _06671_ vssd1 vssd1 vccd1 vccd1 _06674_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_55_1095 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15470_ _05133_ net54 vssd1 vssd1 vccd1 vccd1 _01604_ sky130_fd_sc_hd__nor2_2
X_12682_ net307 _07546_ vssd1 vssd1 vccd1 vccd1 _07547_ sky130_fd_sc_hd__nor2_1
XANTENNA__12784__B net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16256__B net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_117_3903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14421_ net984 _04194_ ag2.body\[532\] net814 _08581_ vssd1 vssd1 vccd1 vccd1 _08582_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_65_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11633_ obsg2.obstacleArray\[33\] obsg2.obstacleArray\[37\] net510 vssd1 vssd1 vccd1
+ vccd1 _06606_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_13_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09625__C1 _04570_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14057__A net1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_854 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17140_ ag2.body\[264\] net885 vssd1 vssd1 vccd1 vccd1 _02819_ sky130_fd_sc_hd__xor2_1
XANTENNA__19364__CLK clknet_leaf_102_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14352_ net1028 ag2.body\[405\] vssd1 vssd1 vccd1 vccd1 _08513_ sky130_fd_sc_hd__nand2_1
X_11564_ obsg2.obstacleArray\[78\] net631 net510 obsg2.obstacleArray\[74\] net759
+ vssd1 vssd1 vccd1 vccd1 _06537_ sky130_fd_sc_hd__o221a_1
XFILLER_0_53_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_876 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11983__B1 net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13303_ net331 _07483_ net302 vssd1 vssd1 vccd1 vccd1 _07835_ sky130_fd_sc_hd__nor3_1
X_17071_ ag2.body\[26\] net723 net928 _03985_ vssd1 vssd1 vccd1 vccd1 _02750_ sky130_fd_sc_hd__a2bb2o_1
X_10515_ ag2.body\[98\] net1187 vssd1 vssd1 vccd1 vccd1 _05488_ sky130_fd_sc_hd__xnor2_1
X_14283_ net1033 _04038_ _04040_ net1012 _08442_ vssd1 vssd1 vccd1 vccd1 _08444_ sky130_fd_sc_hd__a221o_1
X_11495_ _06463_ _06466_ vssd1 vssd1 vccd1 vccd1 _06468_ sky130_fd_sc_hd__or2_1
X_16022_ _01689_ _01694_ vssd1 vssd1 vccd1 vccd1 _01701_ sky130_fd_sc_hd__and2_1
XFILLER_0_81_1612 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10446_ _05398_ _05399_ _05405_ _05411_ _05418_ vssd1 vssd1 vccd1 vccd1 _05419_ sky130_fd_sc_hd__a32o_1
X_13234_ net283 _07426_ _07805_ net1859 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[386\]
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_72_2520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11735__B1 net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_72_2531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16123__C1 _01742_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10377_ ag2.body\[107\] net1164 vssd1 vssd1 vccd1 vccd1 _05350_ sky130_fd_sc_hd__xor2_1
X_13165_ net232 _07773_ _07774_ net1727 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[348\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_21_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12116_ img_gen.tracker.frame\[144\] net627 net593 img_gen.tracker.frame\[153\] vssd1
+ vssd1 vccd1 vccd1 _07088_ sky130_fd_sc_hd__a22o_1
X_17973_ net45 _03595_ vssd1 vssd1 vccd1 vccd1 _03596_ sky130_fd_sc_hd__nor2_1
X_13096_ net243 _07740_ _07741_ net1797 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[312\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_97_1107 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12024__B net1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16924_ ag2.body\[368\] net884 vssd1 vssd1 vccd1 vccd1 _02603_ sky130_fd_sc_hd__xor2_1
XFILLER_0_104_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19712_ clknet_leaf_135_clk _00656_ net1301 vssd1 vssd1 vccd1 vccd1 control.body\[686\]
+ sky130_fd_sc_hd__dfrtp_1
X_12047_ img_gen.tracker.frame\[255\] net610 net593 img_gen.tracker.frame\[261\] _07018_
+ vssd1 vssd1 vccd1 vccd1 _07019_ sky130_fd_sc_hd__a221o_1
XANTENNA__12160__B1 net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_2903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19643_ clknet_leaf_133_clk _00587_ net1391 vssd1 vssd1 vccd1 vccd1 control.body\[745\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11863__B net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16855_ ag2.body\[202\] net863 vssd1 vssd1 vccd1 vccd1 _02534_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_85_2914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_1596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15806_ ag2.body\[282\] net206 _01641_ ag2.body\[274\] vssd1 vssd1 vccd1 vccd1 _01052_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_66_2324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19574_ clknet_leaf_118_clk net2414 net1388 vssd1 vssd1 vccd1 vccd1 control.body\[820\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_66_2335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16786_ _02453_ _02455_ _02457_ net498 net432 vssd1 vssd1 vccd1 vccd1 _02465_ sky130_fd_sc_hd__o221a_1
XFILLER_0_1_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13998_ ag2.body\[134\] net212 _08160_ ag2.body\[126\] vssd1 vssd1 vccd1 vccd1 _00215_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__09459__A2 net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_2346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18525_ clknet_leaf_138_clk img_gen.updater.update.next\[2\] net1293 vssd1 vssd1
+ vccd1 vccd1 img_gen.updater.commands.mode\[2\] sky130_fd_sc_hd__dfrtp_2
X_15737_ ag2.body\[349\] net198 _01633_ ag2.body\[341\] vssd1 vssd1 vccd1 vccd1 _00991_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_88_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12949_ img_gen.tracker.frame\[235\] net660 vssd1 vssd1 vccd1 vccd1 _07672_ sky130_fd_sc_hd__and2_1
XFILLER_0_75_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12975__A net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_72_clk clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_72_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_14_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18456_ _04696_ _04791_ _08144_ _03845_ vssd1 vssd1 vccd1 vccd1 _03945_ sky130_fd_sc_hd__a31o_1
XFILLER_0_47_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15668_ _04472_ net67 vssd1 vssd1 vccd1 vccd1 _01626_ sky130_fd_sc_hd__and2_2
XFILLER_0_5_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17407_ _03987_ net868 net858 _03988_ vssd1 vssd1 vccd1 vccd1 _03086_ sky130_fd_sc_hd__a22o_1
X_14619_ net806 ag2.body\[61\] ag2.body\[62\] net798 _08778_ vssd1 vssd1 vccd1 vccd1
+ _08780_ sky130_fd_sc_hd__o221a_1
XANTENNA__12215__B2 net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18387_ _03805_ _03873_ _03795_ vssd1 vssd1 vccd1 vccd1 _03877_ sky130_fd_sc_hd__a21oi_1
X_15599_ ag2.body\[465\] net122 _01619_ ag2.body\[457\] vssd1 vssd1 vccd1 vccd1 _00867_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_28_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_79_2718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_79_2729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17338_ _03010_ _03015_ vssd1 vssd1 vccd1 vccd1 _03017_ sky130_fd_sc_hd__or2_1
XFILLER_0_83_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17154__B2 net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18731__CLK clknet_leaf_142_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload100 clknet_leaf_98_clk vssd1 vssd1 vccd1 vccd1 clkload100/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_126_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkload111 clknet_leaf_58_clk vssd1 vssd1 vccd1 vccd1 clkload111/Y sky130_fd_sc_hd__bufinv_16
XANTENNA__19857__CLK clknet_leaf_93_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17269_ _04083_ net951 net699 ag2.body\[254\] vssd1 vssd1 vccd1 vccd1 _02948_ sky130_fd_sc_hd__o22a_1
XANTENNA__16362__C1 net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload122 clknet_leaf_79_clk vssd1 vssd1 vccd1 vccd1 clkload122/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_113_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkload133 clknet_leaf_74_clk vssd1 vssd1 vccd1 vccd1 clkload133/Y sky130_fd_sc_hd__inv_8
X_19008_ clknet_leaf_0_clk img_gen.tracker.next_frame\[446\] net1245 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[446\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_71_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09919__B1 net1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire477_X net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20280_ clknet_leaf_35_clk net2160 net1348 vssd1 vssd1 vccd1 vccd1 control.divider.count\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18103__B1 net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10942__B net1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_127_4210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16665__B1 net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08973_ ag2.body\[63\] vssd1 vssd1 vccd1 vccd1 _03998_ sky130_fd_sc_hd__inv_2
XANTENNA__14140__A1 net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold17 img_gen.control.detect4.Q\[0\] vssd1 vssd1 vccd1 vccd1 net1579 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_32_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14140__B2 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold28 _01427_ vssd1 vssd1 vccd1 vccd1 net1590 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_32_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14729__A1_N net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16121__S net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold39 img_gen.tracker.frame\[396\] vssd1 vssd1 vccd1 vccd1 net1601 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1009_A net1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12151__B1 net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1040 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09524__A net1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15245__B net53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout469_A _06648_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_49_1810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09525_ net1051 control.body\[839\] vssd1 vssd1 vccd1 vccd1 _04498_ sky130_fd_sc_hd__or2_1
XFILLER_0_6_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12454__A1 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1280_A net1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_63_clk clknet_4_13__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_63_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout257_X net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19387__CLK clknet_leaf_102_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_26_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09456_ _04416_ _04428_ vssd1 vssd1 vccd1 vccd1 _04429_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_26_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout424_X net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout803_A net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09387_ sound_gen.osc1.stayCount\[10\] _04363_ _04356_ net270 vssd1 vssd1 vccd1 vccd1
+ _01409_ sky130_fd_sc_hd__o211a_1
XANTENNA__15943__A2 net195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_3210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1166_X net1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_95_3221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20616_ net1559 vssd1 vssd1 vccd1 vccd1 gpio_oeb[28] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_95_3232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16804__B net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12109__B net1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11965__B1 net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17696__A2 net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_91_3107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20547_ clknet_leaf_105_clk _01412_ _00021_ vssd1 vssd1 vccd1 vccd1 sound_gen.osc1.stayCount\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11013__B net1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16353__C1 net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14605__A net1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1333_X net1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10300_ net1144 control.body\[699\] vssd1 vssd1 vccd1 vccd1 _05273_ sky130_fd_sc_hd__xor2_1
XFILLER_0_50_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11280_ _06244_ _06249_ _06251_ _06252_ vssd1 vssd1 vccd1 vccd1 _06253_ sky130_fd_sc_hd__or4_2
X_20478_ clknet_leaf_39_clk _01365_ net1352 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[114\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_104_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout793_X net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10231_ _05200_ _05201_ _05202_ _05203_ vssd1 vssd1 vccd1 vccd1 _05204_ sky130_fd_sc_hd__or4_1
XANTENNA__17448__A2 net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16105__C1 net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_1375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10162_ ag2.body\[583\] net1052 vssd1 vssd1 vccd1 vccd1 _05135_ sky130_fd_sc_hd__xor2_1
XANTENNA_fanout960_X net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17635__B net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_89_3025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1004 net1005 vssd1 vssd1 vccd1 vccd1 net1004 sky130_fd_sc_hd__buf_4
XFILLER_0_98_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16120__A2 net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_3036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_3047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1015 net1019 vssd1 vssd1 vccd1 vccd1 net1015 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_101_1527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14131__A1 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1026 net1029 vssd1 vssd1 vccd1 vccd1 net1026 sky130_fd_sc_hd__clkbuf_8
Xfanout1037 net1042 vssd1 vssd1 vccd1 vccd1 net1037 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_101_1549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10093_ _05058_ _05059_ _05064_ _05065_ vssd1 vssd1 vccd1 vccd1 _05066_ sky130_fd_sc_hd__a22o_1
X_14970_ control.body\[1028\] net157 net51 control.body\[1020\] vssd1 vssd1 vccd1
+ vccd1 _00310_ sky130_fd_sc_hd__a22o_1
XFILLER_0_41_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1048 net1053 vssd1 vssd1 vccd1 vccd1 net1048 sky130_fd_sc_hd__buf_2
XANTENNA__14340__A net996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1059 net1063 vssd1 vssd1 vccd1 vccd1 net1059 sky130_fd_sc_hd__buf_4
XANTENNA__12779__B _07592_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13921_ ag2.body\[65\] net134 _08152_ ag2.body\[57\] vssd1 vssd1 vccd1 vccd1 _00146_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__15155__B net53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16640_ obsg2.obstacleArray\[54\] net444 vssd1 vssd1 vccd1 vccd1 _02319_ sky130_fd_sc_hd__or2_1
XFILLER_0_92_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13852_ _05671_ net55 vssd1 vssd1 vccd1 vccd1 _08134_ sky130_fd_sc_hd__nor2_2
XFILLER_0_134_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18466__B net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12803_ net239 _07603_ _07604_ net2050 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[156\]
+ sky130_fd_sc_hd__a22o_1
X_16571_ obsg2.obstacleArray\[126\] obsg2.obstacleArray\[127\] net444 vssd1 vssd1
+ vccd1 vccd1 _02250_ sky130_fd_sc_hd__mux2_1
X_13783_ _08091_ vssd1 vssd1 vccd1 vccd1 _08092_ sky130_fd_sc_hd__inv_2
X_10995_ ag2.body\[343\] net1067 vssd1 vssd1 vccd1 vccd1 _05968_ sky130_fd_sc_hd__xor2_1
Xclkbuf_leaf_54_clk clknet_4_12__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_54_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_85_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18310_ _03804_ _03805_ _03795_ vssd1 vssd1 vccd1 vccd1 _03806_ sky130_fd_sc_hd__o21ba_1
X_15522_ ag2.body\[542\] net156 _01609_ ag2.body\[534\] vssd1 vssd1 vccd1 vccd1 _00800_
+ sky130_fd_sc_hd__a22o_1
X_12734_ net237 _07570_ _07571_ net2076 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[120\]
+ sky130_fd_sc_hd__a22o_1
X_19290_ clknet_leaf_98_clk _00234_ net1444 vssd1 vssd1 vccd1 vccd1 control.body\[1096\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_32_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_106_Left_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18241_ obsg2.obstacleArray\[117\] _03759_ net527 vssd1 vssd1 vccd1 vccd1 _01368_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_112_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18754__CLK clknet_leaf_15_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15453_ ag2.body\[592\] net89 _01602_ net2478 vssd1 vssd1 vccd1 vccd1 _00738_ sky130_fd_sc_hd__a22o_1
X_12665_ net267 _07536_ _07537_ net1785 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[85\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_132_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14404_ net1027 net925 vssd1 vssd1 vccd1 vccd1 _08565_ sky130_fd_sc_hd__or2_1
XFILLER_0_112_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18172_ _03608_ _03705_ obsg2.obstacleArray\[83\] vssd1 vssd1 vccd1 vccd1 _03725_
+ sky130_fd_sc_hd__a21oi_1
X_11616_ obsg2.obstacleArray\[48\] obsg2.obstacleArray\[52\] net511 vssd1 vssd1 vccd1
+ vccd1 _06589_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_1420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15384_ control.body\[658\] net69 _01595_ net2226 vssd1 vssd1 vccd1 vccd1 _00676_
+ sky130_fd_sc_hd__a22o_1
X_12596_ net666 _07499_ vssd1 vssd1 vccd1 vccd1 _07500_ sky130_fd_sc_hd__nor2_1
XFILLER_0_114_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17123_ ag2.body\[517\] net952 vssd1 vssd1 vccd1 vccd1 _02802_ sky130_fd_sc_hd__or2_1
X_14335_ net818 ag2.body\[427\] ag2.body\[428\] net812 _08495_ vssd1 vssd1 vccd1 vccd1
+ _08496_ sky130_fd_sc_hd__a221o_1
XFILLER_0_107_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11547_ _06485_ _06514_ _06519_ _06497_ vssd1 vssd1 vccd1 vccd1 _06520_ sky130_fd_sc_hd__a211o_1
XANTENNA__14515__A net993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19975__RESET_B net1478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17054_ _04003_ net888 net968 _04007_ _02732_ vssd1 vssd1 vccd1 vccd1 _02733_ sky130_fd_sc_hd__a221o_1
Xhold509 img_gen.tracker.frame\[158\] vssd1 vssd1 vccd1 vccd1 net2071 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09609__A net1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_2003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14266_ net999 ag2.body\[8\] vssd1 vssd1 vccd1 vccd1 _08427_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_55_2014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11478_ _06447_ _06448_ _06449_ _06450_ vssd1 vssd1 vccd1 vccd1 _06451_ sky130_fd_sc_hd__a22o_1
XANTENNA__19904__RESET_B net1464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10762__B net1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11708__B1 net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16005_ net850 net882 vssd1 vssd1 vccd1 vccd1 _01684_ sky130_fd_sc_hd__and2b_1
XANTENNA__17439__A2 net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13217_ _07798_ net263 _07796_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[376\]
+ sky130_fd_sc_hd__mux2_1
XANTENNA__12680__D net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10429_ net1110 control.body\[1069\] vssd1 vssd1 vccd1 vccd1 _05402_ sky130_fd_sc_hd__nand2_1
XANTENNA__17826__A net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14197_ _08351_ _08352_ _08353_ _08357_ vssd1 vssd1 vccd1 vccd1 _08358_ sky130_fd_sc_hd__or4b_1
XFILLER_0_122_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_115_Left_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14070__A1_N net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13148_ img_gen.tracker.frame\[340\] net644 vssd1 vssd1 vccd1 vccd1 _07766_ sky130_fd_sc_hd__and2_1
XANTENNA__17545__B net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10931__A1 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10931__B2 net1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17956_ net345 _03581_ vssd1 vssd1 vccd1 vccd1 _03582_ sky130_fd_sc_hd__nor2_2
X_13079_ img_gen.tracker.frame\[304\] net660 vssd1 vssd1 vccd1 vccd1 _07733_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_68_2408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_1360 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16907_ _04076_ net873 net707 ag2.body\[245\] _02579_ vssd1 vssd1 vccd1 vccd1 _02586_
+ sky130_fd_sc_hd__a221o_1
XANTENNA__12684__A1 net245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17887_ _03521_ _03522_ _03524_ _03526_ vssd1 vssd1 vccd1 vccd1 _03527_ sky130_fd_sc_hd__o22a_1
XANTENNA__11109__A_N net1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19626_ clknet_leaf_123_clk net2550 net1407 vssd1 vssd1 vccd1 vccd1 control.body\[760\]
+ sky130_fd_sc_hd__dfrtp_1
X_16838_ _04023_ net873 net712 ag2.body\[100\] _02513_ vssd1 vssd1 vccd1 vccd1 _02517_
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_73_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16769_ obsg2.obstacleArray\[11\] net502 net488 obsg2.obstacleArray\[10\] vssd1 vssd1
+ vccd1 vccd1 _02448_ sky130_fd_sc_hd__a22o_1
X_19557_ clknet_leaf_116_clk _00501_ net1389 vssd1 vssd1 vccd1 vccd1 control.body\[835\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_124_Left_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_45_clk clknet_4_7__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_45_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_92_1582 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09310_ sound_gen.osc1.count\[6\] _04325_ vssd1 vssd1 vccd1 vccd1 _04329_ sky130_fd_sc_hd__or2_1
XFILLER_0_130_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18508_ net1517 net1511 vssd1 vssd1 vccd1 vccd1 _00039_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_17_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19488_ clknet_leaf_113_clk net2534 net1399 vssd1 vssd1 vccd1 vccd1 control.body\[910\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10937__B net1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09241_ net958 vssd1 vssd1 vccd1 vccd1 _04266_ sky130_fd_sc_hd__inv_2
XFILLER_0_91_817 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13313__B net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18439_ _03816_ _03913_ _03926_ _03927_ _03811_ vssd1 vssd1 vccd1 vccd1 _03928_ sky130_fd_sc_hd__a2111o_1
XANTENNA__15925__A2 net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09172_ ag2.body\[538\] vssd1 vssd1 vccd1 vccd1 _04197_ sky130_fd_sc_hd__inv_2
XANTENNA__13936__B2 ag2.body\[71\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20401_ clknet_leaf_25_clk _01288_ net1345 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[37\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__11947__B1 net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16335__C1 net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16116__S net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout217_A net218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14425__A net1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20332_ clknet_leaf_20_clk _01223_ net1364 vssd1 vssd1 vccd1 vccd1 ag2.apple_cord\[0\]
+ sky130_fd_sc_hd__dfstp_1
XPHY_EDGE_ROW_133_Left_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10672__B net1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20263_ clknet_leaf_43_clk net1629 net1372 vssd1 vssd1 vccd1 vccd1 control.body_update.direction\[1\]
+ sky130_fd_sc_hd__dfrtp_1
Xoutput18 net18 vssd1 vssd1 vccd1 vccd1 gpio_out[17] sky130_fd_sc_hd__buf_2
Xoutput29 net29 vssd1 vssd1 vccd1 vccd1 gpio_out[4] sky130_fd_sc_hd__buf_2
XANTENNA_fanout1126_A net1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20194_ clknet_leaf_54_clk _01138_ net1454 vssd1 vssd1 vccd1 vccd1 ag2.body\[192\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_25_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout586_A net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08956_ ag2.body\[17\] vssd1 vssd1 vccd1 vccd1 _03981_ sky130_fd_sc_hd__inv_2
XANTENNA__18627__CLK clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12124__B1 net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout374_X net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout753_A net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1495_A net1504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout920_A control.body_update.curr_length\[1\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__18777__CLK clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15703__B net63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout541_X net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_36_clk clknet_4_5__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_36_clk
+ sky130_fd_sc_hd__clkbuf_8
X_09508_ ag2.body\[403\] net772 net747 ag2.body\[407\] vssd1 vssd1 vccd1 vccd1 _04481_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_79_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11635__C1 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10780_ net1047 control.body\[631\] vssd1 vssd1 vccd1 vccd1 _05753_ sky130_fd_sc_hd__or2_1
XFILLER_0_78_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09843__A2 _04791_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10847__B net1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09439_ net1043 net1198 vssd1 vssd1 vccd1 vccd1 _04412_ sky130_fd_sc_hd__xor2_1
XANTENNA__15377__B1 _01594_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout806_X net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_908 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13927__A1 ag2.body\[71\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13927__B2 ag2.body\[63\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12450_ net1217 net1192 net1167 net1144 vssd1 vssd1 vccd1 vccd1 _07410_ sky130_fd_sc_hd__a31o_1
XFILLER_0_124_407 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11938__B1 net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11401_ ag2.body\[574\] net1080 vssd1 vssd1 vccd1 vccd1 _06374_ sky130_fd_sc_hd__xor2_1
XFILLER_0_90_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12381_ img_gen.updater.commands.count\[16\] _07345_ _07267_ _07227_ vssd1 vssd1
+ vccd1 vccd1 _07346_ sky130_fd_sc_hd__o211a_1
XANTENNA__10863__A _05827_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14120_ net1018 ag2.body\[374\] vssd1 vssd1 vccd1 vccd1 _08281_ sky130_fd_sc_hd__nand2_1
X_11332_ net1071 control.body\[662\] vssd1 vssd1 vccd1 vccd1 _06305_ sky130_fd_sc_hd__xor2_1
XANTENNA__11678__B net1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10582__B net1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1162 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14051_ net824 ag2.body\[186\] ag2.body\[190\] net799 _08208_ vssd1 vssd1 vccd1 vccd1
+ _08212_ sky130_fd_sc_hd__o221a_1
XANTENNA__19402__CLK clknet_leaf_103_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11263_ net773 control.body\[770\] control.body\[772\] net762 vssd1 vssd1 vccd1 vccd1
+ _06236_ sky130_fd_sc_hd__a2bb2o_1
X_13002_ net275 _07694_ _07695_ net1942 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[263\]
+ sky130_fd_sc_hd__a22o_1
X_10214_ net1179 control.body\[994\] vssd1 vssd1 vccd1 vccd1 _05187_ sky130_fd_sc_hd__xnor2_1
X_11194_ net1052 control.body\[879\] vssd1 vssd1 vccd1 vccd1 _06167_ sky130_fd_sc_hd__or2_1
XFILLER_0_24_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10374__C1 net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1213 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14104__A1 net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17810_ net925 _08124_ vssd1 vssd1 vccd1 vccd1 _03478_ sky130_fd_sc_hd__or2_1
XFILLER_0_105_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10145_ _04238_ _04759_ _05109_ _05113_ _05117_ vssd1 vssd1 vccd1 vccd1 _05118_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_20_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14104__B2 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18790_ clknet_leaf_17_clk img_gen.tracker.next_frame\[228\] net1319 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[228\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__12115__B1 net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17741_ _02816_ _02819_ _02824_ _03419_ vssd1 vssd1 vccd1 vccd1 _03420_ sky130_fd_sc_hd__o31a_1
X_10076_ _05039_ _05047_ _05048_ vssd1 vssd1 vccd1 vccd1 _05049_ sky130_fd_sc_hd__nor3_1
X_14953_ control.body\[1044\] net169 _01546_ net2085 vssd1 vssd1 vccd1 vccd1 _00294_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12666__A1 net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17054__B1 net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13904_ ag2.body\[50\] net118 _08150_ ag2.body\[42\] vssd1 vssd1 vccd1 vccd1 _00131_
+ sky130_fd_sc_hd__a22o_1
X_17672_ ag2.body\[452\] net960 vssd1 vssd1 vccd1 vccd1 _03351_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_37_1506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_1566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14884_ control.body\[1111\] net179 _01538_ net2270 vssd1 vssd1 vccd1 vccd1 _00233_
+ sky130_fd_sc_hd__a22o_1
X_16623_ obsg2.obstacleArray\[36\] obsg2.obstacleArray\[37\] net441 vssd1 vssd1 vccd1
+ vccd1 _02302_ sky130_fd_sc_hd__mux2_1
XANTENNA__16801__B1 _02057_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19411_ clknet_leaf_105_clk _00355_ net1432 vssd1 vssd1 vccd1 vccd1 control.body\[977\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_134_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13835_ net677 _08103_ vssd1 vssd1 vccd1 vccd1 _08129_ sky130_fd_sc_hd__nor2_1
XFILLER_0_114_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_27_clk clknet_4_4__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_27_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__11633__S net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_471 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16554_ obsg2.obstacleArray\[110\] net442 vssd1 vssd1 vccd1 vccd1 _02233_ sky130_fd_sc_hd__or2_1
XANTENNA__11626__C1 net1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19342_ clknet_leaf_104_clk _00286_ net1431 vssd1 vssd1 vccd1 vccd1 control.body\[1052\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_130_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13766_ _08065_ _08079_ _08080_ net320 img_gen.updater.commands.count\[6\] vssd1
+ vssd1 vccd1 vccd1 _00063_ sky130_fd_sc_hd__a32o_1
XFILLER_0_43_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10978_ net1077 control.body\[758\] vssd1 vssd1 vccd1 vccd1 _05951_ sky130_fd_sc_hd__nand2_1
XFILLER_0_84_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14229__B net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15505_ ag2.body\[559\] net113 _01607_ ag2.body\[551\] vssd1 vssd1 vccd1 vccd1 _00785_
+ sky130_fd_sc_hd__a22o_1
X_12717_ net237 _07562_ _07563_ net1998 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[111\]
+ sky130_fd_sc_hd__a22o_1
X_19273_ clknet_leaf_21_clk _00217_ net1363 vssd1 vssd1 vccd1 vccd1 ag2.appleSet sky130_fd_sc_hd__dfstp_1
XANTENNA__15368__B1 _01593_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16485_ net401 _02160_ _02159_ net366 vssd1 vssd1 vccd1 vccd1 _02164_ sky130_fd_sc_hd__a211o_1
XANTENNA__11641__A2 net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15907__A2 net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13697_ _04425_ _04637_ track.highScore\[2\] vssd1 vssd1 vccd1 vccd1 _08038_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_84_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18224_ _03666_ net40 vssd1 vssd1 vccd1 vccd1 _03751_ sky130_fd_sc_hd__nor2_1
XANTENNA__13918__A1 ag2.body\[63\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15436_ ag2.body\[609\] net83 _01600_ ag2.body\[601\] vssd1 vssd1 vccd1 vccd1 _00723_
+ sky130_fd_sc_hd__a22o_1
X_12648_ net337 _07527_ vssd1 vssd1 vccd1 vccd1 _07528_ sky130_fd_sc_hd__nor2_1
XFILLER_0_81_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18155_ net522 _03716_ vssd1 vssd1 vccd1 vccd1 _01325_ sky130_fd_sc_hd__and2_1
XFILLER_0_25_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16317__C1 _01919_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15367_ net2441 net68 _01593_ control.body\[667\] vssd1 vssd1 vccd1 vccd1 _00661_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_87_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14245__A net1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12579_ net294 _07488_ _07489_ net1885 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[47\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_68_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17106_ _03979_ net939 net930 _03980_ _02782_ vssd1 vssd1 vccd1 vccd1 _02785_ sky130_fd_sc_hd__a221o_1
XFILLER_0_41_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14318_ _08468_ _08473_ _08477_ _08478_ vssd1 vssd1 vccd1 vccd1 _08479_ sky130_fd_sc_hd__or4_2
X_18086_ net299 _03603_ vssd1 vssd1 vccd1 vccd1 _03673_ sky130_fd_sc_hd__or2_1
XFILLER_0_13_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15298_ control.body\[742\] net76 _01585_ net2512 vssd1 vssd1 vccd1 vccd1 _00600_
+ sky130_fd_sc_hd__a22o_1
Xhold306 img_gen.tracker.frame\[467\] vssd1 vssd1 vccd1 vccd1 net1868 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10492__B net1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold317 img_gen.tracker.frame\[137\] vssd1 vssd1 vccd1 vccd1 net1879 sky130_fd_sc_hd__dlygate4sd3_1
Xhold328 img_gen.tracker.frame\[81\] vssd1 vssd1 vccd1 vccd1 net1890 sky130_fd_sc_hd__dlygate4sd3_1
X_17037_ ag2.body\[124\] net713 net934 _04032_ _02714_ vssd1 vssd1 vccd1 vccd1 _02716_
+ sky130_fd_sc_hd__o221a_1
Xhold339 img_gen.tracker.frame\[301\] vssd1 vssd1 vccd1 vccd1 net1901 sky130_fd_sc_hd__dlygate4sd3_1
X_14249_ net837 ag2.body\[537\] ag2.body\[538\] net828 _08407_ vssd1 vssd1 vccd1 vccd1
+ _08410_ sky130_fd_sc_hd__a221o_1
XFILLER_0_7_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17394__A2_N net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout808 net809 vssd1 vssd1 vccd1 vccd1 net808 sky130_fd_sc_hd__buf_4
XFILLER_0_0_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17275__B net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout819 _03968_ vssd1 vssd1 vccd1 vccd1 net819 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_68_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16096__A1 net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09790_ net1133 control.body\[948\] vssd1 vssd1 vccd1 vccd1 _04763_ sky130_fd_sc_hd__xor2_1
XFILLER_0_20_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18988_ clknet_leaf_9_clk img_gen.tracker.next_frame\[426\] net1271 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[426\] sky130_fd_sc_hd__dfrtp_1
Xhold1006 control.body\[717\] vssd1 vssd1 vccd1 vccd1 net2568 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1017 control.body\[966\] vssd1 vssd1 vccd1 vccd1 net2579 sky130_fd_sc_hd__dlygate4sd3_1
X_17939_ net539 net460 net488 vssd1 vssd1 vccd1 vccd1 _03569_ sky130_fd_sc_hd__nand3_1
Xhold1028 control.body\[656\] vssd1 vssd1 vccd1 vccd1 net2590 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13308__B net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13854__B1 _08134_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1039 control.body\[663\] vssd1 vssd1 vccd1 vccd1 net2601 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_119_1618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1390 net1392 vssd1 vssd1 vccd1 vccd1 net1390 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_108_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09802__A net1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19609_ clknet_leaf_119_clk net2373 net1392 vssd1 vssd1 vccd1 vccd1 control.body\[791\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_5_Right_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11880__A2 net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_18_clk clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_18_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__11617__C1 net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_1494 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11093__B1 _06028_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13043__B _07546_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15359__B1 _01592_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout334_A _07423_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1076_A net1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09224_ control.body\[969\] vssd1 vssd1 vccd1 vccd1 _04249_ sky130_fd_sc_hd__inv_2
XFILLER_0_31_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09155_ ag2.body\[497\] vssd1 vssd1 vccd1 vccd1 _04180_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_1069 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout501_A _01708_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1243_A net1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14155__A net1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09086_ ag2.body\[324\] vssd1 vssd1 vccd1 vccd1 _04111_ sky130_fd_sc_hd__inv_2
XFILLER_0_71_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20315_ clknet_leaf_44_clk obsrand1.next_randY\[1\] net1381 vssd1 vssd1 vccd1 vccd1
+ ag2.randCord\[1\] sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_9_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14334__B2 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1031_X net1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1410_A net1415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold840 control.body\[814\] vssd1 vssd1 vccd1 vccd1 net2402 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1129_X net1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold851 control.body\[812\] vssd1 vssd1 vccd1 vccd1 net2413 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1508_A net9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold862 control.body\[636\] vssd1 vssd1 vccd1 vccd1 net2424 sky130_fd_sc_hd__dlygate4sd3_1
X_20246_ clknet_leaf_69_clk _01190_ net1497 vssd1 vssd1 vccd1 vccd1 ag2.body\[148\]
+ sky130_fd_sc_hd__dfrtp_4
Xhold873 control.body\[841\] vssd1 vssd1 vccd1 vccd1 net2435 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold884 control.body\[1068\] vssd1 vssd1 vccd1 vccd1 net2446 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__17185__B net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout491_X net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout870_A net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold895 control.body\[888\] vssd1 vssd1 vccd1 vccd1 net2457 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout589_X net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17753__X _03432_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20177_ clknet_leaf_82_clk _01121_ net1479 vssd1 vssd1 vccd1 vccd1 ag2.body\[223\]
+ sky130_fd_sc_hd__dfrtp_4
X_09988_ _04950_ _04953_ _04955_ _04960_ vssd1 vssd1 vccd1 vccd1 _04961_ sky130_fd_sc_hd__or4_2
XFILLER_0_102_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08939_ net1044 vssd1 vssd1 vccd1 vccd1 _03964_ sky130_fd_sc_hd__inv_2
XANTENNA__12122__B net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout756_X net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11950_ img_gen.tracker.frame\[100\] net601 net585 img_gen.tracker.frame\[106\] vssd1
+ vssd1 vccd1 vccd1 _06922_ sky130_fd_sc_hd__o22a_1
XFILLER_0_98_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17587__A1 ag2.body\[58\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17587__B2 ag2.body\[63\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10901_ net1218 control.body\[672\] vssd1 vssd1 vccd1 vccd1 _05874_ sky130_fd_sc_hd__xor2_1
XANTENNA__15598__B1 _01619_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11961__B net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1442 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout923_X net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11871__A2 net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11881_ _06851_ _06852_ vssd1 vssd1 vccd1 vccd1 _06853_ sky130_fd_sc_hd__nand2_1
X_13620_ _07987_ _07988_ vssd1 vssd1 vccd1 vccd1 control.divider.next_count\[6\] sky130_fd_sc_hd__nor2_1
XANTENNA__11608__C1 net1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_3976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09431__B net1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10832_ ag2.body\[307\] net1165 vssd1 vssd1 vccd1 vccd1 _05805_ sky130_fd_sc_hd__xor2_1
XFILLER_0_71_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_120_3987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout35_X net35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10577__B net1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_3998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_3397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13551_ ssdec1.in\[1\] ssdec1.in\[0\] vssd1 vssd1 vccd1 vccd1 _07933_ sky130_fd_sc_hd__or2_1
X_10763_ net1058 control.body\[895\] vssd1 vssd1 vccd1 vccd1 _05736_ sky130_fd_sc_hd__and2b_1
XFILLER_0_13_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12502_ net2016 net650 _07446_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[13\]
+ sky130_fd_sc_hd__and3_1
X_16270_ obsg2.obstacleArray\[28\] obsg2.obstacleArray\[29\] net411 vssd1 vssd1 vccd1
+ vccd1 _01949_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13482_ net230 _07904_ _07905_ net1707 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[534\]
+ sky130_fd_sc_hd__a22o_1
X_10694_ ag2.body\[144\] net788 net1113 _04043_ _05666_ vssd1 vssd1 vccd1 vccd1 _05667_
+ sky130_fd_sc_hd__o221a_1
XANTENNA__16562__A2 net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_1213 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15221_ net2593 net93 _01576_ control.body\[794\] vssd1 vssd1 vccd1 vccd1 _00532_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_30_1171 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14573__A1 net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12433_ img_gen.updater.commands.rR1.rainbowRNG\[13\] _07319_ _07338_ _07378_ _07394_
+ vssd1 vssd1 vccd1 vccd1 _07395_ sky130_fd_sc_hd__a221o_1
XANTENNA__14573__B2 net1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10593__A net1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15152_ control.body\[869\] net98 _01568_ control.body\[861\] vssd1 vssd1 vccd1 vccd1
+ _00471_ sky130_fd_sc_hd__a22o_1
X_12364_ _07264_ _07274_ _07329_ _07266_ vssd1 vssd1 vccd1 vccd1 _07330_ sky130_fd_sc_hd__a211o_1
XANTENNA__16314__A2 net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_922 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_484 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14103_ net987 _04213_ _04217_ net1006 vssd1 vssd1 vccd1 vccd1 _08264_ sky130_fd_sc_hd__a22o_1
XANTENNA__11201__B net1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11315_ _06282_ _06287_ _04985_ vssd1 vssd1 vccd1 vccd1 _06288_ sky130_fd_sc_hd__or3b_4
X_19960_ clknet_leaf_62_clk _00904_ net1382 vssd1 vssd1 vccd1 vccd1 ag2.body\[438\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__14325__B2 net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15083_ net2648 net147 _01561_ net2330 vssd1 vssd1 vccd1 vccd1 _00409_ sky130_fd_sc_hd__a22o_1
X_12295_ _04392_ _07257_ _07232_ vssd1 vssd1 vccd1 vccd1 img_gen.updater.update.next\[2\]
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_10_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14034_ net1031 ag2.body\[501\] vssd1 vssd1 vccd1 vccd1 _08195_ sky130_fd_sc_hd__xor2_1
X_18911_ clknet_leaf_142_clk img_gen.tracker.next_frame\[349\] net1258 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[349\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_31_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09446__X _04419_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17095__B net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11246_ ag2.body\[195\] net1155 vssd1 vssd1 vccd1 vccd1 _06219_ sky130_fd_sc_hd__nand2_1
XFILLER_0_129_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19891_ clknet_leaf_85_clk _00835_ net1462 vssd1 vssd1 vccd1 vccd1 ag2.body\[497\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__20054__RESET_B net1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18842_ clknet_leaf_4_clk img_gen.tracker.next_frame\[280\] net1277 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[280\] sky130_fd_sc_hd__dfrtp_1
X_11177_ _06145_ _06146_ _06147_ _06149_ vssd1 vssd1 vccd1 vccd1 _06150_ sky130_fd_sc_hd__or4_1
XFILLER_0_98_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10128_ net1170 control.body\[706\] vssd1 vssd1 vccd1 vccd1 _05101_ sky130_fd_sc_hd__xor2_1
XANTENNA__12568__B_N _07483_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15985_ _03967_ _08120_ vssd1 vssd1 vccd1 vccd1 _01669_ sky130_fd_sc_hd__nor2_1
X_18773_ clknet_leaf_16_clk img_gen.tracker.next_frame\[211\] net1315 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[211\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__17027__B1 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17724_ obsg2.obstacleArray\[128\] obsg2.obstacleArray\[129\] obsg2.obstacleArray\[130\]
+ obsg2.obstacleArray\[131\] net958 net538 vssd1 vssd1 vccd1 vccd1 _03403_ sky130_fd_sc_hd__mux4_1
X_10059_ _04173_ net1233 net1155 _04175_ _05031_ vssd1 vssd1 vccd1 vccd1 _05032_ sky130_fd_sc_hd__a221o_1
X_14936_ control.body\[1061\] net167 _01544_ net2167 vssd1 vssd1 vccd1 vccd1 _00279_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_19_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18000__A net45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09622__A net1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17655_ ag2.body\[105\] net876 vssd1 vssd1 vccd1 vccd1 _03334_ sky130_fd_sc_hd__xor2_1
XANTENNA__11464__A2_N net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14867_ _04947_ net51 vssd1 vssd1 vccd1 vccd1 _01537_ sky130_fd_sc_hd__and2b_2
XANTENNA__16786__C1 net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11862__A2 net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13818_ _08112_ _08114_ _08113_ _08111_ vssd1 vssd1 vccd1 vccd1 _08115_ sky130_fd_sc_hd__or4b_1
X_16606_ obsg2.obstacleArray\[80\] obsg2.obstacleArray\[81\] net447 vssd1 vssd1 vccd1
+ vccd1 _02285_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_1601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17586_ ag2.body\[60\] net962 vssd1 vssd1 vccd1 vccd1 _03265_ sky130_fd_sc_hd__xnor2_1
XANTENNA__13064__A1 net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14798_ net1042 ag2.body\[292\] vssd1 vssd1 vccd1 vccd1 _01469_ sky130_fd_sc_hd__xor2_1
XFILLER_0_97_290 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10487__B net1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16537_ _01737_ _02203_ _02215_ vssd1 vssd1 vccd1 vccd1 _02216_ sky130_fd_sc_hd__o21a_1
XANTENNA__11075__B1 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19325_ clknet_leaf_100_clk net2320 net1445 vssd1 vssd1 vccd1 vccd1 control.body\[1067\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13749_ img_gen.updater.commands.count\[2\] img_gen.updater.commands.count\[1\] img_gen.updater.commands.count\[0\]
+ vssd1 vssd1 vccd1 vccd1 _08068_ sky130_fd_sc_hd__and3_1
XANTENNA__17735__D1 _02652_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16468_ obsg2.obstacleArray\[60\] obsg2.obstacleArray\[61\] obsg2.obstacleArray\[62\]
+ obsg2.obstacleArray\[63\] net454 net397 vssd1 vssd1 vccd1 vccd1 _02147_ sky130_fd_sc_hd__mux4_1
X_19256_ clknet_leaf_75_clk _00200_ net1484 vssd1 vssd1 vccd1 vccd1 ag2.body\[119\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__20425__CLK clknet_leaf_37_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18207_ obsg2.obstacleArray\[100\] _03742_ net522 vssd1 vssd1 vccd1 vccd1 _01351_
+ sky130_fd_sc_hd__o21a_1
X_15419_ control.body\[626\] net81 _01598_ ag2.body\[618\] vssd1 vssd1 vccd1 vccd1
+ _00708_ sky130_fd_sc_hd__a22o_1
X_19187_ clknet_leaf_53_clk _00131_ net1365 vssd1 vssd1 vccd1 vccd1 ag2.body\[50\]
+ sky130_fd_sc_hd__dfrtp_4
X_16399_ obsg2.obstacleArray\[104\] obsg2.obstacleArray\[105\] net454 vssd1 vssd1
+ vccd1 vccd1 _02078_ sky130_fd_sc_hd__mux2_1
XANTENNA__19237__RESET_B net1480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11378__A1 _04427_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18138_ net48 _03554_ _03704_ obsg2.obstacleArray\[66\] vssd1 vssd1 vccd1 vccd1 _03708_
+ sky130_fd_sc_hd__a31o_1
XANTENNA__19598__CLK clknet_leaf_118_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_218 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold103 img_gen.tracker.frame\[397\] vssd1 vssd1 vccd1 vccd1 net1665 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_130_4283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_1476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16902__B net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_130_4294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14316__A1 net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold114 img_gen.tracker.frame\[73\] vssd1 vssd1 vccd1 vccd1 net1676 sky130_fd_sc_hd__dlygate4sd3_1
X_18069_ net300 _03586_ vssd1 vssd1 vccd1 vccd1 _03662_ sky130_fd_sc_hd__nand2_1
XANTENNA__14316__B2 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold125 img_gen.tracker.frame\[309\] vssd1 vssd1 vccd1 vccd1 net1687 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09991__A1 net1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09991__B2 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_7_clk clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_7_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__10008__A net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold136 img_gen.tracker.frame\[123\] vssd1 vssd1 vccd1 vccd1 net1698 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14703__A net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold147 img_gen.tracker.frame\[521\] vssd1 vssd1 vccd1 vccd1 net1709 sky130_fd_sc_hd__dlygate4sd3_1
X_20100_ clknet_leaf_79_clk _01044_ net1489 vssd1 vssd1 vccd1 vccd1 ag2.body\[290\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_22_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold158 img_gen.tracker.frame\[418\] vssd1 vssd1 vccd1 vccd1 net1720 sky130_fd_sc_hd__dlygate4sd3_1
X_09911_ ag2.body\[128\] net1235 vssd1 vssd1 vccd1 vccd1 _04884_ sky130_fd_sc_hd__xor2_1
Xhold169 img_gen.tracker.frame\[9\] vssd1 vssd1 vccd1 vccd1 net1731 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12878__A1 net245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10950__B net1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout605 net608 vssd1 vssd1 vccd1 vccd1 net605 sky130_fd_sc_hd__clkbuf_4
X_20031_ clknet_leaf_66_clk _00975_ net1473 vssd1 vssd1 vccd1 vccd1 ag2.body\[365\]
+ sky130_fd_sc_hd__dfrtp_4
Xfanout616 net617 vssd1 vssd1 vccd1 vccd1 net616 sky130_fd_sc_hd__clkbuf_4
XANTENNA__17266__B1 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout627 net628 vssd1 vssd1 vccd1 vccd1 net627 sky130_fd_sc_hd__clkbuf_4
X_09842_ _04811_ _04812_ _04813_ _04814_ _04810_ vssd1 vssd1 vccd1 vccd1 _04815_ sky130_fd_sc_hd__a221o_1
Xfanout638 _04470_ vssd1 vssd1 vccd1 vccd1 net638 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_123_1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout649 net651 vssd1 vssd1 vccd1 vccd1 net649 sky130_fd_sc_hd__clkbuf_2
XANTENNA__14619__A2 ag2.body\[61\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09773_ ag2.body\[239\] net1061 vssd1 vssd1 vccd1 vccd1 _04746_ sky130_fd_sc_hd__or2_1
XFILLER_0_119_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout284_A net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17018__B1 net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_4098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_1403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_1448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_1_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18230__A2 _03539_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1193_A net1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_920 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout549_A net550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13054__A net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13055__A1 net246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout716_A _04265_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout337_X net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1458_A net1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1079_X net1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18815__CLK clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10684__Y _05657_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_989 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_466 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09207_ net1095 vssd1 vssd1 vccd1 vccd1 _04232_ sky130_fd_sc_hd__clkinv_4
XANTENNA__14555__A1 net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14555__B2 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_1278 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout504_X net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_488 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11369__A1 _06331_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11369__B2 _06314_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11302__A net1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09138_ ag2.body\[462\] vssd1 vssd1 vccd1 vccd1 _04163_ sky130_fd_sc_hd__inv_2
XANTENNA__12030__A2 net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17908__B _03533_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18965__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11021__B net1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09982__A1 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_113_3780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09982__B2 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09069_ ag2.body\[275\] vssd1 vssd1 vccd1 vccd1 _04094_ sky130_fd_sc_hd__inv_2
XANTENNA__14613__A net996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11100_ ag2.body\[428\] net1127 vssd1 vssd1 vccd1 vccd1 _06073_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_103_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12080_ net473 _07050_ _07051_ vssd1 vssd1 vccd1 vccd1 _07052_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout873_X net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold670 control.body\[1057\] vssd1 vssd1 vccd1 vccd1 net2232 sky130_fd_sc_hd__dlygate4sd3_1
Xhold681 control.body\[769\] vssd1 vssd1 vccd1 vccd1 net2243 sky130_fd_sc_hd__dlygate4sd3_1
Xhold692 control.body\[868\] vssd1 vssd1 vccd1 vccd1 net2254 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__17257__B1 net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11031_ net1135 control.body\[1044\] vssd1 vssd1 vccd1 vccd1 _06004_ sky130_fd_sc_hd__or2_1
X_20229_ clknet_leaf_66_clk _01173_ net1476 vssd1 vssd1 vccd1 vccd1 ag2.body\[163\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_102_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_95_1216 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15770_ ag2.body\[314\] net209 _01637_ ag2.body\[306\] vssd1 vssd1 vccd1 vccd1 _01020_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__09713__Y _04686_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_107_3573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12097__A2 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12982_ net232 _07686_ _07687_ net1913 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[252\]
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_107_3584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14721_ _08876_ _08877_ _08878_ _08879_ _08874_ vssd1 vssd1 vccd1 vccd1 _08882_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_107_3595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11933_ img_gen.tracker.frame\[175\] net548 vssd1 vssd1 vccd1 vccd1 _06905_ sky130_fd_sc_hd__or2_1
XFILLER_0_38_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11844__A2 net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_103_3459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10588__A net1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17440_ _03116_ _03117_ _03118_ vssd1 vssd1 vccd1 vccd1 _03119_ sky130_fd_sc_hd__and3_1
XFILLER_0_73_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14652_ net829 ag2.body\[146\] ag2.body\[150\] net802 _08812_ vssd1 vssd1 vccd1 vccd1
+ _08813_ sky130_fd_sc_hd__a221o_1
XFILLER_0_38_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11864_ img_gen.tracker.frame\[196\] net607 net552 img_gen.tracker.frame\[199\] _06835_
+ vssd1 vssd1 vccd1 vccd1 _06836_ sky130_fd_sc_hd__o221a_1
X_13603_ control.divider.count\[19\] _07950_ _07974_ _07977_ vssd1 vssd1 vccd1 vccd1
+ _07978_ sky130_fd_sc_hd__a22o_1
XFILLER_0_28_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17371_ _03019_ _03023_ _03048_ vssd1 vssd1 vccd1 vccd1 _03050_ sky130_fd_sc_hd__and3b_1
XFILLER_0_95_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10815_ net1061 control.body\[1095\] vssd1 vssd1 vccd1 vccd1 _05788_ sky130_fd_sc_hd__or2_1
XANTENNA__14794__A1 net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14583_ net829 ag2.body\[82\] vssd1 vssd1 vccd1 vccd1 _08744_ sky130_fd_sc_hd__nor2_1
XFILLER_0_89_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_2780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11795_ net574 _06753_ _06756_ net467 vssd1 vssd1 vccd1 vccd1 _06767_ sky130_fd_sc_hd__a211o_1
XANTENNA__10100__B net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14794__B2 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_2791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16322_ obsg2.obstacleArray\[64\] obsg2.obstacleArray\[65\] net410 vssd1 vssd1 vccd1
+ vccd1 _02001_ sky130_fd_sc_hd__mux2_1
X_19110_ clknet_leaf_0_clk img_gen.tracker.next_frame\[548\] net1245 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[548\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_94_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13534_ _07627_ _07807_ vssd1 vssd1 vccd1 vccd1 _07925_ sky130_fd_sc_hd__or2_1
X_10746_ ag2.body\[498\] net1184 vssd1 vssd1 vccd1 vccd1 _05719_ sky130_fd_sc_hd__xor2_1
XFILLER_0_40_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1592 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19041_ clknet_leaf_6_clk img_gen.tracker.next_frame\[479\] net1267 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[479\] sky130_fd_sc_hd__dfrtp_1
X_16253_ obsg2.obstacleArray\[60\] obsg2.obstacleArray\[61\] net407 vssd1 vssd1 vccd1
+ vccd1 _01932_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13465_ net338 _07486_ net331 net313 vssd1 vssd1 vccd1 vccd1 _07898_ sky130_fd_sc_hd__and4bb_1
X_10677_ ag2.body\[345\] net1211 vssd1 vssd1 vccd1 vccd1 _05650_ sky130_fd_sc_hd__xor2_1
XFILLER_0_10_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_11_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11212__A net1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15204_ control.body\[819\] net92 _01574_ net2466 vssd1 vssd1 vccd1 vccd1 _00517_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_63_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12416_ img_gen.updater.commands.rR1.rainbowRNG\[5\] net248 _07377_ vssd1 vssd1 vccd1
+ vccd1 _07378_ sky130_fd_sc_hd__a21o_1
XFILLER_0_51_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16184_ obsg2.obstacleArray\[34\] obsg2.obstacleArray\[35\] net421 vssd1 vssd1 vccd1
+ vccd1 _01863_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_73_clk_X clknet_leaf_73_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13396_ net283 _07870_ _07871_ net2011 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[482\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_112_218 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16299__A1 net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20235__RESET_B net1499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15135_ control.body\[886\] net107 _01566_ net2316 vssd1 vssd1 vccd1 vccd1 _00456_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_23_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12347_ net387 _07313_ vssd1 vssd1 vccd1 vccd1 _07314_ sky130_fd_sc_hd__or2_1
XFILLER_0_45_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14523__A net1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19943_ clknet_leaf_46_clk _00887_ net1376 vssd1 vssd1 vccd1 vccd1 ag2.body\[453\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_103_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15066_ _04552_ _05076_ net65 vssd1 vssd1 vccd1 vccd1 _01560_ sky130_fd_sc_hd__and3_2
XANTENNA__11866__B net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12278_ _07232_ _07247_ vssd1 vssd1 vccd1 vccd1 _07248_ sky130_fd_sc_hd__nor2_1
XANTENNA__10770__B net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14017_ net1036 _04162_ ag2.body\[462\] net800 vssd1 vssd1 vccd1 vccd1 _08178_ sky130_fd_sc_hd__o22a_1
XANTENNA_clkbuf_leaf_88_clk_X clknet_leaf_88_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11229_ net1076 control.body\[862\] vssd1 vssd1 vccd1 vccd1 _06202_ sky130_fd_sc_hd__or2_1
X_19874_ clknet_leaf_82_clk _00818_ net1479 vssd1 vssd1 vccd1 vccd1 ag2.body\[512\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_4_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19120__CLK clknet_leaf_141_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18825_ clknet_leaf_2_clk img_gen.tracker.next_frame\[263\] net1249 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[263\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__17553__B net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_131_clk_X clknet_leaf_131_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16471__A1 net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18756_ clknet_leaf_15_clk img_gen.tracker.next_frame\[194\] net1312 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[194\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__13285__A1 net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12088__A2 net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15968_ ag2.body\[139\] net212 _01658_ ag2.body\[131\] vssd1 vssd1 vccd1 vccd1 _01197_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_91_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17707_ obsg2.obstacleArray\[130\] net448 vssd1 vssd1 vccd1 vccd1 _03386_ sky130_fd_sc_hd__or2_1
X_14919_ control.body\[1078\] net170 _01542_ net2205 vssd1 vssd1 vccd1 vccd1 _00264_
+ sky130_fd_sc_hd__a22o_1
X_18687_ clknet_leaf_28_clk img_gen.tracker.next_frame\[125\] net1337 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[125\] sky130_fd_sc_hd__dfrtp_1
X_15899_ ag2.body\[206\] net133 _01650_ ag2.body\[198\] vssd1 vssd1 vccd1 vccd1 _01136_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11835__A2 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15641__X _01623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17420__B1 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17638_ ag2.body\[163\] net852 vssd1 vssd1 vccd1 vccd1 _03317_ sky130_fd_sc_hd__nand2_1
XFILLER_0_77_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18838__CLK clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16774__A2 net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_1418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10010__B net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17569_ ag2.body\[579\] net716 net689 ag2.body\[583\] _03247_ vssd1 vssd1 vccd1 vccd1
+ _03248_ sky130_fd_sc_hd__a221o_1
XFILLER_0_74_934 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19308_ clknet_leaf_99_clk _00252_ net1445 vssd1 vssd1 vccd1 vccd1 control.body\[1082\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20580_ clknet_leaf_107_clk _01437_ _00044_ vssd1 vssd1 vccd1 vccd1 sound_gen.osc1.count\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_136_4470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_4481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16526__A2 net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_132_4334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_132_4345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19239_ clknet_leaf_83_clk _00183_ net1480 vssd1 vssd1 vccd1 vccd1 ag2.body\[102\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_132_4356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11122__A net1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_1573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_41_1584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17487__B1 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14433__A net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1039_A net1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09527__A net1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10680__B net1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_1327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout402 net403 vssd1 vssd1 vccd1 vccd1 net402 sky130_fd_sc_hd__clkbuf_4
XANTENNA__17239__B1 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout413 _01901_ vssd1 vssd1 vccd1 vccd1 net413 sky130_fd_sc_hd__buf_4
XANTENNA__13049__A net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout424 net425 vssd1 vssd1 vccd1 vccd1 net424 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_54_1967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout435 net436 vssd1 vssd1 vccd1 vccd1 net435 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout1206_A net1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20014_ clknet_leaf_59_clk _00958_ net1467 vssd1 vssd1 vccd1 vccd1 ag2.body\[380\]
+ sky130_fd_sc_hd__dfrtp_4
Xfanout446 net448 vssd1 vssd1 vccd1 vccd1 net446 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_96_1514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input4_A gpio_in[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout457 net458 vssd1 vssd1 vccd1 vccd1 net457 sky130_fd_sc_hd__buf_2
X_09825_ net1179 control.body\[922\] vssd1 vssd1 vccd1 vccd1 _04798_ sky130_fd_sc_hd__or2_1
XANTENNA__13991__B net67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18451__A2 _04791_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout468 _06648_ vssd1 vssd1 vccd1 vccd1 net468 sky130_fd_sc_hd__clkbuf_4
XANTENNA__17463__B net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout666_A net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09756_ ag2.body\[212\] net1140 vssd1 vssd1 vccd1 vccd1 _04729_ sky130_fd_sc_hd__or2_1
XANTENNA__13276__A1 net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17750__Y _03429_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09687_ _04656_ _04657_ _04658_ _04659_ vssd1 vssd1 vccd1 vccd1 _04660_ sky130_fd_sc_hd__or4_2
XANTENNA__11826__A2 net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout454_X net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout833_A net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14298__A2_N net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1196_X net1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13028__A1 net238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16765__A2 net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19841__RESET_B net1414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19763__CLK clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11016__B net1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15973__B1 net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_0__f_clk_A clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout621_X net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout719_X net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout42 net43 vssd1 vssd1 vccd1 vccd1 net42 sky130_fd_sc_hd__buf_2
X_10600_ _04236_ _04237_ _04238_ _04946_ _05178_ vssd1 vssd1 vccd1 vccd1 _05573_ sky130_fd_sc_hd__o41a_2
XFILLER_0_49_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout53 net54 vssd1 vssd1 vccd1 vccd1 net53 sky130_fd_sc_hd__clkbuf_8
X_11580_ net760 _06552_ _06549_ _06485_ vssd1 vssd1 vccd1 vccd1 _06553_ sky130_fd_sc_hd__o211a_1
Xfanout64 _08131_ vssd1 vssd1 vccd1 vccd1 net64 sky130_fd_sc_hd__clkbuf_2
XANTENNA__17714__A1 net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout75 net79 vssd1 vssd1 vccd1 vccd1 net75 sky130_fd_sc_hd__buf_2
XFILLER_0_37_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout86 net87 vssd1 vssd1 vccd1 vccd1 net86 sky130_fd_sc_hd__buf_2
X_10531_ net1133 control.body\[916\] vssd1 vssd1 vccd1 vccd1 _05504_ sky130_fd_sc_hd__nand2_1
XFILLER_0_9_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout97 net100 vssd1 vssd1 vccd1 vccd1 net97 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_52_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12773__D _07486_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_115_3820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17919__A net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_115_3831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17190__A2 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_115_3842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13250_ net2025 net648 _07811_ _07812_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[395\]
+ sky130_fd_sc_hd__a31o_1
X_10462_ _04686_ _05424_ _05429_ _05434_ vssd1 vssd1 vccd1 vccd1 _05435_ sky130_fd_sc_hd__or4_4
XFILLER_0_17_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13200__A1 net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout990_X net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17638__B net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_3706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_111_3717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12201_ net317 _07170_ net480 vssd1 vssd1 vccd1 vccd1 _07173_ sky130_fd_sc_hd__a21o_1
XANTENNA__09955__A1 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13181_ net1866 net646 _07781_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[357\]
+ sky130_fd_sc_hd__and3_1
XANTENNA__09955__B2 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10393_ net1135 control.body\[1060\] vssd1 vssd1 vccd1 vccd1 _05366_ sky130_fd_sc_hd__nand2_1
XFILLER_0_33_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14343__A net1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19143__CLK clknet_leaf_132_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12132_ img_gen.tracker.frame\[552\] net622 net605 img_gen.tracker.frame\[555\] _07103_
+ vssd1 vssd1 vccd1 vccd1 _07104_ sky130_fd_sc_hd__o221a_1
XANTENNA__16150__B1 net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11686__B net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12063_ net559 _07034_ net468 vssd1 vssd1 vccd1 vccd1 _07035_ sky130_fd_sc_hd__o21a_1
X_16940_ ag2.body\[524\] net711 net936 _04192_ _02618_ vssd1 vssd1 vccd1 vccd1 _02619_
+ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_109_3635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_2470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_3646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11014_ ag2.body\[596\] net1120 vssd1 vssd1 vccd1 vccd1 _05987_ sky130_fd_sc_hd__xor2_1
XANTENNA__09724__X _04697_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_3657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16871_ ag2.body\[465\] net730 net858 _04165_ vssd1 vssd1 vccd1 vccd1 _02550_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__19293__CLK clknet_leaf_98_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout980 net982 vssd1 vssd1 vccd1 vccd1 net980 sky130_fd_sc_hd__clkbuf_8
X_18610_ clknet_leaf_146_clk img_gen.tracker.next_frame\[48\] net1241 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[48\] sky130_fd_sc_hd__dfrtp_1
Xfanout991 net995 vssd1 vssd1 vccd1 vccd1 net991 sky130_fd_sc_hd__clkbuf_8
X_15822_ ag2.body\[264\] net201 _01643_ ag2.body\[256\] vssd1 vssd1 vccd1 vccd1 _01066_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_5_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09443__Y _04416_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19590_ clknet_leaf_118_clk _00534_ net1386 vssd1 vssd1 vccd1 vccd1 control.body\[804\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_5_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13267__A1 net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19929__RESET_B net1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15753_ ag2.body\[331\] net215 _01635_ ag2.body\[323\] vssd1 vssd1 vccd1 vccd1 _01005_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_87_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18541_ clknet_leaf_135_clk _00067_ net1298 vssd1 vssd1 vccd1 vccd1 img_gen.updater.commands.count\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14804__A2_N ag2.body\[290\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12965_ net232 _07678_ _07679_ net2119 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[243\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11817__A2 net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16205__A1 _01743_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_83_2842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15461__X _01603_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_83_2853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11916_ net467 _06879_ _06882_ vssd1 vssd1 vccd1 vccd1 _06888_ sky130_fd_sc_hd__or3_1
X_14704_ net1038 ag2.body\[236\] vssd1 vssd1 vccd1 vccd1 _08865_ sky130_fd_sc_hd__xor2_1
X_18472_ net724 _03953_ _03957_ vssd1 vssd1 vccd1 vccd1 _01425_ sky130_fd_sc_hd__a21oi_1
X_15684_ ag2.body\[398\] net141 _01627_ ag2.body\[390\] vssd1 vssd1 vccd1 vccd1 _00944_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__10111__A net1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13019__A1 net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_83_2864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12896_ _07448_ net339 net386 vssd1 vssd1 vccd1 vccd1 _07647_ sky130_fd_sc_hd__and3b_2
XFILLER_0_34_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_2263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17423_ ag2.body\[113\] net876 vssd1 vssd1 vccd1 vccd1 _03102_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_64_2274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14635_ net832 ag2.body\[577\] _04212_ net1035 _08793_ vssd1 vssd1 vccd1 vccd1 _08796_
+ sky130_fd_sc_hd__a221o_1
X_11847_ _06812_ _06814_ _06816_ _06818_ net560 net473 vssd1 vssd1 vccd1 vccd1 _06819_
+ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_64_2285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_2138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10518__A2_N net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_60_2149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20487__RESET_B net1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14566_ net986 _04126_ ag2.body\[359\] net797 vssd1 vssd1 vccd1 vccd1 _08727_ sky130_fd_sc_hd__a22o_1
X_17354_ ag2.body\[3\] _03032_ vssd1 vssd1 vccd1 vccd1 _03033_ sky130_fd_sc_hd__nor2_1
XFILLER_0_126_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17705__A1 net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16508__A2 _02059_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11778_ img_gen.tracker.frame\[158\] net626 net603 img_gen.tracker.frame\[161\] _06749_
+ vssd1 vssd1 vccd1 vccd1 _06750_ sky130_fd_sc_hd__o221a_1
XFILLER_0_3_1440 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17116__A2_N net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_844 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14519__A1 net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16305_ obsg2.obstacleArray\[100\] net404 _01983_ net418 vssd1 vssd1 vccd1 vccd1
+ _01984_ sky130_fd_sc_hd__o211a_1
X_13517_ img_gen.tracker.frame\[557\] net657 _07917_ vssd1 vssd1 vccd1 vccd1 _07918_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_125_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14519__B2 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17285_ ag2.body\[308\] net966 vssd1 vssd1 vccd1 vccd1 _02964_ sky130_fd_sc_hd__xor2_1
XFILLER_0_43_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10729_ ag2.body\[248\] net787 net746 ag2.body\[255\] vssd1 vssd1 vccd1 vccd1 _05702_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__17829__A net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14497_ net991 _04086_ ag2.body\[259\] net820 vssd1 vssd1 vccd1 vccd1 _08658_ sky130_fd_sc_hd__a22o_1
XANTENNA__12038__A net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16236_ _01913_ _01914_ net415 vssd1 vssd1 vccd1 vccd1 _01915_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19024_ clknet_leaf_1_clk img_gen.tracker.next_frame\[462\] net1246 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[462\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_899 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13448_ net257 _07890_ _07891_ net1633 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[514\]
+ sky130_fd_sc_hd__a22o_1
Xclkload12 clknet_leaf_143_clk vssd1 vssd1 vccd1 vccd1 clkload12/Y sky130_fd_sc_hd__clkinv_8
XTAP_TAPCELL_ROW_77_2657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload23 clknet_leaf_13_clk vssd1 vssd1 vccd1 vccd1 clkload23/Y sky130_fd_sc_hd__inv_6
XTAP_TAPCELL_ROW_77_2668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12980__B _07505_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload34 clknet_leaf_140_clk vssd1 vssd1 vccd1 vccd1 clkload34/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_23_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_1447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_77_2679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload45 clknet_leaf_27_clk vssd1 vssd1 vccd1 vccd1 clkload45/Y sky130_fd_sc_hd__inv_6
XANTENNA__17469__B1 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload56 clknet_leaf_39_clk vssd1 vssd1 vccd1 vccd1 clkload56/Y sky130_fd_sc_hd__clkinv_8
X_16167_ obsg2.obstacleArray\[13\] net430 vssd1 vssd1 vccd1 vccd1 _01846_ sky130_fd_sc_hd__or2_1
Xclkload67 clknet_leaf_42_clk vssd1 vssd1 vccd1 vccd1 clkload67/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_109_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13379_ net228 _07864_ _07865_ net1896 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[471\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__10781__A net1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_58_2078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload78 clknet_leaf_120_clk vssd1 vssd1 vccd1 vccd1 clkload78/Y sky130_fd_sc_hd__clkinv_4
XTAP_TAPCELL_ROW_58_2089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10556__A2 _05509_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15118_ control.body\[903\] net146 _01554_ net2523 vssd1 vssd1 vccd1 vccd1 _00441_
+ sky130_fd_sc_hd__a22o_1
Xclkload89 clknet_leaf_107_clk vssd1 vssd1 vccd1 vccd1 clkload89/Y sky130_fd_sc_hd__clkinvlp_4
XANTENNA_clkbuf_leaf_53_clk_A clknet_4_6__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16098_ _01728_ _01751_ _01759_ _01767_ _01776_ vssd1 vssd1 vccd1 vccd1 _01777_ sky130_fd_sc_hd__o32a_1
XFILLER_0_107_1160 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19926_ clknet_leaf_51_clk _00870_ net1369 vssd1 vssd1 vccd1 vccd1 ag2.body\[468\]
+ sky130_fd_sc_hd__dfrtp_4
X_15049_ net2631 net163 _01558_ net2383 vssd1 vssd1 vccd1 vccd1 _00378_ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_4_11__f_clk_A clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17283__B net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19857_ clknet_leaf_93_clk _00801_ net1412 vssd1 vssd1 vccd1 vccd1 ag2.body\[543\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_3_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09610_ _04575_ _04576_ _04578_ _04579_ vssd1 vssd1 vccd1 vccd1 _04583_ sky130_fd_sc_hd__or4_1
XANTENNA__17641__B1 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_4013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_68_clk_A clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18808_ clknet_leaf_4_clk img_gen.tracker.next_frame\[246\] net1259 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[246\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_121_4024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19788_ clknet_leaf_127_clk _00732_ net1328 vssd1 vssd1 vccd1 vccd1 ag2.body\[602\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_30_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18660__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19786__CLK clknet_leaf_127_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09532__A_N net1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_111_clk_A clknet_4_10__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09541_ net1063 control.body\[1031\] vssd1 vssd1 vccd1 vccd1 _04514_ sky130_fd_sc_hd__or2_1
X_18739_ clknet_leaf_142_clk img_gen.tracker.next_frame\[177\] net1261 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[177\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_92_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15812__A _04985_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09472_ net917 net913 vssd1 vssd1 vccd1 vccd1 _04445_ sky130_fd_sc_hd__nor2_4
XTAP_TAPCELL_ROW_138_4521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_1466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16747__A2 net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09882__B1 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_4532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_4565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19252__RESET_B net1484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_4576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_4407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_126_clk_A clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_134_4418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13332__A net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20632_ net1549 vssd1 vssd1 vccd1 vccd1 gpio_out[27] sky130_fd_sc_hd__buf_2
XFILLER_0_4_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_956 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10675__B net1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14329__A1_N net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15707__B1 _01629_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12593__D _07312_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload6 clknet_4_12__leaf_clk vssd1 vssd1 vccd1 vccd1 clkload6/Y sky130_fd_sc_hd__clkinvlp_4
X_20563_ clknet_leaf_109_clk toggle1.nextDisplayOut\[3\] net1420 vssd1 vssd1 vccd1
+ vccd1 ssdec1.in\[3\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__17172__A2 net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19166__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1156_A ag2.y\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_574 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11992__B2 net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09809__X _04782_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20494_ clknet_leaf_24_clk _01381_ net1360 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[130\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_116_398 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_3160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_3171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1323_A net1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16132__B1 _01728_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_1271 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout783_A net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_1439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout210 net218 vssd1 vssd1 vccd1 vccd1 net210 sky130_fd_sc_hd__buf_2
XANTENNA__13497__A1 net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1111_X net1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1208 net1213 vssd1 vssd1 vccd1 vccd1 net1208 sky130_fd_sc_hd__buf_4
Xfanout221 net222 vssd1 vssd1 vccd1 vccd1 net221 sky130_fd_sc_hd__buf_1
Xfanout1219 net1221 vssd1 vssd1 vccd1 vccd1 net1219 sky130_fd_sc_hd__buf_4
XFILLER_0_61_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1209_X net1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout232 net233 vssd1 vssd1 vccd1 vccd1 net232 sky130_fd_sc_hd__clkbuf_4
Xfanout243 net244 vssd1 vssd1 vccd1 vccd1 net243 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout950_A obsg2.randCord\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20293__CLK clknet_leaf_37_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout571_X net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout254 net260 vssd1 vssd1 vccd1 vccd1 net254 sky130_fd_sc_hd__buf_2
Xfanout265 net266 vssd1 vssd1 vccd1 vccd1 net265 sky130_fd_sc_hd__buf_2
XANTENNA__16435__A1 net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout669_X net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout276 net279 vssd1 vssd1 vccd1 vccd1 net276 sky130_fd_sc_hd__clkbuf_4
XANTENNA__17761__X _03440_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17632__B1 net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09808_ _04551_ _04759_ _04766_ _04771_ _04780_ vssd1 vssd1 vccd1 vccd1 _04781_ sky130_fd_sc_hd__o32a_1
Xfanout287 net288 vssd1 vssd1 vccd1 vccd1 net287 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_138_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout298 _03546_ vssd1 vssd1 vccd1 vccd1 net298 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_104_3510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16986__A2 net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09739_ ag2.body\[354\] net1185 vssd1 vssd1 vccd1 vccd1 _04712_ sky130_fd_sc_hd__xor2_1
XFILLER_0_74_1620 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1480_X net1480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout836_X net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_3_4_0_clk_X clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11027__A net1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12750_ net305 _07578_ vssd1 vssd1 vccd1 vccd1 _07579_ sky130_fd_sc_hd__nor2_1
XFILLER_0_55_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16738__A2 net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09873__B1 _04832_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11701_ _06641_ _06644_ _06671_ vssd1 vssd1 vccd1 vccd1 _06673_ sky130_fd_sc_hd__and3_2
XFILLER_0_70_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14749__A1 net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14749__B2 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12681_ _06671_ _07545_ vssd1 vssd1 vccd1 vccd1 _07546_ sky130_fd_sc_hd__or2_2
X_14420_ net976 _04195_ _04196_ net1021 vssd1 vssd1 vccd1 vccd1 _08581_ sky130_fd_sc_hd__a22o_1
X_11632_ net504 _06602_ _06604_ net1123 vssd1 vssd1 vccd1 vccd1 _06605_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_13_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_117_3904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17950__A4 _03577_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_1383 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14351_ net1000 ag2.body\[400\] vssd1 vssd1 vccd1 vccd1 _08512_ sky130_fd_sc_hd__xor2_1
XFILLER_0_119_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11563_ obsg2.obstacleArray\[72\] obsg2.obstacleArray\[73\] obsg2.obstacleArray\[76\]
+ obsg2.obstacleArray\[77\] net1123 net510 vssd1 vssd1 vccd1 vccd1 _06536_ sky130_fd_sc_hd__mux4_1
XFILLER_0_9_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xwire633 _06461_ vssd1 vssd1 vccd1 vccd1 net633 sky130_fd_sc_hd__buf_4
X_13302_ net281 _07833_ _07834_ net2040 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[425\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_108_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10514_ ag2.body\[102\] net1089 vssd1 vssd1 vccd1 vccd1 _05487_ sky130_fd_sc_hd__xnor2_1
X_17070_ ag2.body\[26\] net722 net688 ag2.body\[31\] vssd1 vssd1 vccd1 vccd1 _02749_
+ sky130_fd_sc_hd__a22o_1
X_14282_ net845 ag2.body\[136\] ag2.body\[143\] net796 _08438_ vssd1 vssd1 vccd1 vccd1
+ _08443_ sky130_fd_sc_hd__a221o_1
XFILLER_0_11_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11494_ _06463_ _06466_ vssd1 vssd1 vccd1 vccd1 _06467_ sky130_fd_sc_hd__nor2_1
XANTENNA__16272__B net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16021_ net355 vssd1 vssd1 vccd1 vccd1 _01700_ sky130_fd_sc_hd__inv_2
XFILLER_0_80_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11697__A net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13233_ net259 _07426_ _07805_ net1750 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[385\]
+ sky130_fd_sc_hd__a22o_1
X_10445_ _04552_ _05415_ _05416_ _05417_ vssd1 vssd1 vccd1 vccd1 _05418_ sky130_fd_sc_hd__and4_1
XFILLER_0_27_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_72_2510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13164_ net668 _07773_ vssd1 vssd1 vccd1 vccd1 _07774_ sky130_fd_sc_hd__nor2_1
X_10376_ ag2.body\[106\] net1187 vssd1 vssd1 vccd1 vccd1 _05349_ sky130_fd_sc_hd__xor2_1
XANTENNA__16699__S net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12115_ img_gen.tracker.frame\[156\] net627 net609 img_gen.tracker.frame\[159\] _07086_
+ vssd1 vssd1 vccd1 vccd1 _07087_ sky130_fd_sc_hd__a221o_1
XFILLER_0_104_1344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_1198 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14360__X _08521_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17972_ net298 _03594_ vssd1 vssd1 vccd1 vccd1 _03595_ sky130_fd_sc_hd__nand2_1
XANTENNA__10106__A net1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13095_ net674 _07740_ vssd1 vssd1 vccd1 vccd1 _07741_ sky130_fd_sc_hd__nor2_1
XFILLER_0_97_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19711_ clknet_leaf_134_clk _00655_ net1306 vssd1 vssd1 vccd1 vccd1 control.body\[685\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09454__X _04427_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16923_ ag2.body\[374\] net940 vssd1 vssd1 vccd1 vccd1 _02602_ sky130_fd_sc_hd__xor2_1
X_12046_ img_gen.tracker.frame\[252\] net628 net554 img_gen.tracker.frame\[258\] vssd1
+ vssd1 vccd1 vccd1 _07018_ sky130_fd_sc_hd__a22o_1
XFILLER_0_137_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19642_ clknet_leaf_133_clk _00586_ net1391 vssd1 vssd1 vccd1 vccd1 control.body\[744\]
+ sky130_fd_sc_hd__dfrtp_1
X_16854_ _02525_ _02530_ _02532_ vssd1 vssd1 vccd1 vccd1 _02533_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_85_2904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20311__Q ag2.randCord\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_2926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15805_ ag2.body\[281\] net206 _01641_ ag2.body\[273\] vssd1 vssd1 vccd1 vccd1 _01051_
+ sky130_fd_sc_hd__a22o_1
X_19573_ clknet_leaf_116_clk _00517_ net1385 vssd1 vssd1 vccd1 vccd1 control.body\[819\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_66_2325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13997_ ag2.body\[133\] net212 _08160_ ag2.body\[125\] vssd1 vssd1 vccd1 vccd1 _00214_
+ sky130_fd_sc_hd__a22o_1
X_16785_ net381 _02452_ vssd1 vssd1 vccd1 vccd1 _02464_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_66_2336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20616__1559 vssd1 vssd1 vccd1 vccd1 net1559 _20616__1559/LO sky130_fd_sc_hd__conb_1
XANTENNA__09459__A3 net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_2347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15632__A _06028_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18524_ clknet_leaf_138_clk img_gen.updater.update.next\[1\] net1299 vssd1 vssd1
+ vccd1 vccd1 img_gen.updater.commands.mode\[1\] sky130_fd_sc_hd__dfrtp_4
X_15736_ ag2.body\[348\] net198 _01633_ ag2.body\[340\] vssd1 vssd1 vccd1 vccd1 _00990_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_73_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12948_ net246 _07670_ _07671_ net1964 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[234\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__16729__A2 net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18455_ _04645_ _03841_ vssd1 vssd1 vccd1 vccd1 _03944_ sky130_fd_sc_hd__nand2b_1
X_15667_ ag2.body\[415\] net143 _01625_ ag2.body\[407\] vssd1 vssd1 vccd1 vccd1 _00929_
+ sky130_fd_sc_hd__a22o_1
X_12879_ net267 _07425_ _07638_ _07640_ net1642 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[196\]
+ sky130_fd_sc_hd__a32o_1
XANTENNA__14248__A net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13152__A net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19189__CLK clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17406_ ag2.body\[44\] net959 vssd1 vssd1 vccd1 vccd1 _03085_ sky130_fd_sc_hd__xor2_1
X_14618_ net817 ag2.body\[59\] ag2.body\[62\] net798 _08774_ vssd1 vssd1 vccd1 vccd1
+ _08779_ sky130_fd_sc_hd__a221o_1
XFILLER_0_51_1461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15598_ ag2.body\[464\] net121 _01619_ ag2.body\[456\] vssd1 vssd1 vccd1 vccd1 _00866_
+ sky130_fd_sc_hd__a22o_1
X_18386_ net326 _03796_ _03797_ _03874_ _03875_ vssd1 vssd1 vccd1 vccd1 _03876_ sky130_fd_sc_hd__o221ai_1
XANTENNA__13412__A1 net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_79_2719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17337_ _03010_ _03013_ vssd1 vssd1 vccd1 vccd1 _03016_ sky130_fd_sc_hd__or2_1
X_14549_ net808 ag2.body\[245\] ag2.body\[247\] net795 _08709_ vssd1 vssd1 vccd1 vccd1
+ _08710_ sky130_fd_sc_hd__a221o_1
XANTENNA__12991__A net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16463__A net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15165__A1 control.body\[848\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload101 clknet_leaf_99_clk vssd1 vssd1 vccd1 vccd1 clkload101/Y sky130_fd_sc_hd__clkinv_2
X_17268_ _04079_ net885 net726 ag2.body\[250\] vssd1 vssd1 vccd1 vccd1 _02947_ sky130_fd_sc_hd__o22a_1
XFILLER_0_71_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkload112 clknet_leaf_59_clk vssd1 vssd1 vccd1 vccd1 clkload112/Y sky130_fd_sc_hd__bufinv_16
XFILLER_0_3_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload123 clknet_leaf_81_clk vssd1 vssd1 vccd1 vccd1 clkload123/Y sky130_fd_sc_hd__inv_4
XFILLER_0_70_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19007_ clknet_leaf_1_clk img_gen.tracker.next_frame\[445\] net1244 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[445\] sky130_fd_sc_hd__dfrtp_1
X_16219_ net537 _01889_ _01897_ _01737_ vssd1 vssd1 vccd1 vccd1 _01898_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_52_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17199_ ag2.body\[182\] net697 net691 ag2.body\[183\] vssd1 vssd1 vccd1 vccd1 _02878_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_113_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_127_4200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_4211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_1276 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15468__A2 net90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08972_ ag2.body\[61\] vssd1 vssd1 vccd1 vccd1 _03997_ sky130_fd_sc_hd__inv_2
XANTENNA__14711__A net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16402__S net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13479__A1 net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19909_ clknet_leaf_56_clk _00853_ net1458 vssd1 vssd1 vccd1 vccd1 ag2.body\[483\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__09805__A net1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold18 control.detect3.Q\[0\] vssd1 vssd1 vccd1 vccd1 net1580 sky130_fd_sc_hd__dlygate4sd3_1
Xhold29 img_gen.tracker.frame\[326\] vssd1 vssd1 vccd1 vccd1 net1591 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_32_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout197_A net200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17614__B1 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_1626 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13046__B net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout364_A _02068_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09524_ net1051 control.body\[839\] vssd1 vssd1 vccd1 vccd1 _04497_ sky130_fd_sc_hd__nand2_1
XFILLER_0_17_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12454__A2 net1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09540__A net1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_208 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09455_ net901 net907 vssd1 vssd1 vccd1 vccd1 _04428_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout531_A net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_26_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_26_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout629_A _06473_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09386_ net273 _04364_ _04377_ vssd1 vssd1 vccd1 vccd1 _01410_ sky130_fd_sc_hd__nor3_1
XANTENNA__13403__A1 net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18556__CLK clknet_leaf_43_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_3211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10217__A1 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20615_ net1558 vssd1 vssd1 vccd1 vccd1 gpio_oeb[27] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_95_3222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10217__B2 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_3233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1061_X net1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19801__CLK clknet_leaf_124_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1440_A net1442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout417_X net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1159_X net1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09539__X _04512_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_91_3108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20546_ clknet_leaf_105_clk _01411_ _00020_ vssd1 vssd1 vccd1 vccd1 sound_gen.osc1.stayCount\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__15156__B2 control.body\[848\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17188__B net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout998_A net999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_1355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20477_ clknet_leaf_39_clk _01364_ net1352 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[113\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__12406__A net1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10230_ ag2.body\[563\] net1150 vssd1 vssd1 vccd1 vccd1 _05203_ sky130_fd_sc_hd__xor2_1
XANTENNA_fanout786_X net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09418__C obsg2.obstacleCount\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10161_ ag2.body\[579\] net1150 vssd1 vssd1 vccd1 vccd1 _05134_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_89_3026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_3037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1005 ag2.randCord\[0\] vssd1 vssd1 vccd1 vccd1 net1005 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_7_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1016 net1018 vssd1 vssd1 vccd1 vccd1 net1016 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_89_3048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1027 net1029 vssd1 vssd1 vccd1 vccd1 net1027 sky130_fd_sc_hd__buf_4
XANTENNA__09715__A net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout953_X net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1038 net1039 vssd1 vssd1 vccd1 vccd1 net1038 sky130_fd_sc_hd__buf_4
X_10092_ net1148 control.body\[795\] vssd1 vssd1 vccd1 vccd1 _05065_ sky130_fd_sc_hd__or2_1
Xfanout1049 net1051 vssd1 vssd1 vccd1 vccd1 net1049 sky130_fd_sc_hd__clkbuf_4
XANTENNA__17605__B1 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09434__B net1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17932__A _01700_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13920_ ag2.body\[64\] net133 _08152_ ag2.body\[56\] vssd1 vssd1 vccd1 vccd1 _00145_
+ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout65_X net65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20039__CLK clknet_leaf_66_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13851_ ag2.body\[15\] net116 _08133_ ag2.body\[7\] vssd1 vssd1 vccd1 vccd1 _00095_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_57_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19920__Q ag2.body\[478\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12802_ net668 _07603_ vssd1 vssd1 vccd1 vccd1 _07604_ sky130_fd_sc_hd__nor2_1
XANTENNA__18466__C net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16570_ obsg2.obstacleArray\[124\] obsg2.obstacleArray\[125\] net444 vssd1 vssd1
+ vccd1 vccd1 _02249_ sky130_fd_sc_hd__mux2_1
X_13782_ img_gen.updater.commands.count\[12\] img_gen.updater.commands.count\[11\]
+ _08088_ vssd1 vssd1 vccd1 vccd1 _08091_ sky130_fd_sc_hd__and3_1
X_10994_ ag2.body\[339\] net1165 vssd1 vssd1 vccd1 vccd1 _05967_ sky130_fd_sc_hd__xor2_1
XFILLER_0_96_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09450__A net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_366 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__20079__RESET_B net1492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12733_ net683 _07570_ vssd1 vssd1 vccd1 vccd1 _07571_ sky130_fd_sc_hd__nor2_1
X_15521_ ag2.body\[541\] net156 _01609_ ag2.body\[533\] vssd1 vssd1 vccd1 vccd1 _00799_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__14068__A net1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10596__A net1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11044__X _06017_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20189__CLK clknet_leaf_88_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18240_ _03681_ net35 vssd1 vssd1 vccd1 vccd1 _03759_ sky130_fd_sc_hd__nor2_1
X_15452_ _05452_ net63 vssd1 vssd1 vccd1 vccd1 _01602_ sky130_fd_sc_hd__and2_2
X_12664_ net245 _07536_ _07537_ net1773 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[84\]
+ sky130_fd_sc_hd__a22o_1
X_14403_ net1027 net925 vssd1 vssd1 vccd1 vccd1 _08564_ sky130_fd_sc_hd__nand2_1
XFILLER_0_65_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11615_ net508 _06585_ _06587_ net475 vssd1 vssd1 vccd1 vccd1 _06588_ sky130_fd_sc_hd__o211a_1
XFILLER_0_108_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11979__X _06951_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18171_ obsg2.obstacleArray\[82\] _03724_ net531 vssd1 vssd1 vccd1 vccd1 _01333_
+ sky130_fd_sc_hd__o21a_1
X_15383_ net2636 net82 _01595_ net2274 vssd1 vssd1 vccd1 vccd1 _00675_ sky130_fd_sc_hd__a22o_1
X_12595_ _07431_ _07498_ vssd1 vssd1 vccd1 vccd1 _07499_ sky130_fd_sc_hd__nor2_1
XFILLER_0_4_1590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11956__A1 net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14334_ net818 ag2.body\[427\] ag2.body\[431\] net792 vssd1 vssd1 vccd1 vccd1 _08495_
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_110_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17122_ ag2.body\[517\] net952 vssd1 vssd1 vccd1 vccd1 _02801_ sky130_fd_sc_hd__nand2_1
X_11546_ net506 _06515_ _06518_ vssd1 vssd1 vccd1 vccd1 _06519_ sky130_fd_sc_hd__o21a_1
XFILLER_0_135_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_564 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17053_ ag2.body\[72\] net739 net945 _04009_ vssd1 vssd1 vccd1 vccd1 _02732_ sky130_fd_sc_hd__a22o_1
X_14265_ net999 ag2.body\[8\] vssd1 vssd1 vccd1 vccd1 _08426_ sky130_fd_sc_hd__or2_1
XFILLER_0_64_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11477_ ag2.body\[493\] net1114 vssd1 vssd1 vccd1 vccd1 _06450_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_55_2004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_2015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16004_ _01678_ _01682_ _01677_ vssd1 vssd1 vccd1 vccd1 _01683_ sky130_fd_sc_hd__a21o_1
XANTENNA__18097__B1 net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13216_ img_gen.tracker.frame\[376\] net658 vssd1 vssd1 vccd1 vccd1 _07798_ sky130_fd_sc_hd__and2_1
XFILLER_0_122_176 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10428_ net1060 control.body\[1071\] vssd1 vssd1 vccd1 vccd1 _05401_ sky130_fd_sc_hd__nand2_1
X_14196_ net834 ag2.body\[161\] ag2.body\[167\] net793 _08356_ vssd1 vssd1 vccd1 vccd1
+ _08357_ sky130_fd_sc_hd__o221a_1
XFILLER_0_42_1416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13147_ net231 _07764_ _07765_ net2147 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[339\]
+ sky130_fd_sc_hd__a22o_1
X_10359_ ag2.body\[293\] net1115 vssd1 vssd1 vccd1 vccd1 _05332_ sky130_fd_sc_hd__and2b_1
XANTENNA__14531__A net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17955_ net957 net460 net539 net537 vssd1 vssd1 vccd1 vccd1 _03581_ sky130_fd_sc_hd__or4b_1
X_13078_ net244 _07731_ _07732_ net1780 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[303\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_40_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12133__B2 net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12029_ _06690_ _07000_ vssd1 vssd1 vccd1 vccd1 _07001_ sky130_fd_sc_hd__nor2_1
X_16906_ ag2.body\[242\] net726 net711 ag2.body\[244\] _02580_ vssd1 vssd1 vccd1 vccd1
+ _02585_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_68_2409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_1372 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17886_ _04422_ _04445_ _03523_ _03525_ _04537_ vssd1 vssd1 vccd1 vccd1 _03526_ sky130_fd_sc_hd__o311a_1
X_19625_ clknet_leaf_120_clk _00569_ net1392 vssd1 vssd1 vccd1 vccd1 control.body\[775\]
+ sky130_fd_sc_hd__dfrtp_1
X_16837_ ag2.body\[100\] net712 net700 ag2.body\[102\] _02515_ vssd1 vssd1 vccd1 vccd1
+ _02516_ sky130_fd_sc_hd__a221o_1
XANTENNA__17561__B net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16280__C1 net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15622__A2 net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19556_ clknet_leaf_116_clk _00500_ net1389 vssd1 vssd1 vccd1 vccd1 control.body\[834\]
+ sky130_fd_sc_hd__dfrtp_1
X_16768_ _02441_ _02446_ net381 vssd1 vssd1 vccd1 vccd1 _02447_ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14830__B1 _08645_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18507_ net1517 net1511 vssd1 vssd1 vccd1 vccd1 _00038_ sky130_fd_sc_hd__or2_1
XFILLER_0_38_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18579__CLK clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15719_ ag2.body\[366\] net193 _01630_ ag2.body\[358\] vssd1 vssd1 vccd1 vccd1 _00976_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_18_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19487_ clknet_leaf_112_clk net2335 net1418 vssd1 vssd1 vccd1 vccd1 control.body\[909\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_17_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16699_ _02375_ _02377_ net497 vssd1 vssd1 vccd1 vccd1 _02378_ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19824__CLK clknet_4_9__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10998__A2 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09240_ net850 vssd1 vssd1 vccd1 vccd1 _04265_ sky130_fd_sc_hd__inv_2
X_18438_ _03915_ _08138_ vssd1 vssd1 vccd1 vccd1 _03927_ sky130_fd_sc_hd__and2b_1
XFILLER_0_91_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_1387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13397__B1 net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16905__B net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09171_ ag2.body\[534\] vssd1 vssd1 vccd1 vccd1 _04196_ sky130_fd_sc_hd__inv_2
X_18369_ _03859_ _03860_ _03862_ net434 net1923 vssd1 vssd1 vccd1 vccd1 _01393_ sky130_fd_sc_hd__a32o_1
XANTENNA__14706__A net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17127__A2 net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20400_ clknet_leaf_25_clk _01287_ net1340 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[36\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__10953__B net1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20331_ clknet_leaf_108_clk sound_gen.osc1.freq_nxt\[0\] _00007_ vssd1 vssd1 vccd1
+ vccd1 sound_gen.osc1.freq\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_128_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout112_A net113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11130__A net1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18088__B1 net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20262_ clknet_leaf_43_clk _01206_ net1378 vssd1 vssd1 vccd1 vccd1 control.body_update.direction\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_124_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput19 net19 vssd1 vssd1 vccd1 vccd1 gpio_out[18] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_131_Right_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1051 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19204__CLK clknet_leaf_88_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12372__A1 net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20193_ clknet_leaf_88_clk _01137_ net1459 vssd1 vssd1 vccd1 vccd1 ag2.body\[207\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__12911__A3 _07315_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1021_A net1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11580__C1 _06485_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1119_A net1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10349__A2_N net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08955_ ag2.body\[15\] vssd1 vssd1 vccd1 vccd1 _03980_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout481_A net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19614__RESET_B net1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout579_A net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17752__A _02722_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout367_X net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout746_A net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09507_ _04476_ _04477_ _04479_ vssd1 vssd1 vccd1 vccd1 _04480_ sky130_fd_sc_hd__or3_1
XFILLER_0_94_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1118 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20172__RESET_B net1480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1191 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout534_X net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout913_A net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09438_ ag2.body\[7\] net1055 vssd1 vssd1 vccd1 vccd1 _04411_ sky130_fd_sc_hd__or2_1
XFILLER_0_82_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_213 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_427 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16815__B net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11024__B net1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout701_X net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09369_ sound_gen.osc1.stayCount\[20\] _04368_ vssd1 vssd1 vccd1 vccd1 _04370_ sky130_fd_sc_hd__or2_1
XFILLER_0_118_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14616__A net1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11400_ ag2.body\[575\] net1052 vssd1 vssd1 vccd1 vccd1 _06373_ sky130_fd_sc_hd__or2_1
XFILLER_0_62_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12380_ _07341_ _07344_ _07343_ _07236_ vssd1 vssd1 vccd1 vccd1 _07345_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__12060__B1 net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_1439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11331_ net1094 control.body\[661\] vssd1 vssd1 vccd1 vccd1 _06304_ sky130_fd_sc_hd__nand2_1
XFILLER_0_133_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20529_ clknet_leaf_114_clk _01394_ net1398 vssd1 vssd1 vccd1 vccd1 toggle1.bcd_tens\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_133_975 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20615__1558 vssd1 vssd1 vccd1 vccd1 net1558 _20615__1558/LO sky130_fd_sc_hd__conb_1
XFILLER_0_104_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14050_ _08210_ _08205_ _08209_ vssd1 vssd1 vccd1 vccd1 _08211_ sky130_fd_sc_hd__or3b_1
XFILLER_0_127_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11262_ net762 control.body\[772\] control.body\[773\] net754 _06230_ vssd1 vssd1
+ vccd1 vccd1 _06235_ sky130_fd_sc_hd__o221ai_1
XFILLER_0_132_496 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17646__B net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14622__Y _08783_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16629__A1 net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16550__B net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13001_ _07696_ net251 _07694_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[262\]
+ sky130_fd_sc_hd__mux2_1
X_10213_ net1134 control.body\[996\] vssd1 vssd1 vccd1 vccd1 _05186_ sky130_fd_sc_hd__xnor2_1
XANTENNA__14351__A net1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11193_ net1053 control.body\[879\] vssd1 vssd1 vccd1 vccd1 _06166_ sky130_fd_sc_hd__nand2_1
XFILLER_0_98_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10144_ _05115_ _05116_ _05114_ vssd1 vssd1 vccd1 vccd1 _05117_ sky130_fd_sc_hd__a21o_1
XFILLER_0_101_1325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_393 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17740_ _03002_ _03004_ _02491_ _02545_ vssd1 vssd1 vccd1 vccd1 _03419_ sky130_fd_sc_hd__o211a_1
X_10075_ _05037_ _05038_ _05040_ _05046_ vssd1 vssd1 vccd1 vccd1 _05048_ sky130_fd_sc_hd__or4_1
X_14952_ net2217 net174 _01546_ control.body\[1035\] vssd1 vssd1 vccd1 vccd1 _00293_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12666__A2 _07536_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16549__Y _02228_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13903_ ag2.body\[49\] net118 _08150_ ag2.body\[41\] vssd1 vssd1 vccd1 vccd1 _00130_
+ sky130_fd_sc_hd__a22o_1
X_17671_ ag2.body\[448\] net884 vssd1 vssd1 vccd1 vccd1 _03350_ sky130_fd_sc_hd__xor2_1
XANTENNA__17381__B net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11874__B1 net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14883_ control.body\[1110\] net179 _01538_ net2393 vssd1 vssd1 vccd1 vccd1 _00232_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__18721__CLK clknet_leaf_142_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15182__A _04494_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19410_ clknet_leaf_103_clk _00354_ net1427 vssd1 vssd1 vccd1 vccd1 control.body\[976\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_98_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16622_ obsg2.obstacleArray\[38\] obsg2.obstacleArray\[39\] net441 vssd1 vssd1 vccd1
+ vccd1 _02301_ sky130_fd_sc_hd__mux2_1
X_13834_ control.fsm.temp\[2\] net686 _08128_ vssd1 vssd1 vccd1 vccd1 _00083_ sky130_fd_sc_hd__o21a_1
XFILLER_0_43_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19341_ clknet_leaf_100_clk _00285_ net1444 vssd1 vssd1 vccd1 vccd1 control.body\[1051\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11626__B1 net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16553_ net394 _02231_ _02230_ net359 vssd1 vssd1 vccd1 vccd1 _02232_ sky130_fd_sc_hd__a211o_1
X_13765_ img_gen.updater.commands.count\[6\] _08077_ vssd1 vssd1 vccd1 vccd1 _08080_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_58_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10977_ net1077 control.body\[758\] vssd1 vssd1 vccd1 vccd1 _05950_ sky130_fd_sc_hd__or2_1
XFILLER_0_50_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_1590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11215__A net1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15504_ ag2.body\[558\] net113 _01607_ ag2.body\[550\] vssd1 vssd1 vccd1 vccd1 _00784_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__14229__C net1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19272_ clknet_leaf_70_clk _00216_ net1503 vssd1 vssd1 vccd1 vccd1 ag2.body\[135\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_84_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12716_ net683 _07562_ vssd1 vssd1 vccd1 vccd1 _07563_ sky130_fd_sc_hd__nor2_1
XANTENNA__17640__A1_N net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16484_ obsg2.obstacleArray\[45\] _02059_ net401 _02162_ vssd1 vssd1 vccd1 vccd1
+ _02163_ sky130_fd_sc_hd__o211a_1
XANTENNA__18871__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13696_ net892 _08023_ _08037_ vssd1 vssd1 vccd1 vccd1 track.nextCurrScore\[7\] sky130_fd_sc_hd__a21o_1
XANTENNA__13133__C net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19997__CLK clknet_leaf_66_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18223_ obsg2.obstacleArray\[108\] _03750_ net520 vssd1 vssd1 vccd1 vccd1 _01359_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_84_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12647_ _06672_ _07526_ vssd1 vssd1 vccd1 vccd1 _07527_ sky130_fd_sc_hd__nand2_1
X_15435_ ag2.body\[608\] net85 _01600_ ag2.body\[600\] vssd1 vssd1 vccd1 vccd1 _00722_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_66_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17109__A2 net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14526__A net992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11502__X _06475_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13430__A net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18154_ net47 _03582_ _03704_ obsg2.obstacleArray\[74\] vssd1 vssd1 vccd1 vccd1 _03716_
+ sky130_fd_sc_hd__a31o_1
XANTENNA__12051__B1 net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15366_ control.body\[674\] net76 _01593_ net2336 vssd1 vssd1 vccd1 vccd1 _00660_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_108_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12578_ net268 _07488_ _07489_ net2026 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[46\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_80_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10773__B net1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19227__CLK clknet_leaf_75_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17105_ _03976_ net860 net717 ag2.body\[11\] _02783_ vssd1 vssd1 vccd1 vccd1 _02784_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_0_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11529_ net506 _06498_ _06501_ vssd1 vssd1 vccd1 vccd1 _06502_ sky130_fd_sc_hd__o21a_1
XANTENNA__17837__A net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14317_ _08469_ _08470_ _08471_ _08472_ vssd1 vssd1 vccd1 vccd1 _08478_ sky130_fd_sc_hd__a22o_1
X_18085_ net527 _03672_ vssd1 vssd1 vccd1 vccd1 _01299_ sky130_fd_sc_hd__and2_1
X_15297_ control.body\[741\] net76 _01585_ control.body\[733\] vssd1 vssd1 vccd1 vccd1
+ _00599_ sky130_fd_sc_hd__a22o_1
Xhold307 img_gen.tracker.frame\[363\] vssd1 vssd1 vccd1 vccd1 net1869 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold318 img_gen.tracker.frame\[239\] vssd1 vssd1 vccd1 vccd1 net1880 sky130_fd_sc_hd__dlygate4sd3_1
X_17036_ ag2.body\[123\] net856 vssd1 vssd1 vccd1 vccd1 _02715_ sky130_fd_sc_hd__xnor2_1
Xhold329 img_gen.tracker.frame\[184\] vssd1 vssd1 vccd1 vccd1 net1891 sky130_fd_sc_hd__dlygate4sd3_1
X_14248_ net976 ag2.body\[539\] vssd1 vssd1 vccd1 vccd1 _08409_ sky130_fd_sc_hd__xor2_1
XANTENNA__17556__B net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_258 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11885__A net1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14179_ net806 ag2.body\[197\] ag2.body\[198\] net799 _08339_ vssd1 vssd1 vccd1 vccd1
+ _08340_ sky130_fd_sc_hd__a221o_1
XANTENNA__09626__Y _04599_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout809 net810 vssd1 vssd1 vccd1 vccd1 net809 sky130_fd_sc_hd__clkbuf_8
XANTENNA__11562__C1 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19377__CLK clknet_leaf_93_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18987_ clknet_leaf_8_clk img_gen.tracker.next_frame\[425\] net1271 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[425\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__12106__A1 net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1007 control.body\[992\] vssd1 vssd1 vccd1 vccd1 net2569 sky130_fd_sc_hd__dlygate4sd3_1
X_17938_ net516 _03568_ vssd1 vssd1 vccd1 vccd1 _01256_ sky130_fd_sc_hd__nor2_1
Xhold1018 control.body\[1041\] vssd1 vssd1 vccd1 vccd1 net2580 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1029 control.body\[761\] vssd1 vssd1 vccd1 vccd1 net2591 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13308__C net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1380 net1383 vssd1 vssd1 vccd1 vccd1 net1380 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_84_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10668__A1 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10668__B2 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1391 net1392 vssd1 vssd1 vccd1 vccd1 net1391 sky130_fd_sc_hd__clkbuf_4
XANTENNA__15363__Y _01593_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17869_ net2212 _03503_ vssd1 vssd1 vccd1 vccd1 _01241_ sky130_fd_sc_hd__xor2_1
XANTENNA__10013__B _04985_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19608_ clknet_leaf_119_clk net2288 net1391 vssd1 vssd1 vccd1 vccd1 control.body\[790\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_94_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14803__B1 ag2.body\[295\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19539_ clknet_leaf_115_clk _00483_ net1396 vssd1 vssd1 vccd1 vccd1 control.body\[849\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_1331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11093__A1 _04980_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09223_ control.body\[894\] vssd1 vssd1 vccd1 vccd1 _04248_ sky130_fd_sc_hd__inv_2
XFILLER_0_130_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14436__A net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout327_A net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09154_ ag2.body\[495\] vssd1 vssd1 vccd1 vccd1 _04179_ sky130_fd_sc_hd__inv_2
XFILLER_0_17_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_1151 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09085_ ag2.body\[321\] vssd1 vssd1 vccd1 vccd1 _04110_ sky130_fd_sc_hd__inv_2
XANTENNA__17747__A _03420_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14723__X _08884_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1236_A net1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_603 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20314_ clknet_leaf_44_clk obsrand1.next_randY\[0\] net1381 vssd1 vssd1 vccd1 vccd1
+ ag2.randCord\[0\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_9_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15531__A1 ag2.body\[534\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold830 control.body\[1090\] vssd1 vssd1 vccd1 vccd1 net2392 sky130_fd_sc_hd__dlygate4sd3_1
Xhold841 control.body\[661\] vssd1 vssd1 vccd1 vccd1 net2403 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout696_A _04268_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold852 _00518_ vssd1 vssd1 vccd1 vccd1 net2414 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20245_ clknet_leaf_68_clk _01189_ net1496 vssd1 vssd1 vccd1 vccd1 ag2.body\[147\]
+ sky130_fd_sc_hd__dfrtp_4
Xhold863 control.body\[930\] vssd1 vssd1 vccd1 vccd1 net2425 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold874 control.body\[963\] vssd1 vssd1 vccd1 vccd1 net2436 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1024_X net1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1403_A net1404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold885 control.body\[793\] vssd1 vssd1 vccd1 vccd1 net2447 sky130_fd_sc_hd__dlygate4sd3_1
Xhold896 control.body\[763\] vssd1 vssd1 vccd1 vccd1 net2458 sky130_fd_sc_hd__dlygate4sd3_1
X_20176_ clknet_leaf_82_clk _01120_ net1479 vssd1 vssd1 vccd1 vccd1 ag2.body\[222\]
+ sky130_fd_sc_hd__dfrtp_4
X_09987_ _04956_ _04957_ _04958_ _04959_ vssd1 vssd1 vccd1 vccd1 _04960_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout484_X net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout863_A net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15834__A2 net204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08938_ net1003 vssd1 vssd1 vccd1 vccd1 _03963_ sky130_fd_sc_hd__inv_2
XFILLER_0_102_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18233__B1 net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11019__B net1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout749_X net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17587__A2 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1410 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10900_ net1168 control.body\[674\] vssd1 vssd1 vccd1 vccd1 _05873_ sky130_fd_sc_hd__nand2_1
X_11880_ img_gen.tracker.frame\[1\] net623 net590 img_gen.tracker.frame\[10\] vssd1
+ vssd1 vccd1 vccd1 _06852_ sky130_fd_sc_hd__o22a_1
XFILLER_0_135_1454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11608__B1 net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10831_ ag2.body\[306\] net1186 vssd1 vssd1 vccd1 vccd1 _05804_ sky130_fd_sc_hd__xor2_1
XFILLER_0_131_1318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_120_3977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14270__A1 net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout916_X net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_3988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14270__B2 net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13550_ ssdec1.in\[1\] ssdec1.in\[0\] vssd1 vssd1 vccd1 vccd1 _07932_ sky130_fd_sc_hd__nor2_1
X_10762_ control.body\[895\] net1058 vssd1 vssd1 vccd1 vccd1 _05735_ sky130_fd_sc_hd__and2b_1
XANTENNA__18554__SET_B net1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_3398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16547__B1 net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_11_Right_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1486 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12501_ net2074 net650 _07446_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[12\]
+ sky130_fd_sc_hd__and3_1
X_13481_ net666 _07904_ vssd1 vssd1 vccd1 vccd1 _07905_ sky130_fd_sc_hd__nor2_1
X_10693_ ag2.body\[145\] net1211 vssd1 vssd1 vccd1 vccd1 _05666_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_137_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15220_ control.body\[801\] net93 _01576_ net2215 vssd1 vssd1 vccd1 vccd1 _00531_
+ sky130_fd_sc_hd__a22o_1
X_12432_ _07298_ _07386_ _07389_ _07393_ vssd1 vssd1 vccd1 vccd1 _07394_ sky130_fd_sc_hd__or4_1
XFILLER_0_129_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1183 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__20227__CLK clknet_leaf_66_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12584__A1 net250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15151_ net2254 net106 _01568_ net2295 vssd1 vssd1 vccd1 vccd1 _00470_ sky130_fd_sc_hd__a22o_1
X_12363_ _07228_ _07264_ _07267_ vssd1 vssd1 vccd1 vccd1 _07329_ sky130_fd_sc_hd__and3_1
XFILLER_0_22_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11792__C1 net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14102_ _08259_ _08260_ _08261_ _08262_ vssd1 vssd1 vccd1 vccd1 _08263_ sky130_fd_sc_hd__or4_1
XFILLER_0_133_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11314_ _06283_ _06284_ _06285_ _06286_ vssd1 vssd1 vccd1 vccd1 _06287_ sky130_fd_sc_hd__or4_1
XFILLER_0_121_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15082_ net2609 net147 _01561_ net2306 vssd1 vssd1 vccd1 vccd1 _00408_ sky130_fd_sc_hd__a22o_1
XFILLER_0_121_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12294_ _07262_ vssd1 vssd1 vccd1 vccd1 img_gen.updater.update.next\[1\] sky130_fd_sc_hd__inv_2
XANTENNA__15522__B2 ag2.body\[534\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14033_ net986 ag2.body\[498\] vssd1 vssd1 vccd1 vccd1 _08194_ sky130_fd_sc_hd__or2_1
X_18910_ clknet_leaf_3_clk img_gen.tracker.next_frame\[348\] net1258 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[348\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_103_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11245_ ag2.body\[192\] net1233 vssd1 vssd1 vccd1 vccd1 _06218_ sky130_fd_sc_hd__nand2_1
XFILLER_0_121_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19890_ clknet_leaf_85_clk _00834_ net1463 vssd1 vssd1 vccd1 vccd1 ag2.body\[496\]
+ sky130_fd_sc_hd__dfrtp_4
XPHY_EDGE_ROW_20_Right_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11544__C1 net1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18841_ clknet_leaf_5_clk img_gen.tracker.next_frame\[279\] net1277 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[279\] sky130_fd_sc_hd__dfrtp_1
X_11176_ net1148 control.body\[779\] vssd1 vssd1 vccd1 vccd1 _06149_ sky130_fd_sc_hd__xor2_1
XFILLER_0_98_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10127_ net1193 control.body\[705\] vssd1 vssd1 vccd1 vccd1 _05100_ sky130_fd_sc_hd__xor2_1
XFILLER_0_59_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18772_ clknet_leaf_16_clk img_gen.tracker.next_frame\[210\] net1321 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[210\] sky130_fd_sc_hd__dfrtp_1
X_15984_ ag2.body\[2\] _08119_ vssd1 vssd1 vccd1 vccd1 _01668_ sky130_fd_sc_hd__or2_1
XANTENNA__09504__A2 net1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17723_ net461 _03401_ _01743_ vssd1 vssd1 vccd1 vccd1 _03402_ sky130_fd_sc_hd__a21o_1
XANTENNA__20094__RESET_B net1492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10058_ ag2.body\[481\] net1208 vssd1 vssd1 vccd1 vccd1 _05031_ sky130_fd_sc_hd__xor2_1
X_14935_ net2468 net167 _01544_ control.body\[1052\] vssd1 vssd1 vccd1 vccd1 _00278_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_19_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_236 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13425__A _07567_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17654_ _03327_ _03328_ _03330_ _03332_ vssd1 vssd1 vccd1 vccd1 _03333_ sky130_fd_sc_hd__or4b_2
X_14866_ net742 net59 vssd1 vssd1 vccd1 vccd1 _01536_ sky130_fd_sc_hd__nor2_1
XFILLER_0_76_1397 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1239 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10768__B net1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16605_ obsg2.obstacleArray\[83\] net451 net392 _02283_ vssd1 vssd1 vccd1 vccd1 _02284_
+ sky130_fd_sc_hd__o211a_1
X_13817_ control.detect2.Q\[1\] control.detect2.Q\[0\] vssd1 vssd1 vccd1 vccd1 _08114_
+ sky130_fd_sc_hd__nand2b_2
X_17585_ ag2.body\[56\] net738 net698 ag2.body\[62\] vssd1 vssd1 vccd1 vccd1 _03264_
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_54_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14797_ net823 ag2.body\[291\] _04097_ net1030 _01467_ vssd1 vssd1 vccd1 vccd1 _01468_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_57_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13064__A2 _07723_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19324_ clknet_leaf_103_clk _00268_ net1433 vssd1 vssd1 vccd1 vccd1 control.body\[1066\]
+ sky130_fd_sc_hd__dfrtp_1
X_16536_ net538 _02204_ vssd1 vssd1 vccd1 vccd1 _02215_ sky130_fd_sc_hd__nand2_1
X_13748_ img_gen.updater.commands.count\[1\] img_gen.updater.commands.count\[0\] _08061_
+ img_gen.updater.commands.count\[2\] vssd1 vssd1 vccd1 vccd1 _08067_ sky130_fd_sc_hd__a31o_1
XFILLER_0_46_818 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17735__C1 _03413_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19255_ clknet_leaf_75_clk _00199_ net1483 vssd1 vssd1 vccd1 vccd1 ag2.body\[118\]
+ sky130_fd_sc_hd__dfrtp_4
X_16467_ net403 _02143_ net366 vssd1 vssd1 vccd1 vccd1 _02146_ sky130_fd_sc_hd__o21a_1
XFILLER_0_116_706 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14013__A1 net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10784__A net1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14013__B2 net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13679_ _04641_ _08022_ net434 net911 vssd1 vssd1 vccd1 vccd1 track.nextCurrScore\[3\]
+ sky130_fd_sc_hd__a22o_1
X_18206_ _03649_ net36 vssd1 vssd1 vccd1 vccd1 _03742_ sky130_fd_sc_hd__nor2_1
X_15418_ control.body\[625\] net84 _01598_ ag2.body\[617\] vssd1 vssd1 vccd1 vccd1
+ _00707_ sky130_fd_sc_hd__a22o_1
X_19186_ clknet_leaf_53_clk _00130_ net1365 vssd1 vssd1 vccd1 vccd1 ag2.body\[49\]
+ sky130_fd_sc_hd__dfrtp_4
X_16398_ obsg2.obstacleArray\[106\] obsg2.obstacleArray\[107\] net454 vssd1 vssd1
+ vccd1 vccd1 _02077_ sky130_fd_sc_hd__mux2_1
XANTENNA__11378__A2 _04695_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18137_ net530 _03707_ vssd1 vssd1 vccd1 vccd1 _01316_ sky130_fd_sc_hd__and2_1
XFILLER_0_87_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15349_ net2283 net71 _01591_ control.body\[683\] vssd1 vssd1 vccd1 vccd1 _00645_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_13_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10586__B1 _04494_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_130_4273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold104 img_gen.tracker.frame\[7\] vssd1 vssd1 vccd1 vccd1 net1666 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_130_4284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold115 img_gen.tracker.frame\[281\] vssd1 vssd1 vccd1 vccd1 net1677 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_130_4295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18068_ obsg2.obstacleArray\[42\] _03661_ net520 vssd1 vssd1 vccd1 vccd1 _01293_
+ sky130_fd_sc_hd__o21a_1
XANTENNA__17286__B net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold126 img_gen.tracker.frame\[484\] vssd1 vssd1 vccd1 vccd1 net1688 sky130_fd_sc_hd__dlygate4sd3_1
Xhold137 img_gen.tracker.frame\[493\] vssd1 vssd1 vccd1 vccd1 net1699 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10008__B net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18767__CLK clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold148 img_gen.tracker.frame\[114\] vssd1 vssd1 vccd1 vccd1 net1710 sky130_fd_sc_hd__dlygate4sd3_1
X_09910_ ag2.body\[129\] net1211 vssd1 vssd1 vccd1 vccd1 _04883_ sky130_fd_sc_hd__xor2_1
X_17019_ ag2.body\[331\] net856 vssd1 vssd1 vccd1 vccd1 _02698_ sky130_fd_sc_hd__xor2_1
Xhold159 img_gen.tracker.frame\[383\] vssd1 vssd1 vccd1 vccd1 net1721 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19206__RESET_B net1461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12878__A2 _07425_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout606 net607 vssd1 vssd1 vccd1 vccd1 net606 sky130_fd_sc_hd__clkbuf_4
X_20030_ clknet_leaf_67_clk _00974_ net1472 vssd1 vssd1 vccd1 vccd1 ag2.body\[364\]
+ sky130_fd_sc_hd__dfrtp_4
Xfanout617 net620 vssd1 vssd1 vccd1 vccd1 net617 sky130_fd_sc_hd__clkbuf_4
X_09841_ net1083 control.body\[926\] vssd1 vssd1 vccd1 vccd1 _04814_ sky130_fd_sc_hd__nand2_1
XANTENNA__09743__A2 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout628 _06473_ vssd1 vssd1 vccd1 vccd1 net628 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_96_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout639 net640 vssd1 vssd1 vccd1 vccd1 net639 sky130_fd_sc_hd__buf_4
X_09772_ ag2.body\[239\] net1061 vssd1 vssd1 vccd1 vccd1 _04745_ sky130_fd_sc_hd__nand2_1
XANTENNA__16410__S net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18215__B1 net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_4099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15029__B1 _01555_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout277_A net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17569__A2 net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18230__A3 net37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16777__B1 net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20614__1557 vssd1 vssd1 vccd1 vccd1 net1557 _20614__1557/LO sky130_fd_sc_hd__conb_1
XANTENNA__15821__Y _01643_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13054__B _07720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout444_A net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13055__A2 _07720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1186_A net1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16365__B net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout611_A _06475_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout232_X net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1353_A net1355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout709_A net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15201__B1 _01574_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09206_ net1118 vssd1 vssd1 vccd1 vccd1 _04231_ sky130_fd_sc_hd__inv_2
XANTENNA__19542__CLK clknet_leaf_115_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12566__A1 net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09137_ ag2.body\[460\] vssd1 vssd1 vccd1 vccd1 _04162_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout1141_X net1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09068_ ag2.body\[274\] vssd1 vssd1 vccd1 vccd1 _04093_ sky130_fd_sc_hd__inv_2
XANTENNA__16701__B1 net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_113_3770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17196__B net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout980_A net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_3781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout699_X net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14613__B ag2.body\[56\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold660 control.body\[709\] vssd1 vssd1 vccd1 vccd1 net2222 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10329__B1 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09707__B net1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11526__C1 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout92_A net100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold671 toggle1.bcd_tens\[0\] vssd1 vssd1 vccd1 vccd1 net2233 sky130_fd_sc_hd__dlygate4sd3_1
Xhold682 control.body\[668\] vssd1 vssd1 vccd1 vccd1 net2244 sky130_fd_sc_hd__dlygate4sd3_1
X_11030_ net1135 control.body\[1044\] vssd1 vssd1 vccd1 vccd1 _06003_ sky130_fd_sc_hd__nand2_1
X_20228_ clknet_leaf_66_clk _01172_ net1476 vssd1 vssd1 vccd1 vccd1 ag2.body\[162\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__09734__A2 net1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold693 control.body\[658\] vssd1 vssd1 vccd1 vccd1 net2255 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout866_X net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20159_ clknet_leaf_96_clk _01103_ net1441 vssd1 vssd1 vccd1 vccd1 ag2.body\[237\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__18101__A net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16480__A2 _02059_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12981_ net668 _07686_ vssd1 vssd1 vccd1 vccd1 _07687_ sky130_fd_sc_hd__nor2_1
XANTENNA__10869__A ag2.body\[534\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14491__A1 net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_3574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14491__B2 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_3585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14720_ net1041 _04120_ _04121_ net1024 _08875_ vssd1 vssd1 vccd1 vccd1 _08881_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_107_3596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11932_ img_gen.tracker.frame\[172\] net603 vssd1 vssd1 vccd1 vccd1 _06904_ sky130_fd_sc_hd__or2_1
XFILLER_0_73_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18582__RESET_B net1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14651_ net1004 ag2.body\[144\] vssd1 vssd1 vccd1 vccd1 _08812_ sky130_fd_sc_hd__xor2_1
X_11863_ img_gen.tracker.frame\[193\] net624 vssd1 vssd1 vccd1 vccd1 _06835_ sky130_fd_sc_hd__or2_1
XFILLER_0_39_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13602_ control.divider.count\[19\] _07950_ _07975_ _07976_ vssd1 vssd1 vccd1 vccd1
+ _07977_ sky130_fd_sc_hd__o211a_1
X_10814_ _05783_ _05784_ _05785_ _05786_ _05782_ vssd1 vssd1 vccd1 vccd1 _05787_ sky130_fd_sc_hd__a221o_1
X_17370_ _03020_ _03048_ _03031_ vssd1 vssd1 vccd1 vccd1 _03049_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_67_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14582_ _08739_ _08740_ _08741_ _08742_ vssd1 vssd1 vccd1 vccd1 _08743_ sky130_fd_sc_hd__or4b_1
X_11794_ img_gen.tracker.frame\[371\] net587 net549 img_gen.tracker.frame\[368\] _06765_
+ vssd1 vssd1 vccd1 vccd1 _06766_ sky130_fd_sc_hd__o221a_1
XFILLER_0_28_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_2781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10100__C net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16321_ net416 _01997_ _01999_ net371 vssd1 vssd1 vccd1 vccd1 _02000_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_81_2792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13251__Y _07813_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10745_ ag2.body\[499\] net1162 vssd1 vssd1 vccd1 vccd1 _05718_ sky130_fd_sc_hd__xor2_1
X_13533_ net226 _07923_ _07924_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[566\]
+ sky130_fd_sc_hd__o21bai_1
XFILLER_0_83_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19040_ clknet_leaf_6_clk img_gen.tracker.next_frame\[478\] net1267 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[478\] sky130_fd_sc_hd__dfrtp_1
X_16252_ obsg2.obstacleArray\[62\] obsg2.obstacleArray\[63\] net407 vssd1 vssd1 vccd1
+ vccd1 _01931_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10280__A2 _04446_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13464_ net281 _07896_ _07897_ net1626 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[524\]
+ sky130_fd_sc_hd__a22o_1
X_10676_ ag2.body\[346\] net1185 vssd1 vssd1 vccd1 vccd1 _05649_ sky130_fd_sc_hd__xor2_1
XFILLER_0_42_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16940__B1 net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_990 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15203_ net2611 net94 _01574_ control.body\[810\] vssd1 vssd1 vccd1 vccd1 _00516_
+ sky130_fd_sc_hd__a22o_1
X_12415_ net480 _07171_ _07302_ vssd1 vssd1 vccd1 vccd1 _07377_ sky130_fd_sc_hd__and3b_1
XFILLER_0_106_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16183_ net346 _01861_ _01858_ _01742_ vssd1 vssd1 vccd1 vccd1 _01862_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_11_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13395_ net259 _07870_ _07871_ net1855 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[481\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__10109__A net1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10568__B1 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09457__X _04430_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15134_ net2614 net107 _01566_ control.body\[877\] vssd1 vssd1 vccd1 vccd1 _00455_
+ sky130_fd_sc_hd__a22o_1
X_12346_ net590 _06638_ net439 net565 vssd1 vssd1 vccd1 vccd1 _07313_ sky130_fd_sc_hd__or4_1
XFILLER_0_84_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11780__A2 net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19942_ clknet_leaf_46_clk _00886_ net1375 vssd1 vssd1 vccd1 vccd1 ag2.body\[452\]
+ sky130_fd_sc_hd__dfrtp_2
X_15065_ control.body\[951\] net149 _01559_ control.body\[943\] vssd1 vssd1 vccd1
+ vccd1 _00393_ sky130_fd_sc_hd__a22o_1
XFILLER_0_107_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_75_2596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12277_ _07196_ _07225_ _04274_ vssd1 vssd1 vccd1 vccd1 _07247_ sky130_fd_sc_hd__and3b_1
X_14016_ net1016 _04163_ _04164_ net1008 vssd1 vssd1 vccd1 vccd1 _08177_ sky130_fd_sc_hd__o22a_1
XFILLER_0_103_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11228_ _06199_ _06200_ vssd1 vssd1 vccd1 vccd1 _06201_ sky130_fd_sc_hd__nand2_1
X_19873_ clknet_leaf_94_clk _00817_ net1440 vssd1 vssd1 vccd1 vccd1 ag2.body\[527\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__09931__A_N net1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15259__B1 net50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17799__A2 net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18824_ clknet_leaf_2_clk img_gen.tracker.next_frame\[262\] net1249 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[262\] sky130_fd_sc_hd__dfrtp_1
X_11159_ ag2.body\[602\] net1169 vssd1 vssd1 vccd1 vccd1 _06132_ sky130_fd_sc_hd__xor2_1
XANTENNA__18011__A net45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12978__B net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15354__B net53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18755_ clknet_leaf_15_clk img_gen.tracker.next_frame\[193\] net1312 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[193\] sky130_fd_sc_hd__dfrtp_1
X_15967_ ag2.body\[138\] net213 _01658_ ag2.body\[130\] vssd1 vssd1 vccd1 vccd1 _01196_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__14482__A1 net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19415__CLK clknet_leaf_103_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13285__A2 _07827_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14482__B2 net1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17706_ _01895_ _02047_ _03384_ vssd1 vssd1 vccd1 vccd1 _03385_ sky130_fd_sc_hd__and3b_1
X_14918_ control.body\[1077\] net170 _01542_ net2221 vssd1 vssd1 vccd1 vccd1 _00263_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__16759__B1 net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18686_ clknet_leaf_28_clk img_gen.tracker.next_frame\[124\] net1335 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[124\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_91_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_1183 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15898_ ag2.body\[205\] net133 _01650_ ag2.body\[197\] vssd1 vssd1 vccd1 vccd1 _01135_
+ sky130_fd_sc_hd__a22o_1
X_17637_ _03312_ _03313_ _03314_ _03315_ _03311_ vssd1 vssd1 vccd1 vccd1 _03316_ sky130_fd_sc_hd__a221o_1
X_14849_ _01507_ _01508_ _01513_ _01519_ vssd1 vssd1 vccd1 vccd1 _01520_ sky130_fd_sc_hd__and4_1
XANTENNA__16466__A net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17568_ ag2.body\[583\] net688 net723 ag2.body\[578\] vssd1 vssd1 vccd1 vccd1 _03247_
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_85_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19307_ clknet_leaf_99_clk _00251_ net1445 vssd1 vssd1 vccd1 vccd1 control.body\[1081\]
+ sky130_fd_sc_hd__dfrtp_1
X_16519_ _02194_ _02197_ _02057_ vssd1 vssd1 vccd1 vccd1 _02198_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_74_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_136_4460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_4471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17499_ ag2.body\[232\] net885 vssd1 vssd1 vccd1 vccd1 _03178_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_136_4482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19238_ clknet_leaf_84_clk _00182_ net1481 vssd1 vssd1 vccd1 vccd1 ag2.body\[101\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__20542__CLK clknet_leaf_105_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_132_4335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_4346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_4357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_41_1563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19169_ clknet_leaf_52_clk _00113_ net1366 vssd1 vssd1 vccd1 vccd1 ag2.body\[32\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_41_1585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10559__B1 _04416_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11220__A1 _06180_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10961__B net1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_1442 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11771__A2 net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout403 _02063_ vssd1 vssd1 vccd1 vccd1 net403 sky130_fd_sc_hd__clkbuf_4
XANTENNA__13049__B _07718_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09716__A2 net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout414 _01901_ vssd1 vssd1 vccd1 vccd1 net414 sky130_fd_sc_hd__clkbuf_2
Xfanout425 _01735_ vssd1 vssd1 vccd1 vccd1 net425 sky130_fd_sc_hd__buf_2
XFILLER_0_22_1436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_54_1957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout394_A net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout436 net437 vssd1 vssd1 vccd1 vccd1 net436 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_54_1968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20013_ clknet_leaf_59_clk _00957_ net1467 vssd1 vssd1 vccd1 vccd1 ag2.body\[379\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_54_1979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout447 net448 vssd1 vssd1 vccd1 vccd1 net447 sky130_fd_sc_hd__clkbuf_4
X_09824_ net1058 control.body\[927\] vssd1 vssd1 vccd1 vccd1 _04797_ sky130_fd_sc_hd__nand2_1
Xfanout458 net459 vssd1 vssd1 vccd1 vccd1 net458 sky130_fd_sc_hd__buf_4
XANTENNA_fanout1101_A net1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_1389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout469 _06648_ vssd1 vssd1 vccd1 vccd1 net469 sky130_fd_sc_hd__buf_2
XANTENNA__09543__A net1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15264__B net54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09755_ _04724_ _04725_ _04726_ _04727_ vssd1 vssd1 vccd1 vccd1 _04728_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout182_X net182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout561_A net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout659_A _04394_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13065__A net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11137__X _06110_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17760__A net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09686_ ag2.body\[9\] net1198 vssd1 vssd1 vccd1 vccd1 _04659_ sky130_fd_sc_hd__xor2_1
XFILLER_0_69_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20072__CLK clknet_leaf_73_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1470_A net1478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10201__B net1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1091_X net1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout826_A net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout447_X net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14225__B2 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1189_X net1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15973__A1 net223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12787__A1 net239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout43 net44 vssd1 vssd1 vccd1 vccd1 net43 sky130_fd_sc_hd__buf_2
XFILLER_0_92_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1010 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18932__CLK clknet_leaf_141_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout54 net55 vssd1 vssd1 vccd1 vccd1 net54 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout1356_X net1356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12409__A net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout65 net67 vssd1 vssd1 vccd1 vccd1 net65 sky130_fd_sc_hd__clkbuf_4
XANTENNA__17714__A2 net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout76 net79 vssd1 vssd1 vccd1 vccd1 net76 sky130_fd_sc_hd__clkbuf_2
X_10530_ net1109 control.body\[917\] vssd1 vssd1 vccd1 vccd1 _05503_ sky130_fd_sc_hd__or2_1
XFILLER_0_49_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout87 net89 vssd1 vssd1 vccd1 vccd1 net87 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_98_3297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout98 net100 vssd1 vssd1 vccd1 vccd1 net98 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_115_3821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17919__B net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19199__RESET_B net1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_115_3832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16823__B net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12128__B net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_115_3843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13465__A_N net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10461_ _05430_ _05431_ _05432_ _05433_ vssd1 vssd1 vccd1 vccd1 _05434_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_21_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14624__A net1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_3707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12200_ net480 _07171_ vssd1 vssd1 vccd1 vccd1 _07172_ sky130_fd_sc_hd__or2_1
XANTENNA__11747__C1 net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_3718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11967__B net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13180_ net341 net332 _07515_ vssd1 vssd1 vccd1 vccd1 _07781_ sky130_fd_sc_hd__or3b_1
XANTENNA_clkbuf_3_0_0_clk_X clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10392_ net1181 control.body\[1058\] vssd1 vssd1 vccd1 vccd1 _05365_ sky130_fd_sc_hd__xor2_1
XFILLER_0_62_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout983_X net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19195__Q ag2.body\[58\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12131_ img_gen.tracker.frame\[561\] net588 net549 img_gen.tracker.frame\[558\] vssd1
+ vssd1 vccd1 vccd1 _07103_ sky130_fd_sc_hd__o22a_1
XANTENNA__11762__A2 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17935__A net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09437__B net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11686__C net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12062_ img_gen.tracker.frame\[69\] net593 net554 img_gen.tracker.frame\[66\] _07033_
+ vssd1 vssd1 vccd1 vccd1 _07034_ sky130_fd_sc_hd__a221o_1
Xhold490 img_gen.tracker.frame\[70\] vssd1 vssd1 vccd1 vccd1 net2052 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_19_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11514__A2 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12711__A1 net237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11013_ ag2.body\[592\] net1220 vssd1 vssd1 vccd1 vccd1 _05986_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_70_2460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_3636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_2471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_3647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16870_ ag2.body\[470\] net939 vssd1 vssd1 vccd1 vccd1 _02549_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_109_3658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16989__B1 net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout970 net971 vssd1 vssd1 vccd1 vccd1 net970 sky130_fd_sc_hd__buf_4
Xfanout981 net982 vssd1 vssd1 vccd1 vccd1 net981 sky130_fd_sc_hd__clkbuf_8
XANTENNA__20511__D track.nextHighScore\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15821_ _04986_ net59 vssd1 vssd1 vccd1 vccd1 _01643_ sky130_fd_sc_hd__nor2_4
Xfanout992 net995 vssd1 vssd1 vccd1 vccd1 net992 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_5_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18540_ clknet_leaf_135_clk _00066_ net1298 vssd1 vssd1 vccd1 vccd1 img_gen.updater.commands.count\[9\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_35_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15752_ ag2.body\[330\] net216 _01635_ ag2.body\[322\] vssd1 vssd1 vccd1 vccd1 _01004_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_73_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19588__CLK clknet_leaf_118_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12964_ net668 _07678_ vssd1 vssd1 vccd1 vccd1 _07679_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_87_2990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14703_ net1001 ag2.body\[232\] vssd1 vssd1 vccd1 vccd1 _08864_ sky130_fd_sc_hd__xor2_1
X_18471_ _03956_ vssd1 vssd1 vccd1 vccd1 _03957_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_83_2843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11915_ img_gen.tracker.frame\[355\] net542 _06885_ _06886_ vssd1 vssd1 vccd1 vccd1
+ _06887_ sky130_fd_sc_hd__o211a_1
XANTENNA__11207__B _05254_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14216__A1 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15683_ ag2.body\[397\] net142 _01627_ ag2.body\[389\] vssd1 vssd1 vccd1 vccd1 _00943_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_115_1622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_83_2854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14216__B2 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_83_2865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12895_ net292 _07645_ _07646_ net1691 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[206\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_129_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17422_ ag2.body\[113\] net876 vssd1 vssd1 vccd1 vccd1 _03101_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_64_2264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20565__CLK clknet_leaf_43_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14634_ net817 ag2.body\[579\] ag2.body\[581\] net806 vssd1 vssd1 vccd1 vccd1 _08795_
+ sky130_fd_sc_hd__a22o_1
X_11846_ img_gen.tracker.frame\[515\] net583 net544 img_gen.tracker.frame\[512\] _06817_
+ vssd1 vssd1 vccd1 vccd1 _06818_ sky130_fd_sc_hd__o221a_1
XFILLER_0_51_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_2275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_2286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_2139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17353_ net1044 net1043 ag2.body\[2\] vssd1 vssd1 vccd1 vccd1 _03032_ sky130_fd_sc_hd__or3_1
X_14565_ net1040 ag2.body\[356\] vssd1 vssd1 vccd1 vccd1 _08726_ sky130_fd_sc_hd__xor2_1
X_11777_ img_gen.tracker.frame\[164\] net548 vssd1 vssd1 vccd1 vccd1 _06749_ sky130_fd_sc_hd__or2_1
XANTENNA__17705__A2 net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09643__B2 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16304_ obsg2.obstacleArray\[101\] net413 vssd1 vssd1 vccd1 vccd1 _01983_ sky130_fd_sc_hd__or2_1
XFILLER_0_3_1452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11223__A net1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13516_ net2121 net656 _07917_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[556\]
+ sky130_fd_sc_hd__and3_1
X_10728_ net1159 ag2.body\[251\] vssd1 vssd1 vccd1 vccd1 _05701_ sky130_fd_sc_hd__nand2b_1
X_17284_ ag2.body\[307\] net856 vssd1 vssd1 vccd1 vccd1 _02963_ sky130_fd_sc_hd__xor2_1
XFILLER_0_82_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_856 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14496_ net1039 ag2.body\[260\] vssd1 vssd1 vccd1 vccd1 _08657_ sky130_fd_sc_hd__xor2_1
XANTENNA__16913__B1 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19023_ clknet_leaf_2_clk img_gen.tracker.next_frame\[461\] net1247 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[461\] sky130_fd_sc_hd__dfrtp_1
X_16235_ obsg2.obstacleArray\[34\] obsg2.obstacleArray\[35\] net404 vssd1 vssd1 vccd1
+ vccd1 _01914_ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10659_ _05624_ _05625_ _05628_ _05631_ vssd1 vssd1 vccd1 vccd1 _05632_ sky130_fd_sc_hd__or4_4
X_13447_ net235 _07890_ _07891_ net1960 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[513\]
+ sky130_fd_sc_hd__a22o_1
Xclkload13 clknet_leaf_144_clk vssd1 vssd1 vccd1 vccd1 clkload13/X sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_77_2658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload24 clknet_leaf_14_clk vssd1 vssd1 vccd1 vccd1 clkload24/Y sky130_fd_sc_hd__clkinv_4
XTAP_TAPCELL_ROW_77_2669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload35 clknet_leaf_141_clk vssd1 vssd1 vccd1 vccd1 clkload35/X sky130_fd_sc_hd__clkbuf_8
XANTENNA__12980__C _07638_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload46 clknet_leaf_28_clk vssd1 vssd1 vccd1 vccd1 clkload46/Y sky130_fd_sc_hd__bufinv_16
XFILLER_0_45_1403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__20456__RESET_B net1355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16166_ net349 _01840_ _01844_ _01743_ vssd1 vssd1 vccd1 vccd1 _01845_ sky130_fd_sc_hd__o211a_1
X_13378_ net670 _07864_ vssd1 vssd1 vccd1 vccd1 _07865_ sky130_fd_sc_hd__nor2_1
XANTENNA__17469__B2 ag2.body\[534\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload57 clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 clkload57/Y sky130_fd_sc_hd__clkinv_8
Xclkload68 clknet_leaf_44_clk vssd1 vssd1 vccd1 vccd1 clkload68/Y sky130_fd_sc_hd__inv_4
XTAP_TAPCELL_ROW_58_2079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16677__C1 _02211_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload79 clknet_leaf_121_clk vssd1 vssd1 vccd1 vccd1 clkload79/Y sky130_fd_sc_hd__inv_8
XANTENNA__11753__A2 net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15117_ control.body\[902\] net146 _01554_ control.body\[894\] vssd1 vssd1 vccd1
+ vccd1 _00440_ sky130_fd_sc_hd__a22o_1
X_12329_ _07251_ _07253_ vssd1 vssd1 vccd1 vccd1 _07296_ sky130_fd_sc_hd__nor2_1
X_20613__1556 vssd1 vssd1 vccd1 vccd1 net1556 _20613__1556/LO sky130_fd_sc_hd__conb_1
X_16097_ _01742_ _01771_ _01775_ _01729_ vssd1 vssd1 vccd1 vccd1 _01776_ sky130_fd_sc_hd__a31o_1
XANTENNA__12054__A net1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19925_ clknet_leaf_51_clk _00869_ net1368 vssd1 vssd1 vccd1 vccd1 ag2.body\[467\]
+ sky130_fd_sc_hd__dfrtp_4
X_15048_ _06413_ net59 vssd1 vssd1 vccd1 vccd1 _01558_ sky130_fd_sc_hd__nor2_2
XANTENNA__17564__B net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09634__Y _04607_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19856_ clknet_leaf_92_clk _00800_ net1412 vssd1 vssd1 vccd1 vccd1 ag2.body\[542\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_125_4150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10713__B1 _05685_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17641__A1 ag2.body\[160\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_4003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15084__B net58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18807_ clknet_leaf_3_clk img_gen.tracker.next_frame\[245\] net1258 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[245\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__17641__B2 ag2.body\[166\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19787_ clknet_leaf_127_clk _00731_ net1328 vssd1 vssd1 vccd1 vccd1 ag2.body\[601\]
+ sky130_fd_sc_hd__dfrtp_4
X_16999_ _02674_ _02675_ _02676_ _02677_ vssd1 vssd1 vccd1 vccd1 _02678_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_121_4025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09540_ net1059 control.body\[1031\] vssd1 vssd1 vccd1 vccd1 _04513_ sky130_fd_sc_hd__nand2_1
X_18738_ clknet_leaf_141_clk img_gen.tracker.next_frame\[176\] net1261 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[176\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_30_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10302__A net1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_1419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09471_ _04440_ _04443_ vssd1 vssd1 vccd1 vccd1 _04444_ sky130_fd_sc_hd__or2_1
XFILLER_0_8_1330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18669_ clknet_leaf_10_clk img_gen.tracker.next_frame\[107\] net1273 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[107\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__15812__B net66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09882__A1 ag2.body\[160\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10021__B net1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18955__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_4522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09882__B2 ag2.body\[164\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15404__B1 _01581_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_4533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_138_4566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10956__B net1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_134_4408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20631_ net1548 vssd1 vssd1 vccd1 vccd1 gpio_out[26] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_134_4419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13332__B _07505_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_28_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17157__B1 net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_968 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_823 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11133__A net1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_1647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_15_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20562_ clknet_leaf_109_clk toggle1.nextDisplayOut\[2\] net1421 vssd1 vssd1 vccd1
+ vccd1 ssdec1.in\[2\] sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_24_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload7 clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 clkload7/X sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_24_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_24_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_1249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20493_ clknet_leaf_21_clk _01380_ net1360 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[129\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_15_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10972__A net1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout407_A net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19221__RESET_B net1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1051_A net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14444__A net1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_3150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13194__A1 net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_3161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1149_A net1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_3172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20197__RESET_B net1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11744__A2 net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16132__A1 _01743_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17755__A _03045_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1316_A net1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout200 net218 vssd1 vssd1 vccd1 vccd1 net200 sky130_fd_sc_hd__clkbuf_2
XANTENNA__17474__B net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout211 net214 vssd1 vssd1 vccd1 vccd1 net211 sky130_fd_sc_hd__buf_2
Xfanout1209 net1213 vssd1 vssd1 vccd1 vccd1 net1209 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout397_X net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout776_A _04229_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout222 net223 vssd1 vssd1 vccd1 vccd1 net222 sky130_fd_sc_hd__clkbuf_2
Xfanout233 net247 vssd1 vssd1 vccd1 vccd1 net233 sky130_fd_sc_hd__buf_2
Xfanout244 net247 vssd1 vssd1 vccd1 vccd1 net244 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout1104_X net1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout255 net257 vssd1 vssd1 vccd1 vccd1 net255 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_103_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout266 net269 vssd1 vssd1 vccd1 vccd1 net266 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09570__B1 net1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17632__A1 ag2.body\[161\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09807_ _04773_ _04774_ _04779_ _04772_ vssd1 vssd1 vccd1 vccd1 _04780_ sky130_fd_sc_hd__or4b_1
Xfanout277 net278 vssd1 vssd1 vccd1 vccd1 net277 sky130_fd_sc_hd__clkbuf_4
Xfanout288 net295 vssd1 vssd1 vccd1 vccd1 net288 sky130_fd_sc_hd__buf_2
Xfanout299 _03546_ vssd1 vssd1 vccd1 vccd1 net299 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout943_A obsg2.randCord\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout564_X net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15643__B1 _01623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_3500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09738_ _04704_ _04710_ _04698_ vssd1 vssd1 vccd1 vccd1 _04711_ sky130_fd_sc_hd__or3b_2
XANTENNA__17921__C _03554_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1632 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout55_A net62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1138 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15722__B _01631_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16199__A1 net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout731_X net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17396__B1 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09669_ net639 _04640_ vssd1 vssd1 vccd1 vccd1 _04642_ sky130_fd_sc_hd__nand2b_4
XANTENNA__09873__A1 _04822_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout829_X net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12472__A3 _07306_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1210 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09873__B2 _04845_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11700_ _06642_ _06670_ vssd1 vssd1 vccd1 vccd1 _06672_ sky130_fd_sc_hd__xor2_4
XFILLER_0_35_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1232 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_367 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12680_ net589 _06639_ net435 net563 vssd1 vssd1 vccd1 vccd1 _07545_ sky130_fd_sc_hd__or4_1
XANTENNA__09720__B _04688_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11631_ obsg2.obstacleArray\[34\] net510 net506 _06603_ vssd1 vssd1 vccd1 vccd1 _06604_
+ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_13_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_117_3905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09625__A1 _04587_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_834 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14350_ net1018 ag2.body\[406\] vssd1 vssd1 vccd1 vccd1 _08511_ sky130_fd_sc_hd__or2_1
X_11562_ net505 _06533_ _06534_ net759 vssd1 vssd1 vccd1 vccd1 _06535_ sky130_fd_sc_hd__a211o_1
XANTENNA__19110__CLK clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17649__B net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_1625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_1585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10513_ ag2.body\[100\] net1140 vssd1 vssd1 vccd1 vccd1 _05486_ sky130_fd_sc_hd__xnor2_1
XANTENNA__11983__A2 net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13301_ net256 _07833_ _07834_ net1610 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[424\]
+ sky130_fd_sc_hd__a22o_1
X_14281_ net1003 _04036_ ag2.body\[141\] net809 vssd1 vssd1 vccd1 vccd1 _08442_ sky130_fd_sc_hd__a22o_1
X_11493_ net1102 net1222 vssd1 vssd1 vccd1 vccd1 _06466_ sky130_fd_sc_hd__and2b_1
XFILLER_0_24_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14354__A net1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_174 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16020_ _01695_ _01697_ vssd1 vssd1 vccd1 vccd1 _01699_ sky130_fd_sc_hd__xnor2_2
X_13232_ net232 _07426_ _07805_ net1791 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[384\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11697__B net1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10444_ net1158 control.body\[931\] vssd1 vssd1 vccd1 vccd1 _05417_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_122_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19260__CLK clknet_leaf_73_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_2511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11735__A2 net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13163_ net327 _07505_ _07638_ vssd1 vssd1 vccd1 vccd1 _07773_ sky130_fd_sc_hd__and3_1
XANTENNA__16123__A1 net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10375_ ag2.body\[111\] net1066 vssd1 vssd1 vccd1 vccd1 _05348_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_72_2522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_2533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10943__B1 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12114_ net1215 net1190 img_gen.tracker.frame\[165\] vssd1 vssd1 vccd1 vccd1 _07086_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_27_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18828__CLK clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17971_ net380 _01713_ net481 vssd1 vssd1 vccd1 vccd1 _03594_ sky130_fd_sc_hd__and3_1
XANTENNA__17384__B net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13094_ net387 _07460_ _07638_ vssd1 vssd1 vccd1 vccd1 _07740_ sky130_fd_sc_hd__and3_1
XANTENNA__14685__A1 net1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14685__B2 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19710_ clknet_leaf_134_clk _00654_ net1307 vssd1 vssd1 vccd1 vccd1 control.body\[684\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__17952__X _03579_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12045_ img_gen.tracker.frame\[249\] net593 net554 img_gen.tracker.frame\[246\] _07016_
+ vssd1 vssd1 vccd1 vccd1 _07017_ sky130_fd_sc_hd__a221o_1
X_16922_ _02595_ _02600_ vssd1 vssd1 vccd1 vccd1 _02601_ sky130_fd_sc_hd__nand2b_1
XANTENNA__12602__A _07431_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12160__A2 net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19641_ clknet_leaf_123_clk _00585_ net1406 vssd1 vssd1 vccd1 vccd1 control.body\[759\]
+ sky130_fd_sc_hd__dfrtp_1
X_16853_ ag2.body\[174\] net696 _02520_ _02521_ _02531_ vssd1 vssd1 vccd1 vccd1 _02532_
+ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_85_2905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15804_ ag2.body\[280\] net206 _01641_ ag2.body\[272\] vssd1 vssd1 vccd1 vccd1 _01050_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11218__A net1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19572_ clknet_leaf_116_clk _00516_ net1387 vssd1 vssd1 vccd1 vccd1 control.body\[818\]
+ sky130_fd_sc_hd__dfrtp_1
X_16784_ net462 _02425_ _02436_ net352 vssd1 vssd1 vccd1 vccd1 _02463_ sky130_fd_sc_hd__o211a_1
XFILLER_0_88_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10122__A net1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_2326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13996_ ag2.body\[132\] net213 _08160_ ag2.body\[124\] vssd1 vssd1 vccd1 vccd1 _00213_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__14842__D1 _01512_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_66_2337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18523_ clknet_leaf_135_clk img_gen.updater.update.next\[0\] net1299 vssd1 vssd1
+ vccd1 vccd1 img_gen.updater.commands.mode\[0\] sky130_fd_sc_hd__dfrtp_2
XANTENNA__15191__Y _01573_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_2348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15632__B net64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15735_ ag2.body\[347\] net211 _01633_ ag2.body\[339\] vssd1 vssd1 vccd1 vccd1 _00989_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_1_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12947_ net685 _07670_ vssd1 vssd1 vccd1 vccd1 _07671_ sky130_fd_sc_hd__nor2_1
XANTENNA__17387__B1 net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14529__A net1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18454_ _04642_ _03823_ _03841_ _03942_ vssd1 vssd1 vccd1 vccd1 _03943_ sky130_fd_sc_hd__a211o_1
X_15666_ ag2.body\[414\] net143 _01625_ ag2.body\[406\] vssd1 vssd1 vccd1 vccd1 _00928_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__15937__B2 ag2.body\[167\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12878_ net245 _07425_ _07638_ _07640_ net1854 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[195\]
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_28_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10776__B net1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17405_ ag2.body\[42\] net722 net715 ag2.body\[43\] _03082_ vssd1 vssd1 vccd1 vccd1
+ _03084_ sky130_fd_sc_hd__a221o_1
X_14617_ net817 ag2.body\[59\] _03998_ net1006 vssd1 vssd1 vccd1 vccd1 _08778_ sky130_fd_sc_hd__o22a_1
X_18385_ _03793_ _03805_ vssd1 vssd1 vccd1 vccd1 _03875_ sky130_fd_sc_hd__nor2_1
X_11829_ net385 _06800_ vssd1 vssd1 vccd1 vccd1 _06801_ sky130_fd_sc_hd__nand2_1
X_15597_ _04447_ net57 vssd1 vssd1 vccd1 vccd1 _01619_ sky130_fd_sc_hd__nor2_2
XFILLER_0_5_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17336_ net924 net696 vssd1 vssd1 vccd1 vccd1 _03015_ sky130_fd_sc_hd__and2_1
XFILLER_0_16_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14548_ net1020 ag2.body\[246\] vssd1 vssd1 vccd1 vccd1 _08709_ sky130_fd_sc_hd__xor2_1
XPHY_EDGE_ROW_112_Right_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17267_ _04081_ net863 net707 ag2.body\[253\] _02945_ vssd1 vssd1 vccd1 vccd1 _02946_
+ sky130_fd_sc_hd__o221a_1
X_14479_ net989 ag2.body\[441\] vssd1 vssd1 vccd1 vccd1 _08640_ sky130_fd_sc_hd__xor2_1
XFILLER_0_109_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14264__A net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload102 clknet_leaf_100_clk vssd1 vssd1 vccd1 vccd1 clkload102/Y sky130_fd_sc_hd__bufinv_16
XFILLER_0_125_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkload113 clknet_leaf_60_clk vssd1 vssd1 vccd1 vccd1 clkload113/Y sky130_fd_sc_hd__bufinv_16
XFILLER_0_11_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13176__A1 net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19006_ clknet_leaf_0_clk img_gen.tracker.next_frame\[444\] net1245 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[444\] sky130_fd_sc_hd__dfrtp_1
X_16218_ net503 _01889_ vssd1 vssd1 vccd1 vccd1 _01897_ sky130_fd_sc_hd__nor2_1
Xclkload124 clknet_leaf_82_clk vssd1 vssd1 vccd1 vccd1 clkload124/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_10_1181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09919__A2 net1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17198_ ag2.body\[178\] net861 vssd1 vssd1 vccd1 vccd1 _02877_ sky130_fd_sc_hd__or2_1
XANTENNA__11187__B1 net1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_49_Right_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11400__B net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16149_ obsg2.obstacleArray\[21\] net431 vssd1 vssd1 vccd1 vccd1 _01828_ sky130_fd_sc_hd__or2_1
XANTENNA__17311__B1 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14551__X _08712_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_127_4201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09645__X _04618_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16665__A2 net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17294__B net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08971_ ag2.body\[60\] vssd1 vssd1 vccd1 vccd1 _03996_ sky130_fd_sc_hd__inv_2
XANTENNA__10016__B net1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19908_ clknet_leaf_54_clk _00852_ net1457 vssd1 vssd1 vccd1 vccd1 ag2.body\[482\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_97_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold19 score_detect.N\[0\] vssd1 vssd1 vccd1 vccd1 net1581 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12512__A net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12151__A2 net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19839_ clknet_leaf_92_clk _00783_ net1414 vssd1 vssd1 vccd1 vccd1 ag2.body\[557\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__14428__A1 net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15625__B1 _01621_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14428__B2 net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1638 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_58_Right_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_49_1812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09523_ net1171 control.body\[834\] vssd1 vssd1 vccd1 vccd1 _04496_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_49_1823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09855__A1 net1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10967__A net1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09855__B2 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_879 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13343__A net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1099_A net1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09454_ net900 net905 vssd1 vssd1 vccd1 vccd1 _04427_ sky130_fd_sc_hd__and2_4
XFILLER_0_56_1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11662__A1 net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10686__B net1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_26_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13062__B net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09385_ sound_gen.osc1.stayCount\[11\] _04355_ vssd1 vssd1 vccd1 vccd1 _04377_ sky130_fd_sc_hd__nor2_1
XFILLER_0_30_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout524_A net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14600__A1 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_540 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14600__B2 net1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20614_ net1557 vssd1 vssd1 vccd1 vccd1 gpio_oeb[26] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_95_3212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20378__RESET_B net1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_3223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_3234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16373__B net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_1013 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19283__CLK clknet_leaf_98_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11965__A2 net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20307__RESET_B net1499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20545_ clknet_leaf_105_clk _01410_ _00019_ vssd1 vssd1 vccd1 vccd1 sound_gen.osc1.stayCount\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_61_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16353__A1 obsg2.obstacleArray\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14174__A net1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_140_clk clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_140_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_127_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_91_3109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1054_X net1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_314 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13167__A1 net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_67_Right_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20476_ clknet_leaf_38_clk _01363_ net1354 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[112\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_15_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout893_A net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_144 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__20260__CLK clknet_leaf_43_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12406__B net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16105__A1 net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11310__B net1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_1610 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1221_X net1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_520 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10160_ net910 _04571_ net643 vssd1 vssd1 vccd1 vccd1 _05133_ sky130_fd_sc_hd__o21ai_2
XANTENNA_fanout681_X net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_89_3027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_89_3038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1006 net1007 vssd1 vssd1 vccd1 vccd1 net1006 sky130_fd_sc_hd__buf_4
XANTENNA_fanout779_X net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_89_3049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1017 net1018 vssd1 vssd1 vccd1 vccd1 net1017 sky130_fd_sc_hd__buf_2
X_10091_ net1148 control.body\[795\] vssd1 vssd1 vccd1 vccd1 _05064_ sky130_fd_sc_hd__nand2_1
Xfanout1028 net1029 vssd1 vssd1 vccd1 vccd1 net1028 sky130_fd_sc_hd__buf_4
XFILLER_0_22_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1039 net1042 vssd1 vssd1 vccd1 vccd1 net1039 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_22_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12142__A2 net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17932__B _03531_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13237__B _07425_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout946_X net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_76_Right_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13850_ ag2.body\[14\] net127 _08133_ net1577 vssd1 vssd1 vccd1 vccd1 _00094_ sky130_fd_sc_hd__a22o_1
XFILLER_0_88_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout58_X net58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12801_ net328 _07444_ _07505_ vssd1 vssd1 vccd1 vccd1 _07603_ sky130_fd_sc_hd__and3_1
XANTENNA__10299__D _05271_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15452__B net63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10993_ ag2.body\[340\] net1141 vssd1 vssd1 vccd1 vccd1 _05966_ sky130_fd_sc_hd__xor2_1
X_13781_ _08090_ _08070_ vssd1 vssd1 vccd1 vccd1 _00068_ sky130_fd_sc_hd__and2b_1
XFILLER_0_134_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14349__A net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11102__B1 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1462 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15520_ ag2.body\[540\] net156 _01609_ ag2.body\[532\] vssd1 vssd1 vccd1 vccd1 _00798_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__13253__A _07443_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12732_ net388 _07444_ _07460_ vssd1 vssd1 vccd1 vccd1 _07570_ sky130_fd_sc_hd__and3_1
XANTENNA__09450__B net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20612__1544 vssd1 vssd1 vccd1 vccd1 _20612__1544/HI net1544 sky130_fd_sc_hd__conb_1
XFILLER_0_97_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_52_clk_A clknet_4_6__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15451_ ag2.body\[607\] net86 _01601_ ag2.body\[599\] vssd1 vssd1 vccd1 vccd1 _00737_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_2_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12663_ net680 _07536_ vssd1 vssd1 vccd1 vccd1 _07537_ sky130_fd_sc_hd__nor2_1
XFILLER_0_38_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14402_ net990 net1043 vssd1 vssd1 vccd1 vccd1 _08563_ sky130_fd_sc_hd__xor2_1
X_11614_ net504 _06586_ vssd1 vssd1 vccd1 vccd1 _06587_ sky130_fd_sc_hd__or2_1
X_18170_ _03606_ _03706_ vssd1 vssd1 vccd1 vccd1 _03724_ sky130_fd_sc_hd__nor2_1
XANTENNA__17379__B net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15382_ net2590 net87 _01595_ net2302 vssd1 vssd1 vccd1 vccd1 _00674_ sky130_fd_sc_hd__a22o_1
X_12594_ net327 _07497_ vssd1 vssd1 vccd1 vccd1 _07498_ sky130_fd_sc_hd__or2_2
XFILLER_0_25_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10883__Y _05856_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18333__A2 net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_85_Right_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18379__B1_N track.nextHighScore\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17121_ _02793_ _02794_ _02799_ _02792_ vssd1 vssd1 vccd1 vccd1 _02800_ sky130_fd_sc_hd__or4b_1
X_14333_ net981 _04151_ ag2.body\[429\] net807 _08491_ vssd1 vssd1 vccd1 vccd1 _08494_
+ sky130_fd_sc_hd__a221o_1
X_11545_ net505 _06516_ _06517_ net475 vssd1 vssd1 vccd1 vccd1 _06518_ sky130_fd_sc_hd__o31a_1
XANTENNA_clkbuf_leaf_67_clk_A clknet_4_13__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17541__B1 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1206 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_131_clk clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_131_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_0_1466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_2130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11501__A net1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17052_ _02726_ _02727_ _02728_ _02730_ vssd1 vssd1 vccd1 vccd1 _02731_ sky130_fd_sc_hd__or4_1
XFILLER_0_80_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14264_ net989 ag2.body\[9\] vssd1 vssd1 vccd1 vccd1 _08425_ sky130_fd_sc_hd__or2_1
X_11476_ ag2.body\[493\] net1114 vssd1 vssd1 vccd1 vccd1 _06449_ sky130_fd_sc_hd__nand2_1
Xwire475 _06484_ vssd1 vssd1 vccd1 vccd1 net475 sky130_fd_sc_hd__buf_4
XANTENNA_clkbuf_leaf_110_clk_A clknet_4_10__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_55_2005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16003_ net539 _01681_ _01679_ vssd1 vssd1 vccd1 vccd1 _01682_ sky130_fd_sc_hd__a21o_2
XANTENNA__11708__A2 net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13215_ net240 _07796_ _07797_ net1782 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[375\]
+ sky130_fd_sc_hd__a22o_1
X_10427_ net1060 control.body\[1071\] vssd1 vssd1 vccd1 vccd1 _05400_ sky130_fd_sc_hd__or2_1
X_14195_ net792 ag2.body\[167\] ag2.body\[162\] net827 vssd1 vssd1 vccd1 vccd1 _08356_
+ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__10117__A net1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10358_ net1187 ag2.body\[290\] vssd1 vssd1 vccd1 vccd1 _05331_ sky130_fd_sc_hd__and2b_1
X_13146_ net667 _07764_ vssd1 vssd1 vccd1 vccd1 _07765_ sky130_fd_sc_hd__nor2_1
XFILLER_0_46_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19006__CLK clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17954_ obsg2.obstacleArray\[9\] _03580_ net529 vssd1 vssd1 vccd1 vccd1 _01260_ sky130_fd_sc_hd__o21a_1
X_13077_ net685 _07731_ vssd1 vssd1 vccd1 vccd1 _07732_ sky130_fd_sc_hd__nor2_1
X_10289_ ag2.body\[330\] net1186 vssd1 vssd1 vccd1 vccd1 _05262_ sky130_fd_sc_hd__or2_1
XANTENNA_clkbuf_leaf_125_clk_A clknet_4_9__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_94_Right_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_29_Left_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13330__A1 net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20322__Q obsg2.randCord\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12028_ _06993_ _06999_ net470 vssd1 vssd1 vccd1 vccd1 _07000_ sky130_fd_sc_hd__mux2_1
X_16905_ ag2.body\[243\] net854 vssd1 vssd1 vccd1 vccd1 _02584_ sky130_fd_sc_hd__xor2_1
X_17885_ net920 _04239_ obsg2.obstacleCount\[0\] vssd1 vssd1 vccd1 vccd1 _03525_ sky130_fd_sc_hd__a21bo_1
XANTENNA__11341__B1 _04686_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15607__B1 _01620_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_4_2__f_clk_X clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16836_ ag2.body\[99\] net853 vssd1 vssd1 vccd1 vccd1 _02515_ sky130_fd_sc_hd__xor2_1
X_19624_ clknet_leaf_119_clk _00568_ net1392 vssd1 vssd1 vccd1 vccd1 control.body\[774\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19555_ clknet_leaf_115_clk _00499_ net1397 vssd1 vssd1 vccd1 vccd1 control.body\[833\]
+ sky130_fd_sc_hd__dfrtp_1
X_16767_ _02443_ _02445_ net497 vssd1 vssd1 vccd1 vccd1 _02446_ sky130_fd_sc_hd__mux2_1
X_13979_ ag2.body\[117\] net203 _08158_ ag2.body\[109\] vssd1 vssd1 vccd1 vccd1 _00198_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__10787__A net1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18506_ net1517 net1511 vssd1 vssd1 vccd1 vccd1 _00037_ sky130_fd_sc_hd__or2_1
XFILLER_0_57_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15718_ ag2.body\[365\] net193 _01630_ ag2.body\[357\] vssd1 vssd1 vccd1 vccd1 _00975_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_17_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19486_ clknet_leaf_114_clk _00430_ net1400 vssd1 vssd1 vccd1 vccd1 control.body\[908\]
+ sky130_fd_sc_hd__dfrtp_1
X_16698_ obsg2.obstacleArray\[71\] net502 net493 obsg2.obstacleArray\[68\] _02376_
+ vssd1 vssd1 vccd1 vccd1 _02377_ sky130_fd_sc_hd__a221o_1
XFILLER_0_18_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18437_ _03923_ _03924_ _03925_ vssd1 vssd1 vccd1 vccd1 _03926_ sky130_fd_sc_hd__a21oi_1
X_15649_ ag2.body\[431\] net138 _01623_ ag2.body\[423\] vssd1 vssd1 vccd1 vccd1 _00913_
+ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_1_Left_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17780__B1 _03458_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_38_Left_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09170_ ag2.body\[531\] vssd1 vssd1 vccd1 vccd1 _04195_ sky130_fd_sc_hd__inv_2
XFILLER_0_90_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18368_ _07181_ _03819_ _03861_ _08024_ vssd1 vssd1 vccd1 vccd1 _03862_ sky130_fd_sc_hd__o31a_1
XFILLER_0_5_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16193__B net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11947__A2 net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17319_ ag2.body\[223\] net932 vssd1 vssd1 vccd1 vccd1 _02998_ sky130_fd_sc_hd__xor2_1
X_18299_ net323 net321 _03782_ _03793_ vssd1 vssd1 vccd1 vccd1 _03795_ sky130_fd_sc_hd__a31o_1
XFILLER_0_43_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_122_clk clknet_4_9__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_122_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_43_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12507__A net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13149__A1 net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20330_ clknet_leaf_108_clk sound_gen.osc1.freq_nxt\[2\] _00006_ vssd1 vssd1 vccd1
+ vccd1 sound_gen.osc1.freq\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_71_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20261_ clknet_leaf_43_clk _01205_ net1379 vssd1 vssd1 vccd1 vccd1 ag2.body\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_64_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout105_A net107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12372__A2 net241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09816__A net1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20192_ clknet_leaf_88_clk _01136_ net1459 vssd1 vssd1 vccd1 vccd1 ag2.body\[206\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_12_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_47_Left_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15846__B1 _01644_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13338__A net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08954_ ag2.body\[14\] vssd1 vssd1 vccd1 vccd1 _03979_ sky130_fd_sc_hd__inv_2
XANTENNA__09535__B net1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20232__Q ag2.body\[166\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12124__A2 net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17752__B _02928_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13872__A2 net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout474_A _06647_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12896__B net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16368__B _01918_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09551__A net1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10697__A _04470_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12388__S net1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout262_X net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout641_A _04419_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1383_A net1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout739_A net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09506_ _04146_ net1088 net1065 _04147_ _04478_ vssd1 vssd1 vccd1 vccd1 _04479_ sky130_fd_sc_hd__a221o_1
XFILLER_0_91_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11635__A1 net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_56_Left_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09437_ ag2.body\[7\] net1055 vssd1 vssd1 vccd1 vccd1 _04410_ sky130_fd_sc_hd__nand2_1
XANTENNA__11305__B net1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout527_X net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17771__B1 _03175_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1171_X net1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout906_A net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13801__A net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09368_ _03959_ _04369_ _04351_ net273 vssd1 vssd1 vccd1 vccd1 _01420_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_35_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14616__B ag2.body\[60\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11938__A2 net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17767__X _03446_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20141__RESET_B net1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_113_clk clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_113_clk
+ sky130_fd_sc_hd__clkbuf_8
X_09299_ sound_gen.osc1.keepCounting_nxt _04318_ vssd1 vssd1 vccd1 vccd1 _04319_ sky130_fd_sc_hd__and2_2
XFILLER_0_7_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15129__A2 net107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17523__B1 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12417__A net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_13__f_clk_X clknet_4_13__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1398 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11330_ net1095 control.body\[661\] vssd1 vssd1 vccd1 vccd1 _06303_ sky130_fd_sc_hd__or2_1
X_20528_ clknet_leaf_114_clk _01393_ net1398 vssd1 vssd1 vccd1 vccd1 toggle1.bcd_tens\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_62_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11261_ net753 control.body\[773\] control.body\[775\] net743 vssd1 vssd1 vccd1 vccd1
+ _06234_ sky130_fd_sc_hd__a22o_1
X_20459_ clknet_leaf_38_clk _01346_ net1354 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[95\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_28_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10212_ _05181_ _05182_ _05183_ _05184_ vssd1 vssd1 vccd1 vccd1 _05185_ sky130_fd_sc_hd__a22o_1
X_13000_ img_gen.tracker.frame\[262\] net645 vssd1 vssd1 vccd1 vccd1 _07696_ sky130_fd_sc_hd__and2_1
XFILLER_0_105_1440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11192_ net1151 control.body\[875\] vssd1 vssd1 vccd1 vccd1 _06165_ sky130_fd_sc_hd__nand2_1
XANTENNA__10374__A1 net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10143_ net1099 control.body\[821\] vssd1 vssd1 vccd1 vccd1 _05116_ sky130_fd_sc_hd__or2_1
XFILLER_0_101_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_1237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19179__CLK clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12115__A2 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17662__B net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10074_ _05041_ _05042_ _05043_ _05044_ _05045_ vssd1 vssd1 vccd1 vccd1 _05047_ sky130_fd_sc_hd__a221o_1
X_14951_ net2327 net166 _01546_ control.body\[1034\] vssd1 vssd1 vccd1 vccd1 _00292_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_27_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17054__A2 net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13902_ ag2.body\[48\] net118 _08150_ ag2.body\[40\] vssd1 vssd1 vccd1 vccd1 _00129_
+ sky130_fd_sc_hd__a22o_1
X_17670_ ag2.body\[453\] net950 vssd1 vssd1 vccd1 vccd1 _03349_ sky130_fd_sc_hd__xor2_1
X_14882_ control.body\[1109\] net177 _01538_ control.body\[1101\] vssd1 vssd1 vccd1
+ vccd1 _00231_ sky130_fd_sc_hd__a22o_1
XANTENNA_hold739_X net2301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16621_ _02297_ _02298_ _02299_ net394 net359 vssd1 vssd1 vccd1 vccd1 _02300_ sky130_fd_sc_hd__a221o_1
X_13833_ net1628 net662 _08128_ _08127_ vssd1 vssd1 vccd1 vccd1 _00082_ sky130_fd_sc_hd__a31o_1
XANTENNA__15182__B net53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14079__A net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11055__X _06028_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14812__B2 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19340_ clknet_leaf_103_clk _00284_ net1431 vssd1 vssd1 vccd1 vccd1 control.body\[1050\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_43_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16552_ obsg2.obstacleArray\[100\] obsg2.obstacleArray\[101\] net441 vssd1 vssd1
+ vccd1 vccd1 _02231_ sky130_fd_sc_hd__mux2_1
X_13764_ img_gen.updater.commands.count\[6\] _08077_ vssd1 vssd1 vccd1 vccd1 _08079_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_6_1620 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10976_ _05939_ _05940_ _05944_ _05945_ _05948_ vssd1 vssd1 vccd1 vccd1 _05949_ sky130_fd_sc_hd__o221a_1
XFILLER_0_134_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16014__B1 net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15503_ ag2.body\[557\] net113 _01607_ ag2.body\[549\] vssd1 vssd1 vccd1 vccd1 _00783_
+ sky130_fd_sc_hd__a22o_1
X_19271_ clknet_leaf_71_clk _00215_ net1503 vssd1 vssd1 vccd1 vccd1 ag2.body\[134\]
+ sky130_fd_sc_hd__dfrtp_4
X_12715_ net305 _07561_ vssd1 vssd1 vccd1 vccd1 _07562_ sky130_fd_sc_hd__nor2_1
XFILLER_0_6_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16483_ obsg2.obstacleArray\[44\] net452 vssd1 vssd1 vccd1 vccd1 _02162_ sky130_fd_sc_hd__or2_1
XFILLER_0_31_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14229__D net1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15910__B net54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13695_ track.current_collision net464 _08036_ vssd1 vssd1 vccd1 vccd1 _08037_ sky130_fd_sc_hd__and3_1
XANTENNA__17762__B1 _03110_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18222_ _03664_ net36 vssd1 vssd1 vccd1 vccd1 _03750_ sky130_fd_sc_hd__nor2_1
XFILLER_0_2_1517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15434_ _05287_ net52 vssd1 vssd1 vccd1 vccd1 _01600_ sky130_fd_sc_hd__nor2_2
XFILLER_0_72_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12646_ net438 net472 net563 net555 vssd1 vssd1 vccd1 vccd1 _07526_ sky130_fd_sc_hd__and4_1
XFILLER_0_26_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_1620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18153_ net523 _03715_ vssd1 vssd1 vccd1 vccd1 _01324_ sky130_fd_sc_hd__and2_1
XANTENNA__13430__B _07460_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16317__A1 _01912_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15365_ net2574 net68 _01593_ net2234 vssd1 vssd1 vccd1 vccd1 _00659_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_104_clk clknet_4_10__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_104_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_109_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17514__B1 net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12577_ net247 _07488_ _07489_ net1663 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[45\]
+ sky130_fd_sc_hd__a22o_1
X_17104_ ag2.body\[13\] net948 vssd1 vssd1 vccd1 vccd1 _02783_ sky130_fd_sc_hd__xor2_1
XANTENNA__20317__Q ag2.randCord\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14316_ net988 _03991_ ag2.body\[50\] net824 _08476_ vssd1 vssd1 vccd1 vccd1 _08477_
+ sky130_fd_sc_hd__a221o_1
X_11528_ net504 _06499_ _06500_ net475 vssd1 vssd1 vccd1 vccd1 _06501_ sky130_fd_sc_hd__o31a_1
X_18084_ net352 _03539_ net38 obsg2.obstacleArray\[48\] vssd1 vssd1 vccd1 vccd1 _03672_
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_80_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15296_ net2450 net76 _01585_ control.body\[732\] vssd1 vssd1 vccd1 vccd1 _00598_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold308 img_gen.tracker.frame\[290\] vssd1 vssd1 vccd1 vccd1 net1870 sky130_fd_sc_hd__dlygate4sd3_1
X_17035_ ag2.body\[122\] net866 vssd1 vssd1 vccd1 vccd1 _02714_ sky130_fd_sc_hd__xnor2_1
Xhold319 img_gen.tracker.frame\[231\] vssd1 vssd1 vccd1 vccd1 net1881 sky130_fd_sc_hd__dlygate4sd3_1
X_14247_ net837 ag2.body\[537\] ag2.body\[540\] net814 vssd1 vssd1 vccd1 vccd1 _08408_
+ sky130_fd_sc_hd__a2bb2o_1
X_11459_ ag2.body\[258\] net1187 vssd1 vssd1 vccd1 vccd1 _06432_ sky130_fd_sc_hd__or2_1
XFILLER_0_0_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14542__A net1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18014__A net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09636__A net1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11885__B net1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14178_ net841 ag2.body\[192\] _04060_ net988 vssd1 vssd1 vccd1 vccd1 _08339_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_81_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15828__B1 _01643_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13158__A net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13129_ net243 _07755_ _07756_ net1647 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[330\]
+ sky130_fd_sc_hd__a22o_1
X_18986_ clknet_leaf_8_clk img_gen.tracker.next_frame\[424\] net1271 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[424\] sky130_fd_sc_hd__dfrtp_1
Xhold1008 control.body\[734\] vssd1 vssd1 vccd1 vccd1 net2570 sky130_fd_sc_hd__dlygate4sd3_1
X_17937_ net318 _03567_ obsg2.obstacleArray\[5\] vssd1 vssd1 vccd1 vccd1 _03568_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_59_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1019 control.body\[920\] vssd1 vssd1 vccd1 vccd1 net2581 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12997__A net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13308__D _07486_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1624 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1370 net1505 vssd1 vssd1 vccd1 vccd1 net1370 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_108_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1381 net1382 vssd1 vssd1 vccd1 vccd1 net1381 sky130_fd_sc_hd__clkbuf_4
X_17868_ _03503_ _03514_ vssd1 vssd1 vccd1 vccd1 _01240_ sky130_fd_sc_hd__nor2_1
XANTENNA__11865__A1 net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1392 net1395 vssd1 vssd1 vccd1 vccd1 net1392 sky130_fd_sc_hd__buf_2
XFILLER_0_108_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19607_ clknet_leaf_119_clk _00551_ net1393 vssd1 vssd1 vccd1 vccd1 control.body\[789\]
+ sky130_fd_sc_hd__dfrtp_1
X_16819_ ag2.body\[81\] net734 net701 ag2.body\[86\] _02493_ vssd1 vssd1 vccd1 vccd1
+ _02498_ sky130_fd_sc_hd__o221a_1
XANTENNA__14820__A1_N net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17799_ net969 net957 net948 vssd1 vssd1 vccd1 vccd1 _03471_ sky130_fd_sc_hd__a21o_1
XFILLER_0_117_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14803__A1 net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14803__B2 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1490 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19538_ clknet_leaf_115_clk _00482_ net1397 vssd1 vssd1 vccd1 vccd1 control.body\[848\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_49_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_1463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19469_ clknet_leaf_112_clk _00413_ net1424 vssd1 vssd1 vccd1 vccd1 control.body\[923\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14276__X _08437_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14717__A net1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09222_ control.body\[893\] vssd1 vssd1 vccd1 vccd1 _04247_ sky130_fd_sc_hd__inv_2
XFILLER_0_130_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09153_ ag2.body\[492\] vssd1 vssd1 vccd1 vccd1 _04178_ sky130_fd_sc_hd__inv_2
XFILLER_0_99_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout222_A net223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkload110_A clknet_leaf_88_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17505__B1 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20227__Q ag2.body\[161\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09084_ ag2.body\[320\] vssd1 vssd1 vccd1 vccd1 _04109_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_1163 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20313_ clknet_leaf_44_clk _01213_ net1380 vssd1 vssd1 vccd1 vccd1 ag2.randCord\[7\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_102_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17984__C_N net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold820 control.body\[760\] vssd1 vssd1 vccd1 vccd1 net2382 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10980__A net1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1131_A net1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold831 control.body\[1102\] vssd1 vssd1 vccd1 vccd1 net2393 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold842 control.body\[924\] vssd1 vssd1 vccd1 vccd1 net2404 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1229_A net1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20244_ clknet_leaf_69_clk _01188_ net1496 vssd1 vssd1 vccd1 vccd1 ag2.body\[146\]
+ sky130_fd_sc_hd__dfrtp_4
Xhold853 obsg2.obsNeeded\[2\] vssd1 vssd1 vccd1 vccd1 net2415 sky130_fd_sc_hd__dlygate4sd3_1
Xhold864 control.body\[931\] vssd1 vssd1 vccd1 vccd1 net2426 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10356__A1 ag2.body\[291\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold875 control.body\[1037\] vssd1 vssd1 vccd1 vccd1 net2437 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout591_A net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20611__1543 vssd1 vssd1 vccd1 vccd1 _20611__1543/HI net1543 sky130_fd_sc_hd__conb_1
XFILLER_0_101_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold886 _00539_ vssd1 vssd1 vccd1 vccd1 net2448 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout689_A net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold897 control.body\[955\] vssd1 vssd1 vccd1 vccd1 net2459 sky130_fd_sc_hd__dlygate4sd3_1
X_20175_ clknet_leaf_82_clk _01119_ net1479 vssd1 vssd1 vccd1 vccd1 ag2.body\[221\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_110_681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09986_ net1086 control.body\[1118\] vssd1 vssd1 vccd1 vccd1 _04959_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout1017_X net1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19835__RESET_B net1414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08937_ ag2.goodColl vssd1 vssd1 vccd1 vccd1 _03962_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout856_A net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16379__A net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13845__A2 net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10698__Y _05671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16795__A1 _02075_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout644_X net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_64_Left_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1386_X net1386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10830_ _05799_ _05800_ _05801_ _05802_ vssd1 vssd1 vccd1 vccd1 _05803_ sky130_fd_sc_hd__or4_1
XANTENNA__20393__RESET_B net1355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_120_3978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_120_3989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16826__B net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16547__A1 net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout811_X net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10761_ net756 control.body\[893\] _04248_ net1083 _05733_ vssd1 vssd1 vccd1 vccd1
+ _05734_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_101_3399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14627__A net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16318__S net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17744__B1 _03286_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12500_ _07443_ net306 vssd1 vssd1 vccd1 vccd1 _07446_ sky130_fd_sc_hd__or2_1
XANTENNA__14558__B1 ag2.body\[71\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10692_ ag2.body\[144\] net788 net1113 _04043_ _05662_ vssd1 vssd1 vccd1 vccd1 _05665_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_109_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13480_ net308 _07598_ vssd1 vssd1 vccd1 vccd1 _07904_ sky130_fd_sc_hd__nor2_1
XANTENNA__19198__Q ag2.body\[61\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10874__B net1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12431_ _07391_ _07392_ vssd1 vssd1 vccd1 vccd1 _07393_ sky130_fd_sc_hd__nor2_1
XFILLER_0_63_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15150_ net2433 net99 _01568_ control.body\[859\] vssd1 vssd1 vccd1 vccd1 _00469_
+ sky130_fd_sc_hd__a22o_1
X_12362_ _07282_ _07283_ _07300_ _07328_ vssd1 vssd1 vccd1 vccd1 net10 sky130_fd_sc_hd__a22o_1
XFILLER_0_23_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17657__B net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_73_Left_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14101_ net1026 ag2.body\[589\] vssd1 vssd1 vccd1 vccd1 _08262_ sky130_fd_sc_hd__xor2_1
X_11313_ ag2.body\[273\] net1207 vssd1 vssd1 vccd1 vccd1 _06286_ sky130_fd_sc_hd__xor2_1
X_15081_ control.body\[933\] net148 _01561_ net2281 vssd1 vssd1 vccd1 vccd1 _00407_
+ sky130_fd_sc_hd__a22o_1
X_12293_ _07220_ _07260_ _07261_ _04388_ img_gen.updater.commands.mode\[2\] vssd1
+ vssd1 vccd1 vccd1 _07262_ sky130_fd_sc_hd__a32o_1
XANTENNA__14362__A net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_1550 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_957 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13533__A1 net226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14032_ net986 ag2.body\[498\] vssd1 vssd1 vccd1 vccd1 _08193_ sky130_fd_sc_hd__nand2_1
X_11244_ ag2.body\[192\] net1233 vssd1 vssd1 vccd1 vccd1 _06217_ sky130_fd_sc_hd__or2_1
XANTENNA__09456__A _04416_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_1594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18569__CLK clknet_leaf_15_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18472__A1 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11175_ net1075 control.body\[782\] vssd1 vssd1 vccd1 vccd1 _06148_ sky130_fd_sc_hd__xor2_1
X_18840_ clknet_leaf_14_clk img_gen.tracker.next_frame\[278\] net1276 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[278\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_101_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_1608 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10126_ net1148 control.body\[707\] vssd1 vssd1 vccd1 vccd1 _05099_ sky130_fd_sc_hd__xor2_1
XANTENNA__17392__B net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18771_ clknet_leaf_19_clk img_gen.tracker.next_frame\[209\] net1321 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[209\] sky130_fd_sc_hd__dfrtp_1
X_15983_ _01663_ _01665_ vssd1 vssd1 vccd1 vccd1 _01667_ sky130_fd_sc_hd__nand2b_1
XANTENNA__19505__RESET_B net1404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17027__A2 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17722_ obsg2.obstacleArray\[132\] obsg2.obstacleArray\[133\] obsg2.obstacleArray\[134\]
+ obsg2.obstacleArray\[135\] net427 net378 vssd1 vssd1 vccd1 vccd1 _03401_ sky130_fd_sc_hd__mux4_1
X_10057_ _05027_ _05028_ _05029_ vssd1 vssd1 vccd1 vccd1 _05030_ sky130_fd_sc_hd__a21o_1
X_14934_ net2319 net173 _01544_ control.body\[1051\] vssd1 vssd1 vccd1 vccd1 _00277_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_136_1208 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_82_Left_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_19_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17653_ _03324_ _03325_ _03331_ vssd1 vssd1 vccd1 vccd1 _03332_ sky130_fd_sc_hd__and3_1
XFILLER_0_37_1316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_248 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14865_ _03962_ ag2.appleSet _01535_ vssd1 vssd1 vccd1 vccd1 _00217_ sky130_fd_sc_hd__a21o_1
XANTENNA__16786__B2 net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17983__B1 net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkload0_A clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16604_ obsg2.obstacleArray\[82\] net447 vssd1 vssd1 vccd1 vccd1 _02283_ sky130_fd_sc_hd__or2_1
XFILLER_0_37_1349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13816_ control.detect1.Q\[1\] control.detect1.Q\[0\] vssd1 vssd1 vccd1 vccd1 _08113_
+ sky130_fd_sc_hd__and2b_2
X_17584_ ag2.body\[56\] net738 obsg2.randCord\[1\] _03995_ vssd1 vssd1 vccd1 vccd1
+ _03263_ sky130_fd_sc_hd__a22o_1
XFILLER_0_98_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14796_ net838 ag2.body\[289\] ag2.body\[293\] net809 vssd1 vssd1 vccd1 vccd1 _01467_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_97_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19323_ clknet_leaf_100_clk _00267_ net1444 vssd1 vssd1 vccd1 vccd1 control.body\[1065\]
+ sky130_fd_sc_hd__dfrtp_1
X_16535_ _01733_ _02204_ vssd1 vssd1 vccd1 vccd1 _02214_ sky130_fd_sc_hd__nand2_2
XFILLER_0_15_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11075__A2 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13747_ _07189_ _08065_ _08066_ net320 net2476 vssd1 vssd1 vccd1 vccd1 _00058_ sky130_fd_sc_hd__a32o_1
X_10959_ _05928_ _05929_ _05930_ _05931_ vssd1 vssd1 vccd1 vccd1 _05932_ sky130_fd_sc_hd__a22o_1
XANTENNA__17735__B1 _03412_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18009__A net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13441__A net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19254_ clknet_leaf_75_clk _00198_ net1492 vssd1 vssd1 vccd1 vccd1 ag2.body\[117\]
+ sky130_fd_sc_hd__dfrtp_4
X_16466_ net397 _02144_ vssd1 vssd1 vccd1 vccd1 _02145_ sky130_fd_sc_hd__or2_1
XFILLER_0_112_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13678_ _04638_ _08022_ net434 net915 vssd1 vssd1 vccd1 vccd1 track.nextCurrScore\[2\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_116_718 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18205_ obsg2.obstacleArray\[99\] _03741_ net521 vssd1 vssd1 vccd1 vccd1 _01350_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_128_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13160__B net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15417_ net2654 net81 _01598_ ag2.body\[616\] vssd1 vssd1 vccd1 vccd1 _00706_ sky130_fd_sc_hd__a22o_1
X_19185_ clknet_leaf_53_clk _00129_ net1366 vssd1 vssd1 vccd1 vccd1 ag2.body\[48\]
+ sky130_fd_sc_hd__dfrtp_4
X_12629_ net2052 net644 _07516_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[70\]
+ sky130_fd_sc_hd__and3_1
X_16397_ net463 _02065_ vssd1 vssd1 vccd1 vccd1 _02076_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_109_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_91_Left_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18136_ _03542_ net298 net37 obsg2.obstacleArray\[65\] vssd1 vssd1 vccd1 vccd1 _03707_
+ sky130_fd_sc_hd__a31o_1
X_15348_ net2628 net71 _01591_ control.body\[682\] vssd1 vssd1 vccd1 vccd1 _00644_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__10586__A1 _04425_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11783__B1 net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_130_4274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11896__A net1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_130_4285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18067_ net42 _03660_ vssd1 vssd1 vccd1 vccd1 _03661_ sky130_fd_sc_hd__nor2_1
Xhold105 img_gen.tracker.frame\[165\] vssd1 vssd1 vccd1 vccd1 net1667 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14272__A net1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold116 img_gen.tracker.frame\[147\] vssd1 vssd1 vccd1 vccd1 net1678 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15279_ net2381 net88 _01583_ control.body\[749\] vssd1 vssd1 vccd1 vccd1 _00583_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_130_4296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold127 img_gen.tracker.frame\[108\] vssd1 vssd1 vccd1 vccd1 net1689 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__20321__CLK clknet_leaf_43_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold138 img_gen.tracker.frame\[536\] vssd1 vssd1 vccd1 vccd1 net1700 sky130_fd_sc_hd__dlygate4sd3_1
X_17018_ _04114_ net877 net866 _04115_ _02696_ vssd1 vssd1 vccd1 vccd1 _02697_ sky130_fd_sc_hd__a221o_1
XFILLER_0_112_968 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold149 img_gen.tracker.frame\[289\] vssd1 vssd1 vccd1 vccd1 net1711 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10008__C _04980_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19494__CLK clknet_leaf_113_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12878__A3 _07638_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18463__A1 net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09840_ net1083 control.body\[926\] vssd1 vssd1 vccd1 vccd1 _04813_ sky130_fd_sc_hd__or2_1
Xfanout607 net608 vssd1 vssd1 vccd1 vccd1 net607 sky130_fd_sc_hd__clkbuf_4
XANTENNA__17266__A2 net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout618 net620 vssd1 vssd1 vccd1 vccd1 net618 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_95_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10305__A net1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout629 _06473_ vssd1 vssd1 vccd1 vccd1 net629 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_0_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09771_ ag2.body\[233\] net1206 vssd1 vssd1 vccd1 vccd1 _04744_ sky130_fd_sc_hd__nand2_1
X_18969_ clknet_leaf_6_clk img_gen.tracker.next_frame\[407\] net1267 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[407\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__19246__RESET_B net1482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17018__A2 net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12520__A net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09900__B1 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10510__A1 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10510__B2 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1438 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10040__A net1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11493__A_N net1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1081_A net1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14447__A net992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1179_A net1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09205_ net1152 vssd1 vssd1 vccd1 vccd1 _04230_ sky130_fd_sc_hd__inv_4
XANTENNA_fanout604_A net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout225_X net225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1346_A net1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11369__A3 _06341_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09136_ ag2.body\[456\] vssd1 vssd1 vccd1 vccd1 _04161_ sky130_fd_sc_hd__inv_2
XFILLER_0_72_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14960__B1 _01547_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09067_ ag2.body\[271\] vssd1 vssd1 vccd1 vccd1 _04092_ sky130_fd_sc_hd__inv_2
XFILLER_0_5_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18711__CLK clknet_leaf_144_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_3760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09547__Y _04520_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15504__A2 net113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_113_3771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14182__A net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1134_X net1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_3782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09719__B1 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold650 img_gen.updater.commands.rR1.rainbowRNG\[10\] vssd1 vssd1 vccd1 vccd1 net2212
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10329__A1 net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout973_A net974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11526__B1 net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold661 control.body\[1021\] vssd1 vssd1 vccd1 vccd1 net2223 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout594_X net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold672 control.body\[665\] vssd1 vssd1 vccd1 vccd1 net2234 sky130_fd_sc_hd__dlygate4sd3_1
X_20227_ clknet_leaf_66_clk _01171_ net1476 vssd1 vssd1 vccd1 vccd1 ag2.body\[161\]
+ sky130_fd_sc_hd__dfrtp_4
Xhold683 control.body\[937\] vssd1 vssd1 vccd1 vccd1 net2245 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17257__A2 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold694 _00668_ vssd1 vssd1 vccd1 vccd1 net2256 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__17924__C net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout85_A net91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20158_ clknet_leaf_96_clk _01102_ net1441 vssd1 vssd1 vccd1 vccd1 ag2.body\[236\]
+ sky130_fd_sc_hd__dfrtp_4
X_09969_ _04938_ _04939_ _04940_ _04941_ vssd1 vssd1 vccd1 vccd1 _04942_ sky130_fd_sc_hd__or4_1
XANTENNA_fanout761_X net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout859_X net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20089_ clknet_leaf_77_clk _01033_ net1491 vssd1 vssd1 vccd1 vccd1 ag2.body\[311\]
+ sky130_fd_sc_hd__dfrtp_4
X_12980_ net332 _07505_ _07638_ vssd1 vssd1 vccd1 vccd1 _07686_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_107_3575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10869__B net1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_3586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11931_ net438 _06888_ _06889_ _06661_ vssd1 vssd1 vccd1 vccd1 _06903_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_107_3597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14650_ net977 ag2.body\[147\] vssd1 vssd1 vccd1 vccd1 _08811_ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout40_X net40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11862_ img_gen.tracker.frame\[202\] net591 net566 vssd1 vssd1 vccd1 vccd1 _06834_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_79_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13601_ control.divider.count\[19\] _07950_ _07949_ control.divider.count\[18\] vssd1
+ vssd1 vccd1 vccd1 _07976_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_67_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10813_ net1160 control.body\[1091\] vssd1 vssd1 vccd1 vccd1 _05786_ sky130_fd_sc_hd__or2_1
XFILLER_0_138_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14581_ net843 ag2.body\[488\] ag2.body\[489\] net833 vssd1 vssd1 vccd1 vccd1 _08742_
+ sky130_fd_sc_hd__o22a_1
X_11793_ img_gen.tracker.frame\[362\] net621 net605 img_gen.tracker.frame\[365\] vssd1
+ vssd1 vccd1 vccd1 _06765_ sky130_fd_sc_hd__o22a_1
XANTENNA__10885__A net1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_1550 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16320_ obsg2.obstacleArray\[69\] net414 _01998_ net420 vssd1 vssd1 vccd1 vccd1 _01999_
+ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_81_2782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13532_ img_gen.tracker.frame\[566\] net655 _07923_ vssd1 vssd1 vccd1 vccd1 _07924_
+ sky130_fd_sc_hd__and3_1
XANTENNA__19367__CLK clknet_leaf_93_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10744_ _05713_ _05714_ _05715_ _05716_ vssd1 vssd1 vccd1 vccd1 _05717_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_81_2793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20509__D ag2.goodColl vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_876 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16251_ _01929_ vssd1 vssd1 vccd1 vccd1 _01930_ sky130_fd_sc_hd__inv_2
XFILLER_0_125_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13463_ net256 _07896_ _07897_ net1673 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[523\]
+ sky130_fd_sc_hd__a22o_1
X_10675_ ag2.body\[350\] net1092 vssd1 vssd1 vccd1 vccd1 _05648_ sky130_fd_sc_hd__xor2_1
X_15202_ net2635 net92 _01574_ net2182 vssd1 vssd1 vccd1 vccd1 _00515_ sky130_fd_sc_hd__a22o_1
XFILLER_0_129_1034 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09738__X _04711_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12414_ _07282_ _07367_ _07376_ _07300_ vssd1 vssd1 vccd1 vccd1 net29 sky130_fd_sc_hd__a22o_1
XFILLER_0_35_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09958__B1 _04916_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16182_ _01859_ _01860_ net376 vssd1 vssd1 vccd1 vccd1 _01861_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_11_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14951__B1 _01546_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13394_ net238 _07870_ _07871_ net2015 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[480\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11765__B1 net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15133_ control.body\[884\] net114 _01566_ control.body\[876\] vssd1 vssd1 vccd1
+ vccd1 _00454_ sky130_fd_sc_hd__a22o_1
XANTENNA__18560__Q ag2.x\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12345_ _07306_ _07311_ vssd1 vssd1 vccd1 vccd1 _07312_ sky130_fd_sc_hd__nor2_2
XFILLER_0_65_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14092__A net1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19941_ clknet_leaf_46_clk _00885_ net1376 vssd1 vssd1 vccd1 vccd1 ag2.body\[451\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_107_1354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15064_ control.body\[950\] net149 _01559_ net2456 vssd1 vssd1 vccd1 vccd1 _00392_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_75_2597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12276_ _07242_ _07245_ vssd1 vssd1 vccd1 vccd1 _07246_ sky130_fd_sc_hd__nand2_1
XFILLER_0_120_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14015_ net999 _04161_ _04164_ net1008 _08175_ vssd1 vssd1 vccd1 vccd1 _08176_ sky130_fd_sc_hd__a221o_1
XFILLER_0_107_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11227_ net778 control.body\[857\] _04244_ net1171 vssd1 vssd1 vccd1 vccd1 _06200_
+ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__11612__S0 net1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19872_ clknet_leaf_95_clk _00816_ net1440 vssd1 vssd1 vccd1 vccd1 ag2.body\[526\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_120_1532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09473__X _04446_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18823_ clknet_leaf_2_clk img_gen.tracker.next_frame\[261\] net1250 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[261\] sky130_fd_sc_hd__dfrtp_1
X_11158_ ag2.body\[600\] net1219 vssd1 vssd1 vccd1 vccd1 _06131_ sky130_fd_sc_hd__xor2_1
XANTENNA__13436__A net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10109_ net1157 control.body\[939\] vssd1 vssd1 vccd1 vccd1 _05082_ sky130_fd_sc_hd__nand2_1
XFILLER_0_21_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15966_ ag2.body\[137\] net199 _01658_ ag2.body\[129\] vssd1 vssd1 vccd1 vccd1 _01195_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12340__A net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18754_ clknet_leaf_15_clk img_gen.tracker.next_frame\[192\] net1313 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[192\] sky130_fd_sc_hd__dfrtp_1
X_11089_ ag2.body\[536\] net1228 vssd1 vssd1 vccd1 vccd1 _06062_ sky130_fd_sc_hd__and2b_1
XFILLER_0_65_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17705_ net463 net372 _03383_ _03380_ vssd1 vssd1 vccd1 vccd1 _03384_ sky130_fd_sc_hd__a31o_1
X_14917_ control.body\[1076\] net170 _01542_ net2446 vssd1 vssd1 vccd1 vccd1 _00262_
+ sky130_fd_sc_hd__a22o_1
X_15897_ ag2.body\[204\] net133 _01650_ ag2.body\[196\] vssd1 vssd1 vccd1 vccd1 _01134_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__13690__B1 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18685_ clknet_leaf_28_clk img_gen.tracker.next_frame\[123\] net1337 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[123\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_91_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17636_ ag2.body\[162\] net862 vssd1 vssd1 vccd1 vccd1 _03315_ sky130_fd_sc_hd__nand2_1
XANTENNA__17420__A2 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14848_ _08768_ _08773_ _01514_ _01515_ _01518_ vssd1 vssd1 vccd1 vccd1 _01519_ sky130_fd_sc_hd__o2111a_2
XFILLER_0_114_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_1494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18639__RESET_B net1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17567_ _03240_ _03241_ _03242_ _03243_ vssd1 vssd1 vccd1 vccd1 _03246_ sky130_fd_sc_hd__a22o_1
XANTENNA__17708__B1 net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12339__X _07306_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14779_ net1001 ag2.body\[272\] vssd1 vssd1 vccd1 vccd1 _01450_ sky130_fd_sc_hd__xor2_1
XANTENNA__14267__A net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20610__1542 vssd1 vssd1 vccd1 vccd1 _20610__1542/HI net1542 sky130_fd_sc_hd__conb_1
X_16518_ net364 _02195_ _02196_ _02075_ vssd1 vssd1 vccd1 vccd1 _02197_ sky130_fd_sc_hd__o211a_1
X_19306_ clknet_leaf_99_clk _00250_ net1448 vssd1 vssd1 vccd1 vccd1 control.body\[1080\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_131_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17498_ ag2.body\[238\] net943 vssd1 vssd1 vccd1 vccd1 _03177_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_136_4461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_4472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_136_4483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_1556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16449_ obsg2.obstacleArray\[80\] obsg2.obstacleArray\[81\] net458 vssd1 vssd1 vccd1
+ vccd1 _02128_ sky130_fd_sc_hd__mux2_1
XANTENNA__17578__A ag2.body\[341\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19237_ clknet_leaf_84_clk _00181_ net1480 vssd1 vssd1 vccd1 vccd1 ag2.body\[100\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__18734__CLK clknet_leaf_142_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15195__B1 _01573_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11403__B net1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_132_4336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_132_4347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_132_4358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13745__A1 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19168_ clknet_leaf_52_clk _00112_ net1363 vssd1 vssd1 vccd1 vccd1 ag2.body\[31\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_41_1564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_41_1575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10019__B net1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18119_ net352 net38 _03633_ obsg2.obstacleArray\[60\] vssd1 vssd1 vccd1 vccd1 _03695_
+ sky130_fd_sc_hd__a31o_1
XANTENNA__17487__A2 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16144__C1 net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19099_ clknet_leaf_0_clk img_gen.tracker.next_frame\[537\] net1239 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[537\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_1421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12515__A net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09096__A ag2.body\[342\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16695__B1 net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20505__Q coll.badColl vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_1454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14170__A1 net997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17239__A2 net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout404 net405 vssd1 vssd1 vccd1 vccd1 net404 sky130_fd_sc_hd__clkbuf_4
XANTENNA__14170__B2 net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout415 net417 vssd1 vssd1 vccd1 vccd1 net415 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_54_1958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20012_ clknet_leaf_56_clk _00956_ net1457 vssd1 vssd1 vccd1 vccd1 ag2.body\[378\]
+ sky130_fd_sc_hd__dfrtp_4
Xfanout426 net429 vssd1 vssd1 vccd1 vccd1 net426 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_54_1969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_1486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09824__A net1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09823_ net1058 control.body\[927\] vssd1 vssd1 vccd1 vccd1 _04796_ sky130_fd_sc_hd__or2_1
Xfanout437 _06646_ vssd1 vssd1 vccd1 vccd1 net437 sky130_fd_sc_hd__clkbuf_4
Xfanout448 _02214_ vssd1 vssd1 vccd1 vccd1 net448 sky130_fd_sc_hd__buf_2
Xfanout459 _02060_ vssd1 vssd1 vccd1 vccd1 net459 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_35_1379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_1538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout387_A net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09754_ ag2.body\[215\] net1064 vssd1 vssd1 vccd1 vccd1 _04727_ sky130_fd_sc_hd__or2_1
XANTENNA__10689__B net1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09685_ ag2.body\[12\] net1128 vssd1 vssd1 vccd1 vccd1 _04658_ sky130_fd_sc_hd__xor2_1
XFILLER_0_55_1213 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17947__B1 obsg2.obstacleArray\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout554_A net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1296_A net1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_93_clk clknet_4_11__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_93_clk
+ sky130_fd_sc_hd__clkbuf_8
XPHY_EDGE_ROW_126_Right_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10495__B1 net1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11692__C1 net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout721_A _04265_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout342_X net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14177__A net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout819_A _03968_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1463_A net1464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1084_X net1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20367__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout44 net46 vssd1 vssd1 vccd1 vccd1 net44 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_88_1022 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout55 net62 vssd1 vssd1 vccd1 vccd1 net55 sky130_fd_sc_hd__clkbuf_4
Xfanout66 net67 vssd1 vssd1 vccd1 vccd1 net66 sky130_fd_sc_hd__clkbuf_4
Xfanout77 net79 vssd1 vssd1 vccd1 vccd1 net77 sky130_fd_sc_hd__buf_2
XANTENNA__11313__B net1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout88 net89 vssd1 vssd1 vccd1 vccd1 net88 sky130_fd_sc_hd__buf_2
Xfanout99 net100 vssd1 vssd1 vccd1 vccd1 net99 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout607_X net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_115_3822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17919__C net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_3298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_115_3833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10460_ ag2.body\[452\] net1127 vssd1 vssd1 vccd1 vccd1 _05433_ sky130_fd_sc_hd__xor2_1
XFILLER_0_91_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_115_3844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_21_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_1207 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_3708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09119_ ag2.body\[403\] vssd1 vssd1 vccd1 vccd1 _04144_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_111_3719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10391_ net638 _04632_ net892 vssd1 vssd1 vccd1 vccd1 _05364_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_115_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12130_ img_gen.tracker.frame\[564\] net622 net605 img_gen.tracker.frame\[567\] _07100_
+ vssd1 vssd1 vccd1 vccd1 _07102_ sky130_fd_sc_hd__o221a_1
XANTENNA__16150__A2 net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout976_X net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12061_ img_gen.tracker.frame\[60\] net627 net609 img_gen.tracker.frame\[63\] vssd1
+ vssd1 vccd1 vccd1 _07033_ sky130_fd_sc_hd__a22o_1
XANTENNA__14161__B2 net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16331__S net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold480 img_gen.tracker.frame\[294\] vssd1 vssd1 vccd1 vccd1 net2042 sky130_fd_sc_hd__dlygate4sd3_1
Xhold491 img_gen.tracker.frame\[394\] vssd1 vssd1 vccd1 vccd1 net2053 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_70_2450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11012_ _05975_ _05977_ _05979_ _05984_ vssd1 vssd1 vccd1 vccd1 _05985_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_70_2461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_3637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_2472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_3648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_3659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout960 net961 vssd1 vssd1 vccd1 vccd1 net960 sky130_fd_sc_hd__buf_4
X_15820_ ag2.body\[279\] net206 _01642_ ag2.body\[271\] vssd1 vssd1 vccd1 vccd1 _01065_
+ sky130_fd_sc_hd__a22o_1
Xfanout971 net974 vssd1 vssd1 vccd1 vccd1 net971 sky130_fd_sc_hd__buf_4
Xfanout982 ag2.randCord\[2\] vssd1 vssd1 vccd1 vccd1 net982 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_5_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout993 net994 vssd1 vssd1 vccd1 vccd1 net993 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_5_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15751_ ag2.body\[329\] net215 _01635_ ag2.body\[321\] vssd1 vssd1 vccd1 vccd1 _01003_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__17670__B net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12963_ net341 _07494_ vssd1 vssd1 vccd1 vccd1 _07678_ sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_84_clk clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_84_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_87_2980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_376 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_87_2991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14702_ net1020 ag2.body\[238\] vssd1 vssd1 vccd1 vccd1 _08863_ sky130_fd_sc_hd__xor2_1
X_18470_ net969 _03955_ vssd1 vssd1 vccd1 vccd1 _03956_ sky130_fd_sc_hd__nand2_1
X_11914_ img_gen.tracker.frame\[349\] net626 net569 vssd1 vssd1 vccd1 vccd1 _06886_
+ sky130_fd_sc_hd__o21a_1
XANTENNA__10486__B1 net1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15682_ ag2.body\[396\] net143 _01627_ ag2.body\[388\] vssd1 vssd1 vccd1 vccd1 _00942_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_87_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_83_2844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_2390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12894_ net267 _07645_ _07646_ net1985 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[205\]
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_83_2855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17421_ _04026_ net887 net720 ag2.body\[115\] _03099_ vssd1 vssd1 vccd1 vccd1 _03100_
+ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_83_2866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14633_ net1006 ag2.body\[583\] vssd1 vssd1 vccd1 vccd1 _08794_ sky130_fd_sc_hd__xor2_1
X_11845_ img_gen.tracker.frame\[506\] net617 net599 img_gen.tracker.frame\[509\] vssd1
+ vssd1 vccd1 vccd1 _06817_ sky130_fd_sc_hd__o22a_1
XANTENNA__18757__CLK clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_2265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14087__A net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_2276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_2287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17352_ _03019_ _03022_ vssd1 vssd1 vccd1 vccd1 _03031_ sky130_fd_sc_hd__nand2_1
XANTENNA__11504__A net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14564_ net1004 ag2.body\[352\] vssd1 vssd1 vccd1 vccd1 _08725_ sky130_fd_sc_hd__xor2_1
X_11776_ img_gen.tracker.frame\[155\] net580 net548 img_gen.tracker.frame\[152\] _06747_
+ vssd1 vssd1 vccd1 vccd1 _06748_ sky130_fd_sc_hd__o221a_1
XANTENNA__18363__B1 net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16303_ _01980_ _01981_ net415 vssd1 vssd1 vccd1 vccd1 _01982_ sky130_fd_sc_hd__mux2_1
X_13515_ net2128 net656 _07917_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[555\]
+ sky130_fd_sc_hd__and3_1
X_17283_ ag2.body\[310\] net944 vssd1 vssd1 vccd1 vccd1 _02962_ sky130_fd_sc_hd__xor2_1
XFILLER_0_86_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10727_ ag2.body\[252\] net1136 vssd1 vssd1 vccd1 vccd1 _05700_ sky130_fd_sc_hd__or2_1
XANTENNA__16506__S net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14495_ net1001 ag2.body\[256\] vssd1 vssd1 vccd1 vccd1 _08656_ sky130_fd_sc_hd__xor2_1
XANTENNA__14815__A net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19022_ clknet_leaf_1_clk img_gen.tracker.next_frame\[460\] net1246 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[460\] sky130_fd_sc_hd__dfrtp_1
X_16234_ obsg2.obstacleArray\[32\] obsg2.obstacleArray\[33\] net404 vssd1 vssd1 vccd1
+ vccd1 _01913_ sky130_fd_sc_hd__mux2_1
X_13446_ net682 _07890_ vssd1 vssd1 vccd1 vccd1 _07891_ sky130_fd_sc_hd__nor2_1
XANTENNA__14924__B1 _01543_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10658_ _05626_ _05627_ _05629_ _05630_ vssd1 vssd1 vccd1 vccd1 _05631_ sky130_fd_sc_hd__or4_1
Xclkload14 clknet_leaf_145_clk vssd1 vssd1 vccd1 vccd1 clkload14/Y sky130_fd_sc_hd__inv_8
XANTENNA__11738__B1 net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_2659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload25 clknet_leaf_15_clk vssd1 vssd1 vccd1 vccd1 clkload25/Y sky130_fd_sc_hd__bufinv_16
XFILLER_0_106_570 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16165_ net378 _01843_ _01842_ net347 vssd1 vssd1 vccd1 vccd1 _01844_ sky130_fd_sc_hd__a211o_1
XANTENNA__17469__A2 net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload36 clknet_leaf_17_clk vssd1 vssd1 vccd1 vccd1 clkload36/Y sky130_fd_sc_hd__inv_8
XFILLER_0_134_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkload47 clknet_leaf_29_clk vssd1 vssd1 vccd1 vccd1 clkload47/X sky130_fd_sc_hd__clkbuf_8
XANTENNA__09628__B net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13377_ _07539_ net304 vssd1 vssd1 vccd1 vccd1 _07864_ sky130_fd_sc_hd__nor2_1
Xclkload58 clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 clkload58/Y sky130_fd_sc_hd__inv_8
X_10589_ net1130 control.body\[828\] vssd1 vssd1 vccd1 vccd1 _05562_ sky130_fd_sc_hd__xor2_1
Xclkload69 clknet_leaf_45_clk vssd1 vssd1 vccd1 vccd1 clkload69/Y sky130_fd_sc_hd__inv_6
XFILLER_0_45_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15116_ net2660 net146 _01554_ control.body\[893\] vssd1 vssd1 vccd1 vccd1 _00439_
+ sky130_fd_sc_hd__a22o_1
X_12328_ _07251_ _07254_ _07288_ vssd1 vssd1 vccd1 vccd1 _07295_ sky130_fd_sc_hd__and3_1
X_16096_ net375 _01772_ _01774_ net348 vssd1 vssd1 vccd1 vccd1 _01775_ sky130_fd_sc_hd__a211o_1
XFILLER_0_50_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12054__B net1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14152__A1 net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19924_ clknet_leaf_52_clk _00868_ net1368 vssd1 vssd1 vccd1 vccd1 ag2.body\[466\]
+ sky130_fd_sc_hd__dfrtp_4
X_15047_ control.body\[967\] net163 _01556_ net2220 vssd1 vssd1 vccd1 vccd1 _00377_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__14152__B2 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12259_ _04391_ _07228_ vssd1 vssd1 vccd1 vccd1 _07229_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_10_Left_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19855_ clknet_leaf_91_clk _00799_ net1415 vssd1 vssd1 vccd1 vccd1 ag2.body\[541\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_125_4140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10713__A1 _04600_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11910__B1 net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18806_ clknet_leaf_3_clk img_gen.tracker.next_frame\[244\] net1248 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[244\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__17641__A2 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_4004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_121_4015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19786_ clknet_leaf_127_clk _00730_ net1328 vssd1 vssd1 vccd1 vccd1 ag2.body\[600\]
+ sky130_fd_sc_hd__dfrtp_4
X_16998_ ag2.body\[140\] net966 vssd1 vssd1 vccd1 vccd1 _02677_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_121_4026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19532__CLK clknet_leaf_118_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17580__B net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18737_ clknet_leaf_142_clk img_gen.tracker.next_frame\[175\] net1261 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[175\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_30_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15949_ ag2.body\[154\] net195 _01656_ ag2.body\[146\] vssd1 vssd1 vccd1 vccd1 _01180_
+ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_75_clk clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_75_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_95_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14860__C1 _08542_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15381__A _05856_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09470_ _04435_ _04436_ _04438_ _04442_ vssd1 vssd1 vccd1 vccd1 _04443_ sky130_fd_sc_hd__or4_1
X_18668_ clknet_leaf_10_clk img_gen.tracker.next_frame\[106\] net1273 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[106\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_52_1408 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09882__A2 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_4523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_4534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17619_ _04219_ net858 net688 ag2.body\[607\] _03296_ vssd1 vssd1 vccd1 vccd1 _03298_
+ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_138_4545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18599_ clknet_leaf_17_clk img_gen.tracker.next_frame\[37\] net1318 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[37\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_47_1762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_4567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11414__A net1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20630_ net1547 vssd1 vssd1 vccd1 vccd1 gpio_out[25] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_134_4409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13332__C _07813_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkload74_A clknet_leaf_115_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11977__B1 net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16924__B net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_1648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20561_ clknet_leaf_108_clk toggle1.nextDisplayOut\[1\] net1420 vssd1 vssd1 vccd1
+ vccd1 ssdec1.in\[1\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_15_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14725__A net1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout135_A net144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload8 clknet_leaf_1_clk vssd1 vssd1 vccd1 vccd1 clkload8/Y sky130_fd_sc_hd__inv_6
XTAP_TAPCELL_ROW_24_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20492_ clknet_leaf_24_clk _01379_ net1370 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[128\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__18106__B1 net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11729__B1 net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_3151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_3162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_3173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_1515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16668__B1 net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16151__S net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15340__B1 _01590_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14460__A net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1211_A net1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17880__A2 obsg2.obstacleCount\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout201 net204 vssd1 vssd1 vccd1 vccd1 net201 sky130_fd_sc_hd__buf_2
XFILLER_0_22_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout212 net213 vssd1 vssd1 vccd1 vccd1 net212 sky130_fd_sc_hd__buf_2
XANTENNA_fanout1309_A net1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout223 _07980_ vssd1 vssd1 vccd1 vccd1 net223 sky130_fd_sc_hd__buf_4
XFILLER_0_10_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__20166__RESET_B net1484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout234 net236 vssd1 vssd1 vccd1 vccd1 net234 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout671_A net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout292_X net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout245 net246 vssd1 vssd1 vccd1 vccd1 net245 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11901__B1 net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout769_A net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout256 net257 vssd1 vssd1 vccd1 vccd1 net256 sky130_fd_sc_hd__clkbuf_4
X_09806_ _04775_ _04776_ _04777_ _04778_ vssd1 vssd1 vccd1 vccd1 _04779_ sky130_fd_sc_hd__a22o_1
XFILLER_0_22_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout267 net268 vssd1 vssd1 vccd1 vccd1 net267 sky130_fd_sc_hd__clkbuf_4
XANTENNA__13076__A net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17632__A2 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout278 net279 vssd1 vssd1 vccd1 vccd1 net278 sky130_fd_sc_hd__clkbuf_4
Xfanout289 net295 vssd1 vssd1 vccd1 vccd1 net289 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_104_3501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09737_ _04705_ _04706_ _04707_ _04709_ vssd1 vssd1 vccd1 vccd1 _04710_ sky130_fd_sc_hd__a211o_1
XANTENNA__11308__B net1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout936_A obsg2.randCord\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16387__A net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_66_clk clknet_4_13__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_66_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout557_X net557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09668_ net639 _04640_ vssd1 vssd1 vccd1 vccd1 _04641_ sky130_fd_sc_hd__and2b_1
XFILLER_0_97_858 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09873__A2 _04830_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout724_X net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_379 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09599_ net643 _04571_ vssd1 vssd1 vccd1 vccd1 _04572_ sky130_fd_sc_hd__and2_1
XFILLER_0_132_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11630_ obsg2.obstacleArray\[38\] net631 vssd1 vssd1 vccd1 vccd1 _06603_ sky130_fd_sc_hd__or2_1
XFILLER_0_65_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15803__A_N _04984_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_3906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_13_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09625__A2 _04597_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16834__B net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11968__B1 net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11561_ obsg2.obstacleArray\[71\] net632 net513 obsg2.obstacleArray\[67\] net507
+ vssd1 vssd1 vccd1 vccd1 _06534_ sky130_fd_sc_hd__o221a_1
XFILLER_0_108_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13300_ net235 _07833_ _07834_ net1594 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[423\]
+ sky130_fd_sc_hd__a22o_1
X_10512_ ag2.body\[103\] net1064 vssd1 vssd1 vccd1 vccd1 _05485_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_24_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14280_ net821 ag2.body\[139\] ag2.body\[142\] net803 vssd1 vssd1 vccd1 vccd1 _08441_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_11_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xwire635 _04633_ vssd1 vssd1 vccd1 vccd1 net635 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_110_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11492_ _06461_ _06463_ vssd1 vssd1 vccd1 vccd1 _06465_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_134_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16371__A2 _01947_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19405__CLK clknet_leaf_103_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13231_ net673 _07426_ vssd1 vssd1 vccd1 vccd1 _07805_ sky130_fd_sc_hd__nor2_1
XFILLER_0_134_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17946__A net48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10443_ net1204 control.body\[929\] vssd1 vssd1 vccd1 vccd1 _05416_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_33_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11196__A1 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11196__B2 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_2512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13162_ net277 _07770_ _07771_ net1862 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[347\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_103_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_72_2523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10374_ net923 _05346_ _04432_ net641 vssd1 vssd1 vccd1 vccd1 _05347_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_72_2534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18113__Y _03691_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12113_ img_gen.tracker.frame\[162\] net554 net563 vssd1 vssd1 vccd1 vccd1 _07085_
+ sky130_fd_sc_hd__a21o_1
X_17970_ obsg2.obstacleArray\[12\] _03593_ net529 vssd1 vssd1 vccd1 vccd1 _01263_
+ sky130_fd_sc_hd__o21a_1
X_13093_ net291 _07737_ _07738_ net1952 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[311\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__19555__CLK clknet_leaf_115_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12145__B1 net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12044_ img_gen.tracker.frame\[240\] net627 net609 img_gen.tracker.frame\[243\] vssd1
+ vssd1 vccd1 vccd1 _07016_ sky130_fd_sc_hd__a22o_1
X_16921_ _02597_ _02598_ _02599_ vssd1 vssd1 vccd1 vccd1 _02600_ sky130_fd_sc_hd__and3_1
XANTENNA__12696__A1 net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17084__B1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19640_ clknet_leaf_123_clk _00584_ net1405 vssd1 vssd1 vccd1 vccd1 control.body\[758\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_121_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16852_ ag2.body\[171\] net717 net691 ag2.body\[175\] vssd1 vssd1 vccd1 vccd1 _02531_
+ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_85_2906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout790 net791 vssd1 vssd1 vccd1 vccd1 net790 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_85_2917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15803_ _04984_ net49 vssd1 vssd1 vccd1 vccd1 _01641_ sky130_fd_sc_hd__and2b_2
X_16783_ net462 _02459_ _02461_ _01699_ vssd1 vssd1 vccd1 vccd1 _02462_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_85_2928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19571_ clknet_leaf_116_clk _00515_ net1385 vssd1 vssd1 vccd1 vccd1 control.body\[817\]
+ sky130_fd_sc_hd__dfrtp_1
X_13995_ ag2.body\[131\] net213 _08160_ ag2.body\[123\] vssd1 vssd1 vccd1 vccd1 _00212_
+ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_57_clk clknet_4_12__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_57_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__14842__C1 _01510_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_2327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_66_2338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18522_ clknet_leaf_42_clk net1578 net1372 vssd1 vssd1 vccd1 vccd1 control.detect4.Q\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_15734_ ag2.body\[346\] net212 _01633_ ag2.body\[338\] vssd1 vssd1 vccd1 vccd1 _00988_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__09911__B net1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12946_ _07483_ net339 net335 vssd1 vssd1 vccd1 vccd1 _07670_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_66_2349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15665_ ag2.body\[413\] net142 _01625_ ag2.body\[405\] vssd1 vssd1 vccd1 vccd1 _00927_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_115_1442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18453_ _04635_ _03839_ _03940_ _03941_ vssd1 vssd1 vccd1 vccd1 _03942_ sky130_fd_sc_hd__o31a_1
X_12877_ _07425_ _07638_ net678 vssd1 vssd1 vccd1 vccd1 _07640_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_5_1526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14616_ net1034 ag2.body\[60\] vssd1 vssd1 vccd1 vccd1 _08777_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_8_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17404_ ag2.body\[46\] net937 vssd1 vssd1 vccd1 vccd1 _03083_ sky130_fd_sc_hd__xor2_1
XFILLER_0_111_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18384_ _03799_ _03870_ _03871_ _03872_ net321 vssd1 vssd1 vccd1 vccd1 _03874_ sky130_fd_sc_hd__a32o_1
X_11828_ _06781_ _06787_ _06793_ _06799_ net473 net437 vssd1 vssd1 vccd1 vccd1 _06800_
+ sky130_fd_sc_hd__mux4_1
X_15596_ ag2.body\[479\] net122 _01618_ ag2.body\[471\] vssd1 vssd1 vccd1 vccd1 _00865_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__14070__B1 ag2.body\[213\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17335_ _03013_ vssd1 vssd1 vccd1 vccd1 _03014_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14547_ net975 ag2.body\[243\] vssd1 vssd1 vccd1 vccd1 _08708_ sky130_fd_sc_hd__or2_1
XANTENNA__16236__S net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_1504 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11759_ img_gen.tracker.frame\[278\] net618 net601 img_gen.tracker.frame\[281\] vssd1
+ vssd1 vccd1 vccd1 _06731_ sky130_fd_sc_hd__o22a_1
XFILLER_0_55_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14545__A net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_131 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17266_ _04080_ net873 net721 ag2.body\[251\] vssd1 vssd1 vccd1 vccd1 _02945_ sky130_fd_sc_hd__o22a_1
X_14478_ net1027 ag2.body\[445\] vssd1 vssd1 vccd1 vccd1 _08639_ sky130_fd_sc_hd__xor2_1
XANTENNA__16362__A2 net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload103 clknet_leaf_101_clk vssd1 vssd1 vccd1 vccd1 clkload103/Y sky130_fd_sc_hd__bufinv_16
Xclkload114 clknet_leaf_61_clk vssd1 vssd1 vccd1 vccd1 clkload114/Y sky130_fd_sc_hd__inv_8
X_16217_ net355 _01893_ vssd1 vssd1 vccd1 vccd1 _01896_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_102_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19005_ clknet_leaf_2_clk img_gen.tracker.next_frame\[443\] net1245 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[443\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkload125 clknet_leaf_83_clk vssd1 vssd1 vccd1 vccd1 clkload125/Y sky130_fd_sc_hd__inv_8
X_13429_ net225 _07882_ _07883_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[503\]
+ sky130_fd_sc_hd__o21ai_1
X_17197_ ag2.body\[178\] net861 vssd1 vssd1 vccd1 vccd1 _02876_ sky130_fd_sc_hd__nand2_1
XFILLER_0_10_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14832__X _01503_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_460 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__20055__Q ag2.body\[341\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_1392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16148_ net379 _01826_ _01825_ net349 vssd1 vssd1 vccd1 vccd1 _01827_ sky130_fd_sc_hd__a211o_1
XANTENNA__17575__B net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20062__CLK clknet_leaf_73_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_1402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_127_4202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16079_ _01756_ _01757_ net376 vssd1 vssd1 vccd1 vccd1 _01758_ sky130_fd_sc_hd__mux2_1
X_08970_ ag2.body\[57\] vssd1 vssd1 vccd1 vccd1 _03995_ sky130_fd_sc_hd__inv_2
XFILLER_0_45_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_36_1430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12136__B1 net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19907_ clknet_leaf_54_clk _00851_ net1457 vssd1 vssd1 vccd1 vccd1 ag2.body\[481\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_62_1592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12512__B net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19838_ clknet_leaf_122_clk _00782_ net1414 vssd1 vssd1 vccd1 vccd1 ag2.body\[556\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__17614__A2 net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput1 en vssd1 vssd1 vccd1 vccd1 net1 sky130_fd_sc_hd__buf_1
XANTENNA__12439__A1 net1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11128__B net1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_803 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19769_ clknet_leaf_16_clk _00713_ net1322 vssd1 vssd1 vccd1 vccd1 control.body\[631\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10032__B net1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09522_ net1130 control.body\[836\] vssd1 vssd1 vccd1 vccd1 _04495_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_49_1813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_1824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16000__A net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11111__A1 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09453_ net910 net917 net913 net922 vssd1 vssd1 vccd1 vccd1 _04426_ sky130_fd_sc_hd__and4_1
XANTENNA_fanout252_A net254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_571 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09384_ _04357_ _04376_ vssd1 vssd1 vccd1 vccd1 _01411_ sky130_fd_sc_hd__nor2_1
XFILLER_0_47_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20613_ net1556 vssd1 vssd1 vccd1 vccd1 gpio_oeb[25] sky130_fd_sc_hd__buf_2
XFILLER_0_74_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_95_3213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12611__A1 net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_703 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14455__A net1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1161_A net1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10983__A net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout138_X net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_3224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout517_A net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16373__C net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_3235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16889__B1 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20544_ clknet_leaf_105_clk _01409_ _00018_ vssd1 vssd1 vccd1 vccd1 sound_gen.osc1.stayCount\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_62_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16353__A2 net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1025 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20475_ clknet_leaf_32_clk _01362_ net1352 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[111\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_104_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout305_X net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19578__CLK clknet_leaf_118_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1047_X net1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_780 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1492 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20347__RESET_B net1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout886_A net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1214_X net1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_3028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_7_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1007 net1014 vssd1 vssd1 vccd1 vccd1 net1007 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_89_3039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10090_ net773 control.body\[794\] control.body\[796\] net758 vssd1 vssd1 vccd1 vccd1
+ _05063_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_7_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1018 net1019 vssd1 vssd1 vccd1 vccd1 net1018 sky130_fd_sc_hd__buf_4
XANTENNA__12678__A1 net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1029 ag2.randCord\[5\] vssd1 vssd1 vccd1 vccd1 net1029 sky130_fd_sc_hd__buf_4
XANTENNA_fanout674_X net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17605__A2 net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16388__Y _02067_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout841_X net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout939_X net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_39_clk clknet_4_5__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_39_clk
+ sky130_fd_sc_hd__clkbuf_8
X_12800_ net278 _07601_ _07602_ net1996 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[155\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_134_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13780_ img_gen.updater.commands.count\[11\] _08088_ vssd1 vssd1 vccd1 vccd1 _08090_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_138_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10992_ ag2.body\[338\] net1186 vssd1 vssd1 vccd1 vccd1 _05965_ sky130_fd_sc_hd__xor2_1
XFILLER_0_96_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10877__B net1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12731_ net284 _07568_ _07569_ net1838 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[119\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__16577__C1 net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12850__A1 net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15450_ ag2.body\[606\] net86 _01601_ ag2.body\[598\] vssd1 vssd1 vccd1 vccd1 _00736_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_32_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12662_ net386 _07444_ _07535_ vssd1 vssd1 vccd1 vccd1 _07536_ sky130_fd_sc_hd__and3_1
X_14401_ _08555_ _08557_ _08561_ vssd1 vssd1 vccd1 vccd1 _08562_ sky130_fd_sc_hd__or3_1
XFILLER_0_37_232 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11613_ obsg2.obstacleArray\[58\] obsg2.obstacleArray\[59\] obsg2.obstacleArray\[62\]
+ obsg2.obstacleArray\[63\] net1126 net511 vssd1 vssd1 vccd1 vccd1 _06586_ sky130_fd_sc_hd__mux4_1
XANTENNA__16329__C1 net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15381_ _05856_ net52 vssd1 vssd1 vccd1 vccd1 _01595_ sky130_fd_sc_hd__nor2_2
X_12593_ net471 net569 net542 _07312_ vssd1 vssd1 vccd1 vccd1 _07497_ sky130_fd_sc_hd__or4_1
XANTENNA__10893__A net1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14365__A net996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17120_ _02795_ _02796_ _02797_ _02798_ vssd1 vssd1 vccd1 vccd1 _02799_ sky130_fd_sc_hd__or4_1
XANTENNA__11341__X _06314_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14332_ net835 ag2.body\[425\] ag2.body\[430\] net800 vssd1 vssd1 vccd1 vccd1 _08493_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_78_2710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11544_ obsg2.obstacleArray\[111\] net631 net511 obsg2.obstacleArray\[107\] net1125
+ vssd1 vssd1 vccd1 vccd1 _06517_ sky130_fd_sc_hd__o221a_1
XFILLER_0_80_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_747 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_59_2120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_59_2131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14355__A1 net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17051_ _04085_ net885 net719 ag2.body\[259\] _02729_ vssd1 vssd1 vccd1 vccd1 _02730_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_29_1218 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14355__B2 net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14263_ net989 ag2.body\[9\] vssd1 vssd1 vccd1 vccd1 _08424_ sky130_fd_sc_hd__nand2_1
XANTENNA__11501__B net1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11475_ ag2.body\[491\] net1162 vssd1 vssd1 vccd1 vccd1 _06448_ sky130_fd_sc_hd__or2_1
Xwire476 _06064_ vssd1 vssd1 vccd1 vccd1 net476 sky130_fd_sc_hd__buf_1
XFILLER_0_81_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16002_ net883 net948 vssd1 vssd1 vccd1 vccd1 _01681_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_55_2006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13214_ net675 _07796_ vssd1 vssd1 vccd1 vccd1 _07797_ sky130_fd_sc_hd__nor2_1
X_10426_ net638 _05073_ _04632_ vssd1 vssd1 vccd1 vccd1 _05399_ sky130_fd_sc_hd__a21o_1
X_14194_ net834 ag2.body\[161\] ag2.body\[162\] net826 _08354_ vssd1 vssd1 vccd1 vccd1
+ _08355_ sky130_fd_sc_hd__a221o_1
XFILLER_0_0_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_1110 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13145_ _07493_ net327 net336 vssd1 vssd1 vccd1 vccd1 _07764_ sky130_fd_sc_hd__and3b_1
XANTENNA__09906__B net1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10357_ ag2.body\[292\] net1142 vssd1 vssd1 vccd1 vccd1 _05330_ sky130_fd_sc_hd__and2b_1
XFILLER_0_42_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12613__A net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17953_ _03549_ _03564_ _03579_ net298 vssd1 vssd1 vccd1 vccd1 _03580_ sky130_fd_sc_hd__and4b_1
X_13076_ net343 _07561_ vssd1 vssd1 vccd1 vccd1 _07731_ sky130_fd_sc_hd__nor2_1
X_10288_ ag2.body\[330\] net1186 vssd1 vssd1 vccd1 vccd1 _05261_ sky130_fd_sc_hd__nand2_1
XANTENNA__11229__A net1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09534__B2 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12027_ net577 _06995_ _06998_ vssd1 vssd1 vccd1 vccd1 _06999_ sky130_fd_sc_hd__o21a_1
X_16904_ ag2.body\[240\] net885 vssd1 vssd1 vccd1 vccd1 _02583_ sky130_fd_sc_hd__xor2_1
XANTENNA__10133__A net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17884_ _04422_ _04445_ _03523_ vssd1 vssd1 vccd1 vccd1 _03524_ sky130_fd_sc_hd__o21a_1
XANTENNA__11341__A1 net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19623_ clknet_leaf_123_clk _00567_ net1406 vssd1 vssd1 vccd1 vccd1 control.body\[773\]
+ sky130_fd_sc_hd__dfrtp_1
X_16835_ ag2.body\[101\] net951 vssd1 vssd1 vccd1 vccd1 _02514_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_75_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16280__A1 net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19554_ clknet_leaf_116_clk _00498_ net1397 vssd1 vssd1 vccd1 vccd1 control.body\[832\]
+ sky130_fd_sc_hd__dfrtp_1
X_13978_ ag2.body\[116\] net202 _08158_ ag2.body\[108\] vssd1 vssd1 vccd1 vccd1 _00197_
+ sky130_fd_sc_hd__a22o_1
X_16766_ obsg2.obstacleArray\[7\] net502 net484 obsg2.obstacleArray\[5\] _02444_ vssd1
+ vssd1 vccd1 vccd1 _02445_ sky130_fd_sc_hd__a221o_1
XFILLER_0_73_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1612 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18505_ net1515 net1509 vssd1 vssd1 vccd1 vccd1 _00036_ sky130_fd_sc_hd__or2_1
X_15717_ ag2.body\[364\] net194 _01630_ ag2.body\[356\] vssd1 vssd1 vccd1 vccd1 _00974_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__13163__B _07505_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12929_ net343 _07472_ vssd1 vssd1 vccd1 vccd1 _07662_ sky130_fd_sc_hd__nor2_1
X_16697_ obsg2.obstacleArray\[70\] net488 net484 obsg2.obstacleArray\[69\] vssd1 vssd1
+ vccd1 vccd1 _02376_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_17_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19485_ clknet_leaf_114_clk _00429_ net1399 vssd1 vssd1 vccd1 vccd1 control.body\[907\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_17_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18436_ track.nextHighScore\[3\] _03794_ _03814_ vssd1 vssd1 vccd1 vccd1 _03925_
+ sky130_fd_sc_hd__a21bo_1
X_15648_ ag2.body\[430\] net138 _01623_ ag2.body\[422\] vssd1 vssd1 vccd1 vccd1 _00912_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_115_1272 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16474__B net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20428__CLK clknet_4_6__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11899__A net1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14594__B2 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15579_ _04429_ _04718_ net64 vssd1 vssd1 vccd1 vccd1 _01617_ sky130_fd_sc_hd__and3_2
X_18367_ _08030_ _03834_ _03823_ vssd1 vssd1 vccd1 vccd1 _03861_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_84_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17318_ ag2.body\[220\] net964 vssd1 vssd1 vccd1 vccd1 _02997_ sky130_fd_sc_hd__xor2_1
XFILLER_0_7_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11801__C1 net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16335__A2 net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18298_ _08053_ _03783_ _03792_ vssd1 vssd1 vccd1 vccd1 _03794_ sky130_fd_sc_hd__a21oi_4
XANTENNA__19720__CLK clknet_leaf_132_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14346__A1 net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17586__A ag2.body\[60\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14346__B2 net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17249_ _02922_ _02927_ vssd1 vssd1 vccd1 vccd1 _02928_ sky130_fd_sc_hd__or2_2
XANTENNA__10308__A net1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20260_ clknet_leaf_43_clk _01204_ net1379 vssd1 vssd1 vccd1 vccd1 ag2.body\[2\]
+ sky130_fd_sc_hd__dfstp_4
XFILLER_0_98_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_wire475_X net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10027__B net1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20191_ clknet_leaf_88_clk _01135_ net1459 vssd1 vssd1 vccd1 vccd1 ag2.body\[205\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__12372__A3 net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11580__A1 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08953_ ag2.body\[12\] vssd1 vssd1 vccd1 vccd1 _03978_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_102_Left_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13857__B1 _08134_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10314__Y _05287_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17048__B1 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13321__A2 net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10043__A net1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19100__CLK clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1007_A net1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18260__A2 net37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10978__A net1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout467_A net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12896__C net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10330__X _05303_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10697__B net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09505_ ag2.body\[404\] net1139 vssd1 vssd1 vccd1 vccd1 _04478_ sky130_fd_sc_hd__xor2_1
XFILLER_0_78_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19250__CLK clknet_leaf_75_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12832__A1 net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_817 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout255_X net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout634_A _04697_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1376_A net1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17220__B1 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_144_clk_X clknet_leaf_144_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09436_ ag2.body\[3\] net1153 vssd1 vssd1 vccd1 vccd1 _04409_ sky130_fd_sc_hd__xor2_1
XFILLER_0_94_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10843__B1 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_407 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18818__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_111_Left_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout801_A net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09367_ sound_gen.osc1.stayCount\[20\] _04368_ vssd1 vssd1 vccd1 vccd1 _04369_ sky130_fd_sc_hd__nand2_1
XFILLER_0_136_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1164_X net1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09298_ sound_gen.osc1.count\[7\] _04308_ _04317_ vssd1 vssd1 vccd1 vccd1 _04318_
+ sky130_fd_sc_hd__a21oi_1
XANTENNA__12060__A2 net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09461__B1 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12417__B net1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20527_ clknet_leaf_114_clk _01392_ net1398 vssd1 vssd1 vccd1 vccd1 toggle1.bcd_tens\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_65_1418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09566__X _04539_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11260_ net773 control.body\[770\] _04241_ net1050 _06229_ vssd1 vssd1 vccd1 vccd1
+ _06233_ sky130_fd_sc_hd__a221o_1
X_20458_ clknet_leaf_38_clk _01345_ net1354 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[94\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout791_X net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout889_X net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17287__B1 net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10211_ net1157 control.body\[995\] vssd1 vssd1 vccd1 vccd1 _05184_ sky130_fd_sc_hd__or2_1
XANTENNA__13529__A _07624_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11191_ net1151 control.body\[875\] vssd1 vssd1 vccd1 vccd1 _06164_ sky130_fd_sc_hd__or2_1
X_20389_ clknet_leaf_42_clk _01276_ net1371 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[25\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_31_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10142_ net1099 control.body\[821\] vssd1 vssd1 vccd1 vccd1 _05115_ sky130_fd_sc_hd__nand2_1
XFILLER_0_101_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13248__B net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13816__X _08113_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17039__B1 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10073_ net1119 control.body\[716\] vssd1 vssd1 vccd1 vccd1 _05046_ sky130_fd_sc_hd__xor2_1
X_14950_ net2580 net172 _01546_ net2284 vssd1 vssd1 vccd1 vccd1 _00291_ sky130_fd_sc_hd__a22o_1
XANTENNA__12720__X _07564_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13901_ _05588_ net52 vssd1 vssd1 vccd1 vccd1 _08150_ sky130_fd_sc_hd__nor2_2
X_14881_ control.body\[1108\] net179 _01538_ control.body\[1100\] vssd1 vssd1 vccd1
+ vccd1 _00230_ sky130_fd_sc_hd__a22o_1
XANTENNA__10888__A net1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13264__A net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13832_ net1755 net662 _08126_ _08121_ vssd1 vssd1 vccd1 vccd1 _00081_ sky130_fd_sc_hd__a31o_1
X_16620_ obsg2.obstacleArray\[44\] obsg2.obstacleArray\[45\] net441 vssd1 vssd1 vccd1
+ vccd1 _02299_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_1200 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16551_ obsg2.obstacleArray\[102\] net441 net390 _02229_ vssd1 vssd1 vccd1 vccd1
+ _02230_ sky130_fd_sc_hd__o211a_1
X_13763_ _08077_ _08078_ img_gen.updater.commands.count\[5\] net320 vssd1 vssd1 vccd1
+ vccd1 _00062_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__11626__A2 net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_997 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10975_ _05941_ _05942_ _05943_ _05946_ vssd1 vssd1 vccd1 vccd1 _05948_ sky130_fd_sc_hd__and4_1
XFILLER_0_35_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16014__A1 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_1632 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15502_ ag2.body\[556\] net113 _01607_ ag2.body\[548\] vssd1 vssd1 vccd1 vccd1 _00782_
+ sky130_fd_sc_hd__a22o_1
X_12714_ net335 _07448_ vssd1 vssd1 vccd1 vccd1 _07561_ sky130_fd_sc_hd__or2_2
X_19270_ clknet_leaf_68_clk _00214_ net1498 vssd1 vssd1 vccd1 vccd1 ag2.body\[133\]
+ sky130_fd_sc_hd__dfrtp_2
X_16482_ obsg2.obstacleArray\[46\] obsg2.obstacleArray\[47\] net452 vssd1 vssd1 vccd1
+ vccd1 _02161_ sky130_fd_sc_hd__mux2_1
X_13694_ _08032_ _08034_ vssd1 vssd1 vccd1 vccd1 _08036_ sky130_fd_sc_hd__or2_2
XFILLER_0_6_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18221_ obsg2.obstacleArray\[107\] _03749_ net524 vssd1 vssd1 vccd1 vccd1 _01358_
+ sky130_fd_sc_hd__o21a_1
X_15433_ ag2.body\[623\] net84 _01599_ ag2.body\[615\] vssd1 vssd1 vccd1 vccd1 _00721_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_66_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12645_ net295 _07524_ _07525_ net1929 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[77\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_52_1580 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14095__A net992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12608__A net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18152_ net298 _03579_ net37 obsg2.obstacleArray\[73\] vssd1 vssd1 vccd1 vccd1 _03715_
+ sky130_fd_sc_hd__a31o_1
X_15364_ net2659 net75 _01593_ net2211 vssd1 vssd1 vccd1 vccd1 _00658_ sky130_fd_sc_hd__a22o_1
XFILLER_0_65_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12051__A2 net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13430__C _07813_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12576_ net678 _07488_ vssd1 vssd1 vccd1 vccd1 _07489_ sky130_fd_sc_hd__nor2_1
XFILLER_0_108_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17103_ ag2.body\[10\] net724 net696 ag2.body\[14\] vssd1 vssd1 vccd1 vccd1 _02782_
+ sky130_fd_sc_hd__a22o_1
X_14315_ net1015 ag2.body\[54\] vssd1 vssd1 vccd1 vccd1 _08476_ sky130_fd_sc_hd__xor2_1
XFILLER_0_68_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11527_ obsg2.obstacleArray\[127\] net631 net511 obsg2.obstacleArray\[123\] net1125
+ vssd1 vssd1 vccd1 vccd1 _06500_ sky130_fd_sc_hd__o221a_1
XANTENNA__15919__A _04831_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18083_ obsg2.obstacleArray\[47\] _03671_ net523 vssd1 vssd1 vccd1 vccd1 _01298_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_81_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15295_ control.body\[739\] net76 _01585_ net2386 vssd1 vssd1 vccd1 vccd1 _00597_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_123_432 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16514__S net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10128__A net1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17034_ ag2.body\[125\] net954 vssd1 vssd1 vccd1 vccd1 _02713_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_34_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold309 img_gen.tracker.frame\[257\] vssd1 vssd1 vccd1 vccd1 net1871 sky130_fd_sc_hd__dlygate4sd3_1
X_14246_ net814 ag2.body\[540\] ag2.body\[542\] net804 vssd1 vssd1 vccd1 vccd1 _08407_
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_106_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11458_ ag2.body\[258\] net1187 vssd1 vssd1 vccd1 vccd1 _06431_ sky130_fd_sc_hd__nand2_1
XFILLER_0_7_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10409_ _05376_ _05377_ _05378_ _05381_ vssd1 vssd1 vccd1 vccd1 _05382_ sky130_fd_sc_hd__or4_1
XFILLER_0_46_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14177_ net982 ag2.body\[194\] vssd1 vssd1 vccd1 vccd1 _08338_ sky130_fd_sc_hd__nand2_1
XANTENNA__12343__A net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11389_ net1097 control.body\[645\] vssd1 vssd1 vccd1 vccd1 _06362_ sky130_fd_sc_hd__nand2_1
XANTENNA__11562__A1 net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19123__CLK clknet_leaf_141_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13128_ net684 _07755_ vssd1 vssd1 vccd1 vccd1 _07756_ sky130_fd_sc_hd__nor2_1
XFILLER_0_42_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18985_ clknet_leaf_9_clk img_gen.tracker.next_frame\[423\] net1271 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[423\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__14500__A1 net975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14500__B2 net1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17936_ net47 net296 _03566_ vssd1 vssd1 vccd1 vccd1 _03567_ sky130_fd_sc_hd__and3_1
X_13059_ net338 net330 _07433_ vssd1 vssd1 vccd1 vccd1 _07723_ sky130_fd_sc_hd__and3_2
XANTENNA__18030__A net45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1009 control.body\[1055\] vssd1 vssd1 vccd1 vccd1 net2571 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12997__B net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1360 net1361 vssd1 vssd1 vccd1 vccd1 net1360 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09652__A net1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1371 net1373 vssd1 vssd1 vccd1 vccd1 net1371 sky130_fd_sc_hd__clkbuf_4
Xfanout1382 net1383 vssd1 vssd1 vccd1 vccd1 net1382 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_94_1636 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19273__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17867_ img_gen.updater.commands.rR1.rainbowRNG\[8\] img_gen.updater.commands.rR1.rainbowRNG\[7\]
+ _03501_ net2166 vssd1 vssd1 vccd1 vccd1 _03514_ sky130_fd_sc_hd__a31oi_1
XFILLER_0_108_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1393 net1394 vssd1 vssd1 vccd1 vccd1 net1393 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_17_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13174__A net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19606_ clknet_leaf_120_clk _00550_ net1393 vssd1 vssd1 vccd1 vccd1 control.body\[788\]
+ sky130_fd_sc_hd__dfrtp_1
X_16818_ _04011_ net887 net706 ag2.body\[85\] _02494_ vssd1 vssd1 vccd1 vccd1 _02497_
+ sky130_fd_sc_hd__a221o_1
XANTENNA__13067__A1 net246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17798_ _04261_ net709 net703 vssd1 vssd1 vccd1 vccd1 _03470_ sky130_fd_sc_hd__or3_1
XFILLER_0_108_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14803__A2 ag2.body\[288\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19537_ clknet_leaf_118_clk _00481_ net1394 vssd1 vssd1 vccd1 vccd1 control.body\[863\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11406__B net1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16749_ obsg2.obstacleArray\[63\] net501 net487 obsg2.obstacleArray\[62\] vssd1 vssd1
+ vccd1 vccd1 _02428_ sky130_fd_sc_hd__a22o_1
XANTENNA__11617__A2 net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12814__A1 net239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1355 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10825__B1 net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19468_ clknet_leaf_109_clk _00412_ net1416 vssd1 vssd1 vccd1 vccd1 control.body\[922\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_1328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14717__B ag2.body\[341\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09221_ control.body\[886\] vssd1 vssd1 vccd1 vccd1 _04246_ sky130_fd_sc_hd__inv_2
XFILLER_0_91_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18419_ _04646_ _08032_ _03890_ _03907_ _03908_ vssd1 vssd1 vccd1 vccd1 _03909_ sky130_fd_sc_hd__a32o_1
XANTENNA__14567__B2 net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_714 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19399_ clknet_leaf_102_clk _00343_ net1429 vssd1 vssd1 vccd1 vccd1 control.body\[997\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_130_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_259 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11422__A net1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09152_ ag2.body\[487\] vssd1 vssd1 vccd1 vccd1 _04177_ sky130_fd_sc_hd__inv_2
XFILLER_0_133_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14319__A1 net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11141__B net1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14319__B2 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09083_ ag2.body\[319\] vssd1 vssd1 vccd1 vccd1 _04108_ sky130_fd_sc_hd__inv_2
XANTENNA__16424__S _02076_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10038__A net1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_1175 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20312_ clknet_leaf_44_clk _01212_ net1380 vssd1 vssd1 vccd1 vccd1 ag2.randCord\[6\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_115_988 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_1039 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold810 control.body\[783\] vssd1 vssd1 vccd1 vccd1 net2372 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_936 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold821 control.body\[944\] vssd1 vssd1 vccd1 vccd1 net2383 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold832 _00232_ vssd1 vssd1 vccd1 vccd1 net2394 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold843 control.body\[855\] vssd1 vssd1 vccd1 vccd1 net2405 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__17269__B1 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20243_ clknet_leaf_70_clk _01187_ net1497 vssd1 vssd1 vccd1 vccd1 ag2.body\[145\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_29_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold854 control.body\[633\] vssd1 vssd1 vccd1 vccd1 net2416 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10356__A2 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1124_A net1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold865 control.body\[950\] vssd1 vssd1 vccd1 vccd1 net2427 sky130_fd_sc_hd__dlygate4sd3_1
Xhold876 _00295_ vssd1 vssd1 vccd1 vccd1 net2438 sky130_fd_sc_hd__dlygate4sd3_1
Xhold887 control.body\[844\] vssd1 vssd1 vccd1 vccd1 net2449 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_51_clk_A clknet_4_6__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20174_ clknet_leaf_82_clk _01118_ net1480 vssd1 vssd1 vccd1 vccd1 ag2.body\[220\]
+ sky130_fd_sc_hd__dfrtp_2
Xhold898 _00373_ vssd1 vssd1 vccd1 vccd1 net2460 sky130_fd_sc_hd__dlygate4sd3_1
X_09985_ net1086 control.body\[1118\] vssd1 vssd1 vccd1 vccd1 _04958_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout584_A net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08936_ control.divider.fsm.current_mode\[0\] vssd1 vssd1 vccd1 vccd1 _03961_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout372_X net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout751_A net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14389__A1_N net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1493_A net1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_66_clk_A clknet_4_13__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout849_A net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10501__A net1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13058__A1 net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18640__CLK clknet_leaf_15_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11608__A2 net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12805__A1 net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10220__B net1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_3968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout637_X net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_120_3979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10760_ net1157 control.body\[891\] vssd1 vssd1 vccd1 vccd1 _05733_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_101_3389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14558__A1 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09419_ obsg2.obstacleCount\[3\] _04397_ vssd1 vssd1 vccd1 vccd1 _04398_ sky130_fd_sc_hd__nand2_1
XANTENNA__14558__B2 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10691_ _05658_ _05659_ _05663_ _05237_ vssd1 vssd1 vccd1 vccd1 _05664_ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout804_X net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12428__A net1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_124_clk_A clknet_4_9__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12430_ _06627_ _06629_ _07390_ _07352_ vssd1 vssd1 vccd1 vccd1 _07392_ sky130_fd_sc_hd__a31o_1
XFILLER_0_47_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_911 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13230__A1 net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16842__B net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_864 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12361_ img_gen.updater.commands.rR1.rainbowRNG\[8\] _07319_ _07320_ _07321_ _07327_
+ vssd1 vssd1 vccd1 vccd1 _07328_ sky130_fd_sc_hd__a221o_1
XFILLER_0_63_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14643__A net1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19146__CLK clknet_leaf_51_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14100_ net1034 ag2.body\[588\] vssd1 vssd1 vccd1 vccd1 _08261_ sky130_fd_sc_hd__xor2_1
X_11312_ ag2.body\[277\] net1112 vssd1 vssd1 vccd1 vccd1 _06285_ sky130_fd_sc_hd__xor2_1
X_15080_ net2650 net148 _01561_ net2404 vssd1 vssd1 vccd1 vccd1 _00406_ sky130_fd_sc_hd__a22o_1
X_12292_ img_gen.updater.commands.mode\[2\] img_gen.control.current\[0\] _04388_ _07183_
+ vssd1 vssd1 vccd1 vccd1 _07261_ sky130_fd_sc_hd__or4b_1
XFILLER_0_22_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_139_clk_A clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14031_ net977 ag2.body\[499\] vssd1 vssd1 vccd1 vccd1 _08192_ sky130_fd_sc_hd__xor2_1
XANTENNA__14730__A1 net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11243_ ag2.body\[197\] net1104 vssd1 vssd1 vccd1 vccd1 _06216_ sky130_fd_sc_hd__xor2_1
XANTENNA__13259__A net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_969 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14730__B2 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_19_clk_A clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11174_ net1226 control.body\[776\] vssd1 vssd1 vccd1 vccd1 _06147_ sky130_fd_sc_hd__xor2_1
XANTENNA__10898__A3 _05074_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19296__CLK clknet_leaf_98_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17680__B1 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10125_ _05094_ _05095_ _05096_ _05097_ _05093_ vssd1 vssd1 vccd1 vccd1 _05098_ sky130_fd_sc_hd__a221o_1
XFILLER_0_98_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18770_ clknet_leaf_16_clk img_gen.tracker.next_frame\[208\] net1321 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[208\] sky130_fd_sc_hd__dfrtp_1
X_15982_ _01661_ _01665_ _01666_ _01660_ net1602 vssd1 vssd1 vccd1 vccd1 _01203_ sky130_fd_sc_hd__a32o_1
XANTENNA__13297__A1 net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17721_ _03396_ _03399_ _01728_ vssd1 vssd1 vccd1 vccd1 _03400_ sky130_fd_sc_hd__mux2_1
XANTENNA__18558__Q ag2.x\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10912__B1_N _04447_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20273__CLK clknet_leaf_37_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10056_ ag2.body\[482\] net1177 vssd1 vssd1 vccd1 vccd1 _05029_ sky130_fd_sc_hd__xor2_1
X_14933_ control.body\[1058\] net168 _01544_ net2501 vssd1 vssd1 vccd1 vccd1 _00276_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11066__X _06039_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17432__B1 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11507__A net1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17652_ ag2.body\[35\] net715 net928 _03986_ _03326_ vssd1 vssd1 vccd1 vccd1 _03331_
+ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_19_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14864_ _01506_ _01520_ _01534_ vssd1 vssd1 vccd1 vccd1 _01535_ sky130_fd_sc_hd__and3_2
XANTENNA__10411__A net1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16603_ _02279_ _02280_ _02281_ net392 net360 vssd1 vssd1 vccd1 vccd1 _02282_ sky130_fd_sc_hd__a221o_1
XFILLER_0_86_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13815_ _04276_ control.detect3.Q\[1\] vssd1 vssd1 vccd1 vccd1 _08112_ sky130_fd_sc_hd__nor2_1
XFILLER_0_118_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14797__A1 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17583_ _03258_ _03259_ _03261_ _03257_ vssd1 vssd1 vccd1 vccd1 _03262_ sky130_fd_sc_hd__a211o_1
XANTENNA__14797__B2 net1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14795_ _01459_ _01460_ _01461_ _01465_ vssd1 vssd1 vccd1 vccd1 _01466_ sky130_fd_sc_hd__or4_1
XANTENNA__16509__S net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19322_ clknet_leaf_104_clk _00266_ net1433 vssd1 vssd1 vccd1 vccd1 control.body\[1064\]
+ sky130_fd_sc_hd__dfrtp_1
X_16534_ _01733_ _02204_ vssd1 vssd1 vccd1 vccd1 _02213_ sky130_fd_sc_hd__and2_1
XFILLER_0_85_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13746_ img_gen.updater.commands.count\[1\] img_gen.updater.commands.count\[0\] vssd1
+ vssd1 vccd1 vccd1 _08066_ sky130_fd_sc_hd__nand2_1
X_10958_ ag2.body\[174\] net1081 vssd1 vssd1 vccd1 vccd1 _05931_ sky130_fd_sc_hd__or2_1
XFILLER_0_15_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17735__A1 _03248_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_1451 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18009__B net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14549__A1 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19253_ clknet_leaf_74_clk _00197_ net1500 vssd1 vssd1 vccd1 vccd1 ag2.body\[116\]
+ sky130_fd_sc_hd__dfrtp_4
X_16465_ obsg2.obstacleArray\[56\] obsg2.obstacleArray\[57\] net454 vssd1 vssd1 vccd1
+ vccd1 _02144_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13677_ _04402_ net464 vssd1 vssd1 vccd1 vccd1 _08024_ sky130_fd_sc_hd__nand2_2
XANTENNA__14549__B2 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12338__A net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10889_ net1146 control.body\[651\] vssd1 vssd1 vccd1 vccd1 _05862_ sky130_fd_sc_hd__or2_1
X_18204_ _03647_ net40 vssd1 vssd1 vccd1 vccd1 _03741_ sky130_fd_sc_hd__nor2_1
X_12628_ net2133 net645 _07516_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[69\]
+ sky130_fd_sc_hd__and3_1
X_15416_ _05685_ net63 vssd1 vssd1 vccd1 vccd1 _01598_ sky130_fd_sc_hd__and2_2
X_16396_ net461 _02065_ vssd1 vssd1 vccd1 vccd1 _02075_ sky130_fd_sc_hd__xnor2_4
X_19184_ clknet_leaf_20_clk _00128_ net1365 vssd1 vssd1 vccd1 vccd1 ag2.body\[47\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_13_1372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13221__A1 net241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18135_ _03549_ net41 vssd1 vssd1 vccd1 vccd1 _03706_ sky130_fd_sc_hd__or2_2
X_15347_ control.body\[689\] net75 _01591_ control.body\[681\] vssd1 vssd1 vccd1 vccd1
+ _00643_ sky130_fd_sc_hd__a22o_1
XFILLER_0_41_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12559_ net226 _07477_ _07478_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[38\]
+ sky130_fd_sc_hd__o21bai_1
XANTENNA__14553__A net1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18025__A net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10586__A2 net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09647__A net1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_130_4275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18066_ net300 _03582_ vssd1 vssd1 vccd1 vccd1 _03660_ sky130_fd_sc_hd__nand2_1
XANTENNA__11896__B net1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15278_ net2562 net88 _01583_ control.body\[748\] vssd1 vssd1 vccd1 vccd1 _00582_
+ sky130_fd_sc_hd__a22o_1
Xhold106 img_gen.tracker.frame\[392\] vssd1 vssd1 vccd1 vccd1 net1668 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_130_4286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold117 img_gen.tracker.frame\[175\] vssd1 vssd1 vccd1 vccd1 net1679 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_130_4297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_9_Right_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_622 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold128 img_gen.tracker.frame\[489\] vssd1 vssd1 vccd1 vccd1 net1690 sky130_fd_sc_hd__dlygate4sd3_1
X_17017_ ag2.body\[333\] net954 vssd1 vssd1 vccd1 vccd1 _02696_ sky130_fd_sc_hd__xor2_1
XANTENNA__13169__A net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold139 img_gen.tracker.frame\[408\] vssd1 vssd1 vccd1 vccd1 net1701 sky130_fd_sc_hd__dlygate4sd3_1
X_14229_ net997 net988 net1035 net1007 vssd1 vssd1 vccd1 vccd1 _08390_ sky130_fd_sc_hd__or4_1
XFILLER_0_111_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11535__A1 _06505_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout608 _06476_ vssd1 vssd1 vccd1 vccd1 net608 sky130_fd_sc_hd__clkbuf_4
XANTENNA__18463__A2 net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout619 net620 vssd1 vssd1 vccd1 vccd1 net619 sky130_fd_sc_hd__buf_2
XFILLER_0_61_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_107_Right_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09770_ ag2.body\[233\] net1206 vssd1 vssd1 vccd1 vccd1 _04743_ sky130_fd_sc_hd__or2_1
XANTENNA__12801__A net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18968_ clknet_leaf_6_clk img_gen.tracker.next_frame\[406\] net1269 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[406\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__18663__CLK clknet_leaf_13_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17919_ net957 net539 net462 net537 vssd1 vssd1 vccd1 vccd1 _03553_ sky130_fd_sc_hd__or4b_1
XANTENNA__11838__A2 _06807_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18899_ clknet_leaf_144_clk img_gen.tracker.next_frame\[337\] net1251 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[337\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_52_1897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_1542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1190 net1191 vssd1 vssd1 vccd1 vccd1 net1190 sky130_fd_sc_hd__clkbuf_4
XANTENNA__16777__A2 net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_603 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout165_A net171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout332_A net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1074_A net1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19169__CLK clknet_leaf_52_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09204_ net1174 vssd1 vssd1 vccd1 vccd1 _04229_ sky130_fd_sc_hd__inv_2
XFILLER_0_134_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1248 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13212__A1 net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09135_ ag2.body\[448\] vssd1 vssd1 vccd1 vccd1 _04160_ sky130_fd_sc_hd__inv_2
XANTENNA__15559__A _04686_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10991__A ag2.body\[337\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14463__A net1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout218_X net218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09557__A net1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09066_ ag2.body\[267\] vssd1 vssd1 vccd1 vccd1 _04091_ sky130_fd_sc_hd__inv_2
XANTENNA__16701__A2 net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_113_3761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_3772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_113_3783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout799_A net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17774__A _03440_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold640 img_gen.tracker.frame\[334\] vssd1 vssd1 vccd1 vccd1 net2202 sky130_fd_sc_hd__dlygate4sd3_1
Xhold651 control.body\[766\] vssd1 vssd1 vccd1 vccd1 net2213 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1127_X net1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold662 _00311_ vssd1 vssd1 vccd1 vccd1 net2224 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09844__X _04817_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20226_ clknet_leaf_66_clk _01170_ net1476 vssd1 vssd1 vccd1 vccd1 ag2.body\[160\]
+ sky130_fd_sc_hd__dfrtp_4
Xhold673 control.body\[786\] vssd1 vssd1 vccd1 vccd1 net2235 sky130_fd_sc_hd__dlygate4sd3_1
Xhold684 toggle1.bcd_ones\[1\] vssd1 vssd1 vccd1 vccd1 net2246 sky130_fd_sc_hd__dlygate4sd3_1
Xhold695 control.body\[758\] vssd1 vssd1 vccd1 vccd1 net2257 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout966_A net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17924__D net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout587_X net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09968_ ag2.body\[80\] net1235 vssd1 vssd1 vccd1 vccd1 _04941_ sky130_fd_sc_hd__xor2_1
X_20157_ clknet_leaf_94_clk _01101_ net1441 vssd1 vssd1 vccd1 vccd1 ag2.body\[235\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_42_1590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09899_ _04004_ net1211 net1117 _04008_ _04871_ vssd1 vssd1 vccd1 vccd1 _04872_ sky130_fd_sc_hd__a221o_1
X_20088_ clknet_leaf_78_clk _01032_ net1490 vssd1 vssd1 vccd1 vccd1 ag2.body\[310\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA_fanout754_X net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17414__B1 net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_3576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11930_ net439 _06901_ vssd1 vssd1 vccd1 vccd1 _06902_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_107_3587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_3598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16396__Y _02075_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11046__B net1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11861_ img_gen.tracker.frame\[214\] net591 net552 img_gen.tracker.frame\[211\] _06832_
+ vssd1 vssd1 vccd1 vccd1 _06833_ sky130_fd_sc_hd__o221a_1
XFILLER_0_68_912 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13600_ _03960_ control.divider.count\[16\] control.divider.count\[17\] _07951_ vssd1
+ vssd1 vccd1 vccd1 _07975_ sky130_fd_sc_hd__o211a_1
XFILLER_0_79_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13542__A net226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10812_ net1159 control.body\[1091\] vssd1 vssd1 vccd1 vccd1 _05785_ sky130_fd_sc_hd__nand2_1
X_14580_ net826 ag2.body\[490\] ag2.body\[488\] net842 vssd1 vssd1 vccd1 vccd1 _08741_
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_138_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11792_ img_gen.tracker.frame\[380\] net549 _06763_ net575 vssd1 vssd1 vccd1 vccd1
+ _06764_ sky130_fd_sc_hd__o211a_1
XFILLER_0_32_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13531_ net2116 net656 _07923_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[565\]
+ sky130_fd_sc_hd__and3_1
XANTENNA__17949__A net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10743_ ag2.body\[501\] net1114 vssd1 vssd1 vccd1 vccd1 _05716_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_81_2783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11462__B1 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_1562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_95_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_2794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16250_ _01893_ _01928_ vssd1 vssd1 vccd1 vccd1 _01929_ sky130_fd_sc_hd__nand2_1
X_13462_ net235 _07896_ _07897_ net1640 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[522\]
+ sky130_fd_sc_hd__a22o_1
X_10674_ ag2.body\[351\] net1065 vssd1 vssd1 vccd1 vccd1 _05647_ sky130_fd_sc_hd__xor2_1
XANTENNA__17668__B net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18116__Y _03693_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15201_ net2497 net95 _01574_ control.body\[808\] vssd1 vssd1 vccd1 vccd1 _00514_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_49_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16940__A2 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12413_ img_gen.updater.commands.rR1.rainbowRNG\[12\] _07319_ _07338_ _07368_ _07375_
+ vssd1 vssd1 vccd1 vccd1 _07376_ sky130_fd_sc_hd__a221o_1
X_16181_ obsg2.obstacleArray\[38\] obsg2.obstacleArray\[39\] net423 vssd1 vssd1 vccd1
+ vccd1 _01860_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_11_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09958__B2 _04903_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13393_ net671 _07870_ vssd1 vssd1 vccd1 vccd1 _07871_ sky130_fd_sc_hd__nor2_1
XANTENNA__14373__A net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_1046 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_11_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10568__A2 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15132_ control.body\[883\] net107 _01566_ net2515 vssd1 vssd1 vccd1 vccd1 _00453_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_106_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12344_ net435 _07305_ vssd1 vssd1 vccd1 vccd1 _07311_ sky130_fd_sc_hd__nor2_1
XANTENNA__18591__RESET_B net1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19940_ clknet_leaf_47_clk _00884_ net1376 vssd1 vssd1 vccd1 vccd1 ag2.body\[450\]
+ sky130_fd_sc_hd__dfrtp_4
X_15063_ control.body\[949\] net150 _01559_ net2300 vssd1 vssd1 vccd1 vccd1 _00391_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_49_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12275_ _07243_ _07244_ vssd1 vssd1 vccd1 vccd1 _07245_ sky130_fd_sc_hd__and2b_1
XFILLER_0_82_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10406__A net1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_2598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_1490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14014_ net1027 ag2.body\[461\] vssd1 vssd1 vccd1 vccd1 _08175_ sky130_fd_sc_hd__xor2_1
X_11226_ net778 control.body\[857\] control.body\[863\] net744 vssd1 vssd1 vccd1 vccd1
+ _06199_ sky130_fd_sc_hd__o22a_1
XFILLER_0_120_1500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19871_ clknet_leaf_95_clk _00815_ net1440 vssd1 vssd1 vccd1 vccd1 ag2.body\[525\]
+ sky130_fd_sc_hd__dfrtp_4
X_18822_ clknet_leaf_2_clk img_gen.tracker.next_frame\[260\] net1248 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[260\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__09914__B net1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11157_ ag2.body\[606\] net1073 vssd1 vssd1 vccd1 vccd1 _06130_ sky130_fd_sc_hd__xor2_1
XANTENNA__12621__A net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10108_ net1157 control.body\[939\] vssd1 vssd1 vccd1 vccd1 _05081_ sky130_fd_sc_hd__or2_1
X_18753_ clknet_leaf_144_clk img_gen.tracker.next_frame\[191\] net1255 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[191\] sky130_fd_sc_hd__dfrtp_1
X_15965_ ag2.body\[136\] net212 _01658_ ag2.body\[128\] vssd1 vssd1 vccd1 vccd1 _01194_
+ sky130_fd_sc_hd__a22o_1
X_11088_ ag2.body\[538\] net1180 vssd1 vssd1 vccd1 vccd1 _06061_ sky130_fd_sc_hd__and2b_1
XANTENNA__12340__B _07306_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17704_ _03381_ _03382_ net416 vssd1 vssd1 vccd1 vccd1 _03383_ sky130_fd_sc_hd__mux2_1
XANTENNA__17405__B1 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10039_ net1227 control.body\[896\] vssd1 vssd1 vccd1 vccd1 _05012_ sky130_fd_sc_hd__xor2_1
X_14916_ control.body\[1075\] net170 _01542_ net2183 vssd1 vssd1 vccd1 vccd1 _00261_
+ sky130_fd_sc_hd__a22o_1
X_18684_ clknet_leaf_28_clk img_gen.tracker.next_frame\[122\] net1336 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[122\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__10141__A net1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16759__A2 net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15896_ ag2.body\[203\] net133 _01650_ ag2.body\[195\] vssd1 vssd1 vccd1 vccd1 _01133_
+ sky130_fd_sc_hd__a22o_1
X_17635_ ag2.body\[162\] net862 vssd1 vssd1 vccd1 vccd1 _03314_ sky130_fd_sc_hd__or2_1
X_14847_ _08280_ _08447_ _08914_ _01517_ vssd1 vssd1 vccd1 vccd1 _01518_ sky130_fd_sc_hd__and4_1
XFILLER_0_77_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14548__A net1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_400 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11524__X _06497_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13442__A1 net235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17566_ _04209_ net869 net858 _04210_ _03244_ vssd1 vssd1 vccd1 vccd1 _03245_ sky130_fd_sc_hd__a221o_1
X_14778_ net837 ag2.body\[273\] ag2.body\[275\] net820 vssd1 vssd1 vccd1 vccd1 _01449_
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_114_1359 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10795__B net1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19305_ clknet_leaf_99_clk _00249_ net1448 vssd1 vssd1 vccd1 vccd1 control.body\[1095\]
+ sky130_fd_sc_hd__dfrtp_1
X_16517_ net402 _02188_ _02187_ net366 vssd1 vssd1 vccd1 vccd1 _02196_ sky130_fd_sc_hd__a211o_1
XANTENNA__13171__B net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13729_ _07221_ _07254_ _04391_ vssd1 vssd1 vccd1 vccd1 _00052_ sky130_fd_sc_hd__mux2_1
XANTENNA__12068__A net1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17497_ ag2.body\[238\] net943 vssd1 vssd1 vccd1 vccd1 _03176_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_136_4462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_4473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19236_ clknet_leaf_84_clk _00180_ net1481 vssd1 vssd1 vccd1 vccd1 ag2.body\[99\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_136_4484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16448_ net402 _02126_ _02125_ net367 vssd1 vssd1 vccd1 vccd1 _02127_ sky130_fd_sc_hd__a211o_1
XANTENNA__17578__B net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_4337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_132_4348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_4359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19167_ clknet_leaf_52_clk _00111_ net1363 vssd1 vssd1 vccd1 vccd1 ag2.body\[30\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_41_1565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16379_ net956 _01888_ _02052_ vssd1 vssd1 vccd1 vccd1 _02058_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_41_1576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10559__A2 net1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_1587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18118_ obsg2.obstacleArray\[59\] _03694_ net525 vssd1 vssd1 vccd1 vccd1 _01310_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_30_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_571 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19098_ clknet_leaf_145_clk img_gen.tracker.next_frame\[536\] net1243 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[536\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_1433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15498__A2 net113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1287 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18049_ net301 _03562_ vssd1 vssd1 vccd1 vccd1 _03649_ sky130_fd_sc_hd__nand2_1
XFILLER_0_26_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_91_3090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout405 net406 vssd1 vssd1 vccd1 vccd1 net405 sky130_fd_sc_hd__buf_2
Xfanout416 net417 vssd1 vssd1 vccd1 vccd1 net416 sky130_fd_sc_hd__clkbuf_4
XANTENNA__18202__B net40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout427 net429 vssd1 vssd1 vccd1 vccd1 net427 sky130_fd_sc_hd__buf_2
X_20011_ clknet_leaf_59_clk _00955_ net1467 vssd1 vssd1 vccd1 vccd1 ag2.body\[377\]
+ sky130_fd_sc_hd__dfrtp_4
X_09822_ _04788_ _04790_ _04792_ _04794_ vssd1 vssd1 vccd1 vccd1 _04795_ sky130_fd_sc_hd__nand4_1
XTAP_TAPCELL_ROW_54_1959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout438 net439 vssd1 vssd1 vccd1 vccd1 net438 sky130_fd_sc_hd__buf_2
Xfanout449 net451 vssd1 vssd1 vccd1 vccd1 net449 sky130_fd_sc_hd__clkbuf_4
X_09753_ ag2.body\[215\] net1064 vssd1 vssd1 vccd1 vccd1 _04726_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout282_A _07335_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15670__A2 net195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09684_ ag2.body\[11\] net1152 vssd1 vssd1 vccd1 vccd1 _04657_ sky130_fd_sc_hd__xor2_1
XFILLER_0_55_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17947__A1 net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09840__A net1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10986__A net1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_102_3440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1191_A net1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout547_A net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16080__C1 _01742_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13433__A1 net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18559__CLK clknet_leaf_132_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13984__A2 net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout45 net46 vssd1 vssd1 vccd1 vccd1 net45 sky130_fd_sc_hd__clkbuf_4
Xfanout56 net62 vssd1 vssd1 vccd1 vccd1 net56 sky130_fd_sc_hd__buf_6
XANTENNA_fanout1077_X net1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout67 _08131_ vssd1 vssd1 vccd1 vccd1 net67 sky130_fd_sc_hd__buf_4
XFILLER_0_33_1589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_1183 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17488__B net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout78 net79 vssd1 vssd1 vccd1 vccd1 net78 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout89 net90 vssd1 vssd1 vccd1 vccd1 net89 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_98_3299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_115_3823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_3834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout502_X net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14193__A net1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_115_3845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18124__A1 net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12706__A net225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09118_ ag2.body\[402\] vssd1 vssd1 vccd1 vccd1 _04143_ sky130_fd_sc_hd__inv_2
XFILLER_0_60_631 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_111_3709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10390_ net1060 control.body\[1063\] vssd1 vssd1 vccd1 vccd1 _05363_ sky130_fd_sc_hd__or2_1
XFILLER_0_66_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16686__A1 net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15489__A2 net113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09049_ ag2.body\[239\] vssd1 vssd1 vccd1 vccd1 _04074_ sky130_fd_sc_hd__inv_2
XFILLER_0_130_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_4_4__f_clk clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_4__leaf_clk sky130_fd_sc_hd__clkbuf_16
XANTENNA__14921__A net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12060_ img_gen.tracker.frame\[57\] net593 net554 img_gen.tracker.frame\[54\] _07031_
+ vssd1 vssd1 vccd1 vccd1 _07032_ sky130_fd_sc_hd__a221o_1
Xhold470 img_gen.tracker.frame\[22\] vssd1 vssd1 vccd1 vccd1 net2032 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout871_X net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold481 control.divider.count\[13\] vssd1 vssd1 vccd1 vccd1 net2043 sky130_fd_sc_hd__dlygate4sd3_1
Xhold492 img_gen.tracker.frame\[455\] vssd1 vssd1 vccd1 vccd1 net2054 sky130_fd_sc_hd__dlygate4sd3_1
X_11011_ _05983_ _05981_ _05980_ _05982_ vssd1 vssd1 vccd1 vccd1 _05984_ sky130_fd_sc_hd__and4b_1
X_20209_ clknet_leaf_54_clk _01153_ net1456 vssd1 vssd1 vccd1 vccd1 ag2.body\[191\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_40_1538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_70_2451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_2462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_3638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_2473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_3649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_1163 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16989__A2 net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout950 obsg2.randCord\[5\] vssd1 vssd1 vccd1 vccd1 net950 sky130_fd_sc_hd__buf_4
Xfanout961 net968 vssd1 vssd1 vccd1 vccd1 net961 sky130_fd_sc_hd__buf_4
XANTENNA__11263__A1_N net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout972 net974 vssd1 vssd1 vccd1 vccd1 net972 sky130_fd_sc_hd__buf_4
Xfanout983 net984 vssd1 vssd1 vccd1 vccd1 net983 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_5_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout994 net995 vssd1 vssd1 vccd1 vccd1 net994 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_5_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_5_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15750_ ag2.body\[328\] net215 _01635_ ag2.body\[320\] vssd1 vssd1 vccd1 vccd1 _01002_
+ sky130_fd_sc_hd__a22o_1
X_12962_ net278 _07676_ _07677_ net1948 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[242\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__19334__CLK clknet_leaf_103_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_2970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14701_ _08854_ _08856_ _08861_ vssd1 vssd1 vccd1 vccd1 _08862_ sky130_fd_sc_hd__or3_4
XTAP_TAPCELL_ROW_87_2981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11913_ img_gen.tracker.frame\[352\] net598 net580 img_gen.tracker.frame\[358\] vssd1
+ vssd1 vccd1 vccd1 _06885_ sky130_fd_sc_hd__o22a_1
XANTENNA__11683__B1 net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15681_ ag2.body\[395\] net142 _01627_ ag2.body\[387\] vssd1 vssd1 vccd1 vccd1 _00941_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_115_1602 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12893_ net246 _07645_ _07646_ net1928 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[204\]
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_83_2845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_2391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_2856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17420_ ag2.body\[118\] net701 net695 ag2.body\[119\] vssd1 vssd1 vccd1 vccd1 _03099_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_83_2867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11844_ img_gen.tracker.frame\[518\] net620 net544 img_gen.tracker.frame\[524\] _06815_
+ vssd1 vssd1 vccd1 vccd1 _06816_ sky130_fd_sc_hd__o221a_1
X_14632_ net798 ag2.body\[582\] ag2.body\[580\] net811 vssd1 vssd1 vccd1 vccd1 _08793_
+ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__13424__A1 net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_2266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_2277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_64_2288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14563_ net1032 ag2.body\[357\] vssd1 vssd1 vccd1 vccd1 _08724_ sky130_fd_sc_hd__xor2_1
X_17351_ net925 net924 ag2.body\[7\] _03013_ _03015_ vssd1 vssd1 vccd1 vccd1 _03030_
+ sky130_fd_sc_hd__o32a_1
XANTENNA__11504__B net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11775_ img_gen.tracker.frame\[146\] net621 net603 img_gen.tracker.frame\[149\] vssd1
+ vssd1 vccd1 vccd1 _06747_ sky130_fd_sc_hd__o22a_1
XFILLER_0_51_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_797 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11986__A1 _06945_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16302_ obsg2.obstacleArray\[98\] obsg2.obstacleArray\[99\] net404 vssd1 vssd1 vccd1
+ vccd1 _01981_ sky130_fd_sc_hd__mux2_1
X_13514_ _07615_ _07807_ vssd1 vssd1 vccd1 vccd1 _07917_ sky130_fd_sc_hd__or2_1
X_10726_ ag2.body\[252\] net1136 vssd1 vssd1 vccd1 vccd1 _05699_ sky130_fd_sc_hd__nand2_1
X_14494_ net1022 ag2.body\[262\] vssd1 vssd1 vccd1 vccd1 _08655_ sky130_fd_sc_hd__xor2_1
X_17282_ _02955_ _02956_ _02960_ _02954_ vssd1 vssd1 vccd1 vccd1 _02961_ sky130_fd_sc_hd__a211o_1
XFILLER_0_137_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16913__A2 net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19021_ clknet_leaf_1_clk img_gen.tracker.next_frame\[459\] net1246 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[459\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16233_ net460 _01905_ vssd1 vssd1 vccd1 vccd1 _01912_ sky130_fd_sc_hd__xnor2_4
X_13445_ _07578_ net302 vssd1 vssd1 vccd1 vccd1 _07890_ sky130_fd_sc_hd__nor2_1
XFILLER_0_36_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10657_ ag2.body\[283\] net1164 vssd1 vssd1 vccd1 vccd1 _05630_ sky130_fd_sc_hd__xor2_1
XFILLER_0_3_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkload15 clknet_leaf_146_clk vssd1 vssd1 vccd1 vccd1 clkload15/Y sky130_fd_sc_hd__inv_12
XFILLER_0_51_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkload26 clknet_leaf_131_clk vssd1 vssd1 vccd1 vccd1 clkload26/Y sky130_fd_sc_hd__inv_6
X_16164_ obsg2.obstacleArray\[10\] obsg2.obstacleArray\[11\] net426 vssd1 vssd1 vccd1
+ vccd1 _01843_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13376_ net280 _07862_ _07863_ net1930 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[470\]
+ sky130_fd_sc_hd__a22o_1
Xclkload37 clknet_leaf_18_clk vssd1 vssd1 vccd1 vccd1 clkload37/Y sky130_fd_sc_hd__clkinv_4
X_10588_ net1051 control.body\[831\] vssd1 vssd1 vccd1 vccd1 _05561_ sky130_fd_sc_hd__or2_1
XFILLER_0_106_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkload48 clknet_leaf_30_clk vssd1 vssd1 vccd1 vccd1 clkload48/Y sky130_fd_sc_hd__inv_12
XANTENNA__09628__C _04239_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16677__A1 net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload59 clknet_leaf_23_clk vssd1 vssd1 vccd1 vccd1 clkload59/Y sky130_fd_sc_hd__inv_6
XFILLER_0_23_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15115_ control.body\[900\] net146 _01554_ net2318 vssd1 vssd1 vccd1 vccd1 _00438_
+ sky130_fd_sc_hd__a22o_1
X_12327_ _07289_ _07291_ _07293_ vssd1 vssd1 vccd1 vccd1 _07294_ sky130_fd_sc_hd__nand3_1
X_16095_ obsg2.obstacleArray\[119\] net430 net377 _01773_ vssd1 vssd1 vccd1 vccd1
+ _01774_ sky130_fd_sc_hd__o211a_1
XFILLER_0_11_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19923_ clknet_leaf_51_clk _00867_ net1368 vssd1 vssd1 vccd1 vccd1 ag2.body\[465\]
+ sky130_fd_sc_hd__dfrtp_4
X_15046_ net2579 net164 _01556_ control.body\[958\] vssd1 vssd1 vccd1 vccd1 _00376_
+ sky130_fd_sc_hd__a22o_1
X_12258_ img_gen.updater.commands.cmd_num\[4\] _07188_ _07227_ vssd1 vssd1 vccd1 vccd1
+ _07228_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_107_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11209_ _04446_ _05051_ net636 vssd1 vssd1 vccd1 vccd1 _06182_ sky130_fd_sc_hd__o21a_1
X_19854_ clknet_leaf_93_clk _00798_ net1413 vssd1 vssd1 vccd1 vccd1 ag2.body\[540\]
+ sky130_fd_sc_hd__dfrtp_4
X_12189_ net1222 ag2.apple_cord\[0\] vssd1 vssd1 vccd1 vccd1 _07161_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_125_4130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_125_4141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18805_ clknet_leaf_3_clk img_gen.tracker.next_frame\[243\] net1258 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[243\] sky130_fd_sc_hd__dfrtp_1
X_19785_ clknet_leaf_126_clk _00729_ net1332 vssd1 vssd1 vccd1 vccd1 ag2.body\[615\]
+ sky130_fd_sc_hd__dfrtp_4
X_16997_ ag2.body\[139\] net856 vssd1 vssd1 vccd1 vccd1 _02676_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_121_4005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15652__A2 net139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_121_4027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1482 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_1550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18736_ clknet_leaf_142_clk img_gen.tracker.next_frame\[174\] net1257 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[174\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_30_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15948_ ag2.body\[153\] net195 _01656_ ag2.body\[145\] vssd1 vssd1 vccd1 vccd1 _01179_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_30_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20465__RESET_B net1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14860__B1 _01530_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15381__B net52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18667_ clknet_leaf_11_clk img_gen.tracker.next_frame\[105\] net1282 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[105\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__14278__A net1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15879_ ag2.body\[220\] net192 _01648_ ag2.body\[212\] vssd1 vssd1 vccd1 vccd1 _01118_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_25_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19827__CLK clknet_leaf_124_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_4524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17618_ ag2.body\[603\] net715 net698 ag2.body\[606\] _03290_ vssd1 vssd1 vccd1 vccd1
+ _03297_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_138_4535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18598_ clknet_leaf_13_clk img_gen.tracker.next_frame\[36\] net1318 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[36\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_138_4546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17549_ _04109_ net887 net934 _04112_ _03227_ vssd1 vssd1 vccd1 vccd1 _03228_ sky130_fd_sc_hd__a221o_1
XANTENNA__16493__A net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17157__A2 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_28_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_15_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20560_ clknet_leaf_109_clk toggle1.nextDisplayOut\[0\] net1421 vssd1 vssd1 vccd1
+ vccd1 ssdec1.in\[0\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_43_1649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_24_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload9 clknet_leaf_2_clk vssd1 vssd1 vccd1 vccd1 clkload9/Y sky130_fd_sc_hd__bufinv_16
XFILLER_0_55_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19219_ clknet_leaf_67_clk _00163_ net1495 vssd1 vssd1 vccd1 vccd1 ag2.body\[82\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__17101__B net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20491_ clknet_leaf_38_clk _01378_ net1354 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[127\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__09819__B _04791_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12526__A net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout128_A net219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_3152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_3163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_3174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_1062 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10046__A net1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17755__C _03426_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1037_A net1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09835__A net1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout497_A net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout202 net203 vssd1 vssd1 vccd1 vccd1 net202 sky130_fd_sc_hd__buf_2
XANTENNA__17617__B1 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout213 net214 vssd1 vssd1 vccd1 vccd1 net213 sky130_fd_sc_hd__clkbuf_2
XANTENNA__13357__A net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout224 _03489_ vssd1 vssd1 vccd1 vccd1 net224 sky130_fd_sc_hd__buf_2
XANTENNA_fanout1204_A net1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout235 net236 vssd1 vssd1 vccd1 vccd1 net235 sky130_fd_sc_hd__clkbuf_4
Xfanout246 net247 vssd1 vssd1 vccd1 vccd1 net246 sky130_fd_sc_hd__clkbuf_4
XANTENNA_input2_A gpio_in[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09805_ net1181 control.body\[962\] vssd1 vssd1 vccd1 vccd1 _04778_ sky130_fd_sc_hd__or2_1
Xfanout257 net260 vssd1 vssd1 vccd1 vccd1 net257 sky130_fd_sc_hd__clkbuf_4
XANTENNA__13076__B _07561_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09570__A2 net1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout268 net269 vssd1 vssd1 vccd1 vccd1 net268 sky130_fd_sc_hd__clkbuf_4
Xfanout279 _07335_ vssd1 vssd1 vccd1 vccd1 net279 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout664_A net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout285_X net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15643__A2 net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19230__RESET_B net1482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_3502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09736_ ag2.body\[89\] net781 net775 ag2.body\[90\] _04708_ vssd1 vssd1 vccd1 vccd1
+ _04709_ sky130_fd_sc_hd__a221o_1
XANTENNA__20334__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_12__f_clk clknet_3_6_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_12__leaf_clk
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__09858__B1 net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18042__B1 net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15291__B net52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09667_ net917 net914 net921 net910 vssd1 vssd1 vccd1 vccd1 _04640_ sky130_fd_sc_hd__a31o_4
XANTENNA_fanout452_X net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14188__A net999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17396__A2 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1194_X net1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout929_A obsg2.randCord\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11164__X _06137_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09598_ net890 net900 net904 net896 vssd1 vssd1 vccd1 vccd1 _04571_ sky130_fd_sc_hd__or4b_4
XFILLER_0_55_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20484__CLK clknet_leaf_37_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11324__B net1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout717_X net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11560_ obsg2.obstacleArray\[65\] obsg2.obstacleArray\[69\] net513 vssd1 vssd1 vccd1
+ vccd1 _06533_ sky130_fd_sc_hd__mux2_1
XANTENNA__12090__B1 net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_255 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10511_ _05475_ _05478_ _05482_ _05483_ vssd1 vssd1 vccd1 vccd1 _05484_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_68_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17011__B net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1638 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09729__B net1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11491_ net632 _06463_ vssd1 vssd1 vccd1 vccd1 _06464_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_11_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13230_ net286 _07802_ _07803_ net1721 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[383\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_123_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10442_ _04586_ _05412_ _05413_ _05414_ vssd1 vssd1 vccd1 vccd1 _05415_ sky130_fd_sc_hd__and4_1
XFILLER_0_61_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16203__S0 net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13161_ _07772_ net253 _07770_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[346\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16342__S net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10373_ net907 net920 net916 net912 vssd1 vssd1 vccd1 vccd1 _05346_ sky130_fd_sc_hd__and4bb_2
XANTENNA__14651__A net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_2513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_72_2524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_57_2070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10943__A2 _04230_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12112_ net574 _07080_ _07083_ _06647_ vssd1 vssd1 vccd1 vccd1 _07084_ sky130_fd_sc_hd__o211a_1
XFILLER_0_108_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09745__A net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13092_ _07739_ net265 _07737_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[310\]
+ sky130_fd_sc_hd__mux2_1
XANTENNA__11339__X _06312_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12043_ _06690_ _07013_ _07014_ net439 vssd1 vssd1 vccd1 vccd1 _07015_ sky130_fd_sc_hd__a31o_1
XFILLER_0_44_1482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16920_ _04206_ net869 net710 ag2.body\[564\] vssd1 vssd1 vccd1 vccd1 _02599_ sky130_fd_sc_hd__o22a_1
XFILLER_0_121_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16851_ _02522_ _02523_ _02526_ _02527_ _02529_ vssd1 vssd1 vccd1 vccd1 _02530_ sky130_fd_sc_hd__a221o_1
XANTENNA__18724__CLK clknet_leaf_142_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout780 net781 vssd1 vssd1 vccd1 vccd1 net780 sky130_fd_sc_hd__clkbuf_2
Xfanout791 net797 vssd1 vssd1 vccd1 vccd1 net791 sky130_fd_sc_hd__clkbuf_4
X_15802_ ag2.body\[295\] net207 _01640_ ag2.body\[287\] vssd1 vssd1 vccd1 vccd1 _01049_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_85_2907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_85_2918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19570_ clknet_leaf_118_clk net2498 net1388 vssd1 vssd1 vccd1 vccd1 control.body\[816\]
+ sky130_fd_sc_hd__dfrtp_1
X_16782_ net352 _02384_ _02460_ net460 vssd1 vssd1 vccd1 vccd1 _02461_ sky130_fd_sc_hd__o211a_1
XFILLER_0_92_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_85_2929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13994_ ag2.body\[130\] net213 _08160_ ag2.body\[122\] vssd1 vssd1 vccd1 vccd1 _00211_
+ sky130_fd_sc_hd__a22o_1
X_18521_ clknet_leaf_42_clk net1564 net1372 vssd1 vssd1 vccd1 vccd1 control.detect4.Q\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_66_2328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15733_ ag2.body\[345\] net200 _01633_ ag2.body\[337\] vssd1 vssd1 vccd1 vccd1 _00987_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_77_1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_66_2339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12945_ net293 _07667_ _07668_ net1706 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[233\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__14098__A net1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17387__A2 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18452_ _03839_ _03940_ _03823_ vssd1 vssd1 vccd1 vccd1 _03941_ sky130_fd_sc_hd__a21oi_1
X_15664_ ag2.body\[412\] net143 _01625_ ag2.body\[404\] vssd1 vssd1 vccd1 vccd1 _00926_
+ sky130_fd_sc_hd__a22o_1
X_12876_ net339 net311 vssd1 vssd1 vccd1 vccd1 _07639_ sky130_fd_sc_hd__nand2_8
XANTENNA__18874__CLK clknet_leaf_13_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17403_ ag2.body\[47\] net928 vssd1 vssd1 vccd1 vccd1 _03082_ sky130_fd_sc_hd__xor2_1
X_14615_ net987 ag2.body\[57\] vssd1 vssd1 vccd1 vccd1 _08776_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_51_1431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18383_ _03786_ _03798_ vssd1 vssd1 vccd1 vccd1 _03873_ sky130_fd_sc_hd__or2_1
X_11827_ net571 _06798_ _06796_ vssd1 vssd1 vccd1 vccd1 _06799_ sky130_fd_sc_hd__a21oi_1
X_15595_ ag2.body\[478\] net122 _01618_ ag2.body\[470\] vssd1 vssd1 vccd1 vccd1 _00864_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__14070__B2 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17334_ _03011_ _03012_ vssd1 vssd1 vccd1 vccd1 _03013_ sky130_fd_sc_hd__or2_2
XFILLER_0_16_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11758_ net570 _06729_ _06727_ net471 vssd1 vssd1 vccd1 vccd1 _06730_ sky130_fd_sc_hd__a211o_1
X_14546_ net975 ag2.body\[243\] vssd1 vssd1 vccd1 vccd1 _08707_ sky130_fd_sc_hd__nand2_1
XANTENNA__12081__B1 net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_1516 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10709_ ag2.body\[22\] net1078 vssd1 vssd1 vccd1 vccd1 _05682_ sky130_fd_sc_hd__xor2_1
X_17265_ _02939_ _02940_ _02941_ _02943_ vssd1 vssd1 vccd1 vccd1 _02944_ sky130_fd_sc_hd__a211o_1
XFILLER_0_125_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14477_ net981 ag2.body\[442\] vssd1 vssd1 vccd1 vccd1 _08638_ sky130_fd_sc_hd__xor2_1
X_11689_ _06630_ _06659_ _06658_ vssd1 vssd1 vccd1 vccd1 _06661_ sky130_fd_sc_hd__a21oi_4
XANTENNA__12346__A net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkload104 clknet_leaf_54_clk vssd1 vssd1 vccd1 vccd1 clkload104/Y sky130_fd_sc_hd__bufinv_16
X_19004_ clknet_leaf_2_clk img_gen.tracker.next_frame\[442\] net1247 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[442\] sky130_fd_sc_hd__dfrtp_1
X_16216_ net319 _01894_ vssd1 vssd1 vccd1 vccd1 _01895_ sky130_fd_sc_hd__xnor2_1
Xclkload115 clknet_leaf_62_clk vssd1 vssd1 vccd1 vccd1 clkload115/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_126_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13428_ net1979 net647 _07882_ vssd1 vssd1 vccd1 vccd1 _07883_ sky130_fd_sc_hd__nand3_1
XFILLER_0_107_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17196_ ag2.body\[180\] net960 vssd1 vssd1 vccd1 vccd1 _02875_ sky130_fd_sc_hd__xor2_1
Xclkload126 clknet_leaf_84_clk vssd1 vssd1 vccd1 vccd1 clkload126/Y sky130_fd_sc_hd__inv_4
XANTENNA__11187__A2 net1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11041__D1 net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16147_ obsg2.obstacleArray\[18\] obsg2.obstacleArray\[19\] net429 vssd1 vssd1 vccd1
+ vccd1 _01826_ sky130_fd_sc_hd__mux2_1
X_13359_ net228 _07856_ _07857_ net1853 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[459\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_51_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16252__S net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12633__X _07519_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18033__A net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17311__A2 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09655__A net1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_4203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16078_ obsg2.obstacleArray\[110\] obsg2.obstacleArray\[111\] net422 vssd1 vssd1
+ vccd1 vccd1 _01757_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_36_1420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15873__A2 net161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19906_ clknet_leaf_56_clk _00850_ net1458 vssd1 vssd1 vccd1 vccd1 ag2.body\[480\]
+ sky130_fd_sc_hd__dfrtp_4
X_15029_ control.body\[983\] net167 _01555_ net2492 vssd1 vssd1 vccd1 vccd1 _00361_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_100_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_32_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19837_ clknet_leaf_122_clk _00781_ net1414 vssd1 vssd1 vccd1 vccd1 ag2.body\[555\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_78_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput2 gpio_in[25] vssd1 vssd1 vccd1 vccd1 net2 sky130_fd_sc_hd__clkbuf_1
X_19768_ clknet_leaf_16_clk _00712_ net1316 vssd1 vssd1 vccd1 vccd1 control.body\[630\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_78_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14833__B1 _08315_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1200 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09521_ net891 _04493_ net636 vssd1 vssd1 vccd1 vccd1 _04494_ sky130_fd_sc_hd__o21ai_2
XANTENNA__18024__B1 net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18719_ clknet_leaf_142_clk img_gen.tracker.next_frame\[157\] net1261 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[157\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_49_1803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_49_1814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19699_ clknet_leaf_135_clk _00643_ net1307 vssd1 vssd1 vccd1 vccd1 control.body\[689\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_49_1825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16000__B net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09452_ net917 net913 net922 vssd1 vssd1 vccd1 vccd1 _04425_ sky130_fd_sc_hd__nand3_4
XFILLER_0_56_1375 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16586__B1 net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16935__B net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11426__B1_N _04472_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11144__B net1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09383_ sound_gen.osc1.stayCount\[12\] _04364_ net270 vssd1 vssd1 vccd1 vccd1 _04376_
+ sky130_fd_sc_hd__o21ai_1
XANTENNA__18623__RESET_B net1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14061__A1 net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_583 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14061__B2 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout245_A net246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20612_ net1544 vssd1 vssd1 vccd1 vccd1 gpio_oeb[24] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_99_3350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12072__B1 net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_1140 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_3214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_3225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_715 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16373__D net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16889__B2 ag2.body\[213\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20543_ clknet_leaf_105_clk _01408_ _00017_ vssd1 vssd1 vccd1 vccd1 sound_gen.osc1.stayCount\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout412_A _01902_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10328__X _05301_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15010__B1 _01552_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1154_A net1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20474_ clknet_leaf_33_clk _01361_ net1346 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[110\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__17766__B _03230_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15838__Y _01644_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout200_X net200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10386__B1 _05358_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1419_A net1435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16510__A0 obsg2.obstacleArray\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09565__A net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout781_A net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12127__B2 net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout879_A net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_3029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10063__X _05036_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1008 net1009 vssd1 vssd1 vccd1 vccd1 net1008 sky130_fd_sc_hd__buf_4
XANTENNA__20387__RESET_B net1374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10504__A net1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1019 ag2.randCord\[6\] vssd1 vssd1 vccd1 vccd1 net1019 sky130_fd_sc_hd__buf_4
XANTENNA_fanout1207_X net1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1081 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11886__B1 net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout667_X net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10223__B net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout60_A net61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13534__B _07807_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09719_ ag2.body\[243\] net770 net761 ag2.body\[244\] _04691_ vssd1 vssd1 vccd1 vccd1
+ _04692_ sky130_fd_sc_hd__o221a_1
XANTENNA_fanout834_X net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10991_ ag2.body\[337\] net1211 vssd1 vssd1 vccd1 vccd1 _05964_ sky130_fd_sc_hd__xor2_1
XANTENNA__11102__A2 net1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17721__S _01728_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11335__A net1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12730_ net258 _07568_ _07569_ net1734 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[118\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_38_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16845__B net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12661_ net629 net440 net473 net571 vssd1 vssd1 vccd1 vccd1 _07535_ sky130_fd_sc_hd__and4_2
XANTENNA__14052__A1 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14052__B2 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11612_ obsg2.obstacleArray\[56\] obsg2.obstacleArray\[57\] obsg2.obstacleArray\[60\]
+ obsg2.obstacleArray\[61\] net1125 net511 vssd1 vssd1 vccd1 vccd1 _06585_ sky130_fd_sc_hd__mux4_1
X_14400_ _08559_ _08560_ vssd1 vssd1 vccd1 vccd1 _08561_ sky130_fd_sc_hd__nand2_1
XFILLER_0_77_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12063__B1 net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12592_ net276 net308 _07495_ _07496_ net1749 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[53\]
+ sky130_fd_sc_hd__a32o_1
X_15380_ net2292 net70 _01594_ net2428 vssd1 vssd1 vccd1 vccd1 _00673_ sky130_fd_sc_hd__a22o_1
XFILLER_0_37_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_78_2700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14331_ net998 ag2.body\[424\] vssd1 vssd1 vccd1 vccd1 _08492_ sky130_fd_sc_hd__xnor2_1
X_11543_ obsg2.obstacleArray\[106\] net633 net509 obsg2.obstacleArray\[110\] net759
+ vssd1 vssd1 vccd1 vccd1 _06516_ sky130_fd_sc_hd__o221a_1
XFILLER_0_93_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_2711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10238__X _05211_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_2110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17541__A2 net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_394 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_59_2121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14262_ net981 ag2.body\[10\] vssd1 vssd1 vccd1 vccd1 _08423_ sky130_fd_sc_hd__xor2_1
X_17050_ _04086_ net875 net854 _04088_ vssd1 vssd1 vccd1 vccd1 _02729_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_59_2132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11474_ ag2.body\[491\] net1162 vssd1 vssd1 vccd1 vccd1 _06447_ sky130_fd_sc_hd__nand2_1
XFILLER_0_123_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xwire477 _05999_ vssd1 vssd1 vccd1 vccd1 net477 sky130_fd_sc_hd__clkbuf_2
X_16001_ net871 net939 vssd1 vssd1 vccd1 vccd1 _01680_ sky130_fd_sc_hd__xor2_1
X_13213_ net383 _07627_ vssd1 vssd1 vccd1 vccd1 _07796_ sky130_fd_sc_hd__nor2_1
XFILLER_0_81_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10425_ _05391_ _05395_ _05396_ _05397_ vssd1 vssd1 vccd1 vccd1 _05398_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_55_2007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14193_ net1037 ag2.body\[164\] vssd1 vssd1 vccd1 vccd1 _08354_ sky130_fd_sc_hd__xor2_1
XFILLER_0_106_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_850 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09746__Y _04719_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13144_ net278 _07762_ _07763_ net1950 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[338\]
+ sky130_fd_sc_hd__a22o_1
X_10356_ ag2.body\[291\] net772 _05326_ _05327_ _05328_ vssd1 vssd1 vccd1 vccd1 _05329_
+ sky130_fd_sc_hd__a2111o_1
XANTENNA__15300__A_N _04968_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1280 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_1122 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12613__B _06639_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12118__B2 net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17952_ net380 net462 net495 net481 vssd1 vssd1 vccd1 vccd1 _03579_ sky130_fd_sc_hd__and4_2
X_13075_ net290 _07729_ _07730_ net1739 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[302\]
+ sky130_fd_sc_hd__a22o_1
X_10287_ _05256_ _05257_ _05258_ _05259_ vssd1 vssd1 vccd1 vccd1 _05260_ sky130_fd_sc_hd__a22o_1
X_12026_ img_gen.tracker.frame\[204\] net630 net566 _06997_ vssd1 vssd1 vccd1 vccd1
+ _06998_ sky130_fd_sc_hd__a211o_1
X_16903_ ag2.body\[246\] net943 vssd1 vssd1 vccd1 vccd1 _02582_ sky130_fd_sc_hd__or2_1
XANTENNA__20057__RESET_B net1502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17883_ obsg2.obstacleCount\[1\] obsg2.obstacleCount\[0\] vssd1 vssd1 vccd1 vccd1
+ _03523_ sky130_fd_sc_hd__xor2_4
XANTENNA__16265__C1 net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11341__A2 _04239_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19622_ clknet_leaf_123_clk _00566_ net1407 vssd1 vssd1 vccd1 vccd1 control.body\[772\]
+ sky130_fd_sc_hd__dfrtp_1
X_16834_ ag2.body\[103\] net932 vssd1 vssd1 vccd1 vccd1 _02513_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_73_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19553_ clknet_leaf_115_clk _00497_ net1397 vssd1 vssd1 vccd1 vccd1 control.body\[847\]
+ sky130_fd_sc_hd__dfrtp_1
X_16765_ obsg2.obstacleArray\[4\] net493 net488 obsg2.obstacleArray\[6\] vssd1 vssd1
+ vccd1 vccd1 _02444_ sky130_fd_sc_hd__a22o_1
X_13977_ ag2.body\[115\] net190 _08158_ ag2.body\[107\] vssd1 vssd1 vccd1 vccd1 _00196_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_87_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1624 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18504_ net1515 net1509 vssd1 vssd1 vccd1 vccd1 _00035_ sky130_fd_sc_hd__or2_1
XFILLER_0_57_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15716_ ag2.body\[363\] net193 _01630_ ag2.body\[355\] vssd1 vssd1 vccd1 vccd1 _00973_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_53_1515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19484_ clknet_leaf_114_clk _00428_ net1398 vssd1 vssd1 vccd1 vccd1 control.body\[906\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13163__C _07638_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12928_ net290 _07659_ _07660_ net2033 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[224\]
+ sky130_fd_sc_hd__a22o_1
X_16696_ obsg2.obstacleArray\[64\] net493 net484 obsg2.obstacleArray\[65\] _02374_
+ vssd1 vssd1 vccd1 vccd1 _02375_ sky130_fd_sc_hd__a221o_1
XFILLER_0_92_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_17_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18435_ _03808_ _03911_ _03794_ vssd1 vssd1 vccd1 vccd1 _03924_ sky130_fd_sc_hd__a21oi_1
XANTENNA__19052__CLK clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15647_ ag2.body\[429\] net126 _01623_ ag2.body\[421\] vssd1 vssd1 vccd1 vccd1 _00911_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_29_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16247__S net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12859_ _07431_ _07630_ vssd1 vssd1 vccd1 vccd1 _07631_ sky130_fd_sc_hd__nor2_1
XANTENNA__18309__A1 track.nextHighScore\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18028__A net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15240__B1 _01578_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13460__A _07587_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18366_ _03794_ _03851_ vssd1 vssd1 vccd1 vccd1 _03860_ sky130_fd_sc_hd__nand2_1
XANTENNA__11899__B net1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15578_ _04429_ net64 vssd1 vssd1 vccd1 vccd1 _01616_ sky130_fd_sc_hd__and2_2
XFILLER_0_111_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17317_ ag2.body\[217\] net874 vssd1 vssd1 vccd1 vccd1 _02996_ sky130_fd_sc_hd__xor2_1
XFILLER_0_56_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14529_ net1010 ag2.body\[255\] vssd1 vssd1 vccd1 vccd1 _08690_ sky130_fd_sc_hd__or2_1
X_18297_ track.nextHighScore\[6\] track.nextHighScore\[7\] vssd1 vssd1 vccd1 vccd1
+ _03793_ sky130_fd_sc_hd__or2_2
XFILLER_0_86_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19922__RESET_B net1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17248_ _02924_ _02926_ vssd1 vssd1 vccd1 vccd1 _02927_ sky130_fd_sc_hd__nand2_1
XFILLER_0_113_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17586__B net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17179_ ag2.body\[456\] net737 net696 ag2.body\[462\] _02857_ vssd1 vssd1 vccd1 vccd1
+ _02858_ sky130_fd_sc_hd__a221o_1
XANTENNA__14291__A net996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11565__C1 net1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20190_ clknet_leaf_88_clk _01134_ net1459 vssd1 vssd1 vccd1 vccd1 ag2.body\[204\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_45_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08952_ ag2.body\[11\] vssd1 vssd1 vccd1 vccd1 _03977_ sky130_fd_sc_hd__inv_2
XANTENNA__16710__S net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20480__RESET_B net1355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11139__B net1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11868__B1 net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout195_A net196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18210__B net40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17752__D _02994_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16011__A net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14282__A1 net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout362_A _02222_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14282__B2 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09504_ _04142_ net1209 net757 ag2.body\[405\] vssd1 vssd1 vccd1 vccd1 _04477_ sky130_fd_sc_hd__a22o_1
XFILLER_0_71_1615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09435_ ag2.body\[6\] net1079 vssd1 vssd1 vccd1 vccd1 _04408_ sky130_fd_sc_hd__xor2_1
XANTENNA__10994__A ag2.body\[339\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout627_A net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1369_A net1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09366_ sound_gen.osc1.stayCount\[19\] sound_gen.osc1.stayCount\[18\] _04367_ vssd1
+ vssd1 vccd1 vccd1 _04368_ sky130_fd_sc_hd__and3_1
XANTENNA__12045__B1 net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19545__CLK clknet_leaf_115_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15996__S net223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09297_ sound_gen.osc1.count\[7\] _04308_ _04309_ sound_gen.osc1.count\[6\] _04316_
+ vssd1 vssd1 vccd1 vccd1 _04317_ sky130_fd_sc_hd__o221a_1
XANTENNA__09461__A1 net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout415_X net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17523__A2 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1157_X net1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20526_ clknet_leaf_114_clk _01391_ net1398 vssd1 vssd1 vccd1 vccd1 toggle1.bcd_tens\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__20522__CLK clknet_leaf_93_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16731__B1 net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout996_A net1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20457_ clknet_leaf_38_clk _01344_ net1354 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[93\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout1324_X net1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_628 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10210_ net1161 control.body\[995\] vssd1 vssd1 vccd1 vccd1 _05183_ sky130_fd_sc_hd__nand2_1
XFILLER_0_30_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11190_ _05921_ _06159_ _06161_ _06162_ vssd1 vssd1 vccd1 vccd1 _06163_ sky130_fd_sc_hd__or4_4
XFILLER_0_101_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13529__B _07807_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20388_ clknet_leaf_42_clk _01275_ net1371 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[24\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA_fanout784_X net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16495__C1 net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17716__S net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10141_ net1171 control.body\[818\] vssd1 vssd1 vccd1 vccd1 _05114_ sky130_fd_sc_hd__xor2_1
XFILLER_0_30_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13848__B2 net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11049__B net1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10072_ net1096 control.body\[717\] vssd1 vssd1 vccd1 vccd1 _05045_ sky130_fd_sc_hd__xor2_1
XANTENNA_fanout951_X net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20150__RESET_B net1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13900_ ag2.body\[47\] net118 _08149_ ag2.body\[39\] vssd1 vssd1 vccd1 vccd1 _00128_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__09742__B net1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10521__X _05494_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14880_ control.body\[1107\] net179 _01538_ net2317 vssd1 vssd1 vccd1 vccd1 _00229_
+ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout63_X net63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13831_ _08121_ _08126_ vssd1 vssd1 vccd1 vccd1 _08128_ sky130_fd_sc_hd__and2b_1
XFILLER_0_138_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16550_ obsg2.obstacleArray\[103\] net449 vssd1 vssd1 vccd1 vccd1 _02229_ sky130_fd_sc_hd__or2_1
XFILLER_0_35_1212 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13762_ img_gen.updater.commands.count\[5\] _08075_ _08065_ vssd1 vssd1 vccd1 vccd1
+ _08078_ sky130_fd_sc_hd__o21ai_1
X_10974_ net1108 control.body\[1005\] vssd1 vssd1 vccd1 vccd1 _05947_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_98_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16014__A2 net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15501_ ag2.body\[555\] net113 _01607_ ag2.body\[547\] vssd1 vssd1 vccd1 vccd1 _00781_
+ sky130_fd_sc_hd__a22o_1
X_12713_ net284 _07559_ _07560_ net1650 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[110\]
+ sky130_fd_sc_hd__a22o_1
X_16481_ obsg2.obstacleArray\[36\] obsg2.obstacleArray\[37\] net453 vssd1 vssd1 vccd1
+ vccd1 _02160_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_1644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16067__S net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13693_ _08032_ _08034_ vssd1 vssd1 vccd1 vccd1 _08035_ sky130_fd_sc_hd__nor2_2
XFILLER_0_57_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18220_ _03662_ net40 vssd1 vssd1 vccd1 vccd1 _03749_ sky130_fd_sc_hd__nor2_1
XFILLER_0_35_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12036__B1 net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15432_ ag2.body\[622\] net84 _01599_ ag2.body\[614\] vssd1 vssd1 vccd1 vccd1 _00720_
+ sky130_fd_sc_hd__a22o_1
X_12644_ net264 _07524_ _07525_ net1836 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[76\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__16970__B1 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_931 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_1592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12608__B _07444_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18151_ net523 _03714_ vssd1 vssd1 vccd1 vccd1 _01323_ sky130_fd_sc_hd__and2_1
X_15363_ _05871_ net53 vssd1 vssd1 vccd1 vccd1 _01593_ sky130_fd_sc_hd__nor2_4
X_12575_ net343 net311 _07487_ vssd1 vssd1 vccd1 vccd1 _07488_ sky130_fd_sc_hd__and3_1
XANTENNA__18135__X _03706_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18912__CLK clknet_leaf_142_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17514__A2 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17102_ ag2.body\[8\] net882 vssd1 vssd1 vccd1 vccd1 _02781_ sky130_fd_sc_hd__or2_1
XANTENNA__11795__C1 net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14314_ net832 ag2.body\[49\] _03992_ net980 _08474_ vssd1 vssd1 vccd1 vccd1 _08475_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_48_1617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11526_ obsg2.obstacleArray\[122\] net633 net509 obsg2.obstacleArray\[126\] net759
+ vssd1 vssd1 vccd1 vccd1 _06499_ sky130_fd_sc_hd__o221a_1
X_18082_ net39 _03670_ vssd1 vssd1 vccd1 vccd1 _03671_ sky130_fd_sc_hd__and2_1
XANTENNA__15919__B net61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16722__B1 net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15294_ net2482 net78 _01585_ control.body\[730\] vssd1 vssd1 vccd1 vccd1 _00596_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_53_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17033_ _02706_ _02708_ _02709_ _02711_ vssd1 vssd1 vccd1 vccd1 _02712_ sky130_fd_sc_hd__or4_1
X_11457_ ag2.body\[263\] net1066 vssd1 vssd1 vccd1 vccd1 _06430_ sky130_fd_sc_hd__nand2_1
XFILLER_0_22_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14245_ net1002 ag2.body\[536\] vssd1 vssd1 vccd1 vccd1 _08406_ sky130_fd_sc_hd__xor2_1
XFILLER_0_40_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11547__C1 _06497_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10408_ net1230 control.body\[1072\] vssd1 vssd1 vccd1 vccd1 _05381_ sky130_fd_sc_hd__xor2_1
X_14176_ net982 ag2.body\[194\] vssd1 vssd1 vccd1 vccd1 _08337_ sky130_fd_sc_hd__or2_1
XANTENNA__17278__B2 net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11388_ net1097 control.body\[645\] vssd1 vssd1 vccd1 vccd1 _06361_ sky130_fd_sc_hd__or2_1
X_10339_ _05308_ _05309_ _05310_ _05311_ vssd1 vssd1 vccd1 vccd1 _05312_ sky130_fd_sc_hd__a22o_1
X_13127_ net343 _07587_ vssd1 vssd1 vccd1 vccd1 _07755_ sky130_fd_sc_hd__nor2_1
X_18984_ clknet_leaf_8_clk img_gen.tracker.next_frame\[422\] net1270 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[422\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__13839__A1 net1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17935_ net484 _03540_ _03561_ vssd1 vssd1 vccd1 vccd1 _03566_ sky130_fd_sc_hd__and3_2
X_13058_ net293 _07720_ _07721_ net1840 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[293\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__19418__CLK clknet_leaf_111_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12511__A1 net226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1350 net1351 vssd1 vssd1 vccd1 vccd1 net1350 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12997__C _07515_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12009_ img_gen.tracker.frame\[457\] net614 net540 img_gen.tracker.frame\[463\] _06980_
+ vssd1 vssd1 vccd1 vccd1 _06981_ sky130_fd_sc_hd__o221a_1
XANTENNA__13455__A _07584_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1361 net1362 vssd1 vssd1 vccd1 vccd1 net1361 sky130_fd_sc_hd__clkbuf_4
X_17866_ net2192 _03502_ vssd1 vssd1 vccd1 vccd1 _01239_ sky130_fd_sc_hd__xnor2_1
Xfanout1372 net1373 vssd1 vssd1 vccd1 vccd1 net1372 sky130_fd_sc_hd__clkbuf_4
XANTENNA__16789__B1 net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10522__B1 _05489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1383 net1505 vssd1 vssd1 vccd1 vccd1 net1383 sky130_fd_sc_hd__clkbuf_2
XANTENNA__10798__B net1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1394 net1395 vssd1 vssd1 vccd1 vccd1 net1394 sky130_fd_sc_hd__clkbuf_4
X_16817_ _04011_ net887 net935 _04015_ vssd1 vssd1 vccd1 vccd1 _02496_ sky130_fd_sc_hd__o22a_1
XFILLER_0_108_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13174__B _07607_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19605_ clknet_leaf_120_clk _00549_ net1394 vssd1 vssd1 vccd1 vccd1 control.body\[787\]
+ sky130_fd_sc_hd__dfrtp_1
X_17797_ _04261_ net703 net696 net690 vssd1 vssd1 vccd1 vccd1 _03469_ sky130_fd_sc_hd__or4_1
XANTENNA__13067__A2 _07726_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19536_ clknet_leaf_120_clk _00480_ net1394 vssd1 vssd1 vccd1 vccd1 control.body\[862\]
+ sky130_fd_sc_hd__dfrtp_1
X_16748_ obsg2.obstacleArray\[59\] net501 net487 obsg2.obstacleArray\[58\] _02426_
+ vssd1 vssd1 vccd1 vccd1 _02427_ sky130_fd_sc_hd__a221o_1
XFILLER_0_88_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19467_ clknet_leaf_110_clk _00411_ net1417 vssd1 vssd1 vccd1 vccd1 control.body\[921\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_124_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16679_ net396 _02353_ _02354_ _02355_ net362 vssd1 vssd1 vccd1 vccd1 _02358_ sky130_fd_sc_hd__a221o_1
XANTENNA__14016__A1 net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14016__B2 net1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13190__A net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09220_ control.body\[880\] vssd1 vssd1 vccd1 vccd1 _04245_ sky130_fd_sc_hd__inv_2
X_18418_ _04639_ _03821_ _03848_ vssd1 vssd1 vccd1 vccd1 _03908_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_57_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20545__CLK clknet_leaf_105_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19398_ clknet_leaf_103_clk _00342_ net1427 vssd1 vssd1 vccd1 vccd1 control.body\[996\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_118_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12578__A1 net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09151_ ag2.body\[484\] vssd1 vssd1 vccd1 vccd1 _04176_ sky130_fd_sc_hd__inv_2
XFILLER_0_17_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18592__CLK clknet_leaf_13_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18349_ _03844_ vssd1 vssd1 vccd1 vccd1 _03845_ sky130_fd_sc_hd__inv_2
XFILLER_0_90_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17505__A2 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09667__X _04640_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09082_ ag2.body\[318\] vssd1 vssd1 vccd1 vccd1 _04107_ sky130_fd_sc_hd__inv_2
XFILLER_0_128_1431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20311_ clknet_leaf_44_clk _01211_ net1380 vssd1 vssd1 vccd1 vccd1 ag2.randCord\[5\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_86_1187 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold800 control.body\[641\] vssd1 vssd1 vccd1 vccd1 net2362 sky130_fd_sc_hd__dlygate4sd3_1
Xhold811 _00553_ vssd1 vssd1 vccd1 vccd1 net2373 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12534__A net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold822 control.body\[980\] vssd1 vssd1 vccd1 vccd1 net2384 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11002__A1 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20242_ clknet_leaf_69_clk _01186_ net1496 vssd1 vssd1 vccd1 vccd1 ag2.body\[144\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_130_948 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold833 control.body\[788\] vssd1 vssd1 vccd1 vccd1 net2395 sky130_fd_sc_hd__dlygate4sd3_1
Xhold844 control.body\[1048\] vssd1 vssd1 vccd1 vccd1 net2406 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold855 _00691_ vssd1 vssd1 vccd1 vccd1 net2417 sky130_fd_sc_hd__dlygate4sd3_1
Xhold866 control.body\[663\] vssd1 vssd1 vccd1 vccd1 net2428 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold877 control.body\[777\] vssd1 vssd1 vccd1 vccd1 net2439 sky130_fd_sc_hd__dlygate4sd3_1
X_20173_ clknet_leaf_82_clk _01117_ net1480 vssd1 vssd1 vccd1 vccd1 ag2.body\[219\]
+ sky130_fd_sc_hd__dfrtp_4
Xhold888 control.body\[740\] vssd1 vssd1 vccd1 vccd1 net2450 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold899 control.body\[828\] vssd1 vssd1 vccd1 vccd1 net2461 sky130_fd_sc_hd__dlygate4sd3_1
X_09984_ net1111 control.body\[1117\] vssd1 vssd1 vccd1 vccd1 _04957_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout1117_A ag2.x\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08935_ control.divider.fsm.current_mode\[2\] vssd1 vssd1 vccd1 vccd1 _03960_ sky130_fd_sc_hd__inv_2
XANTENNA__10989__A _04605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16012__Y _01691_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout577_A _06649_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13058__A2 _07720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout365_X net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout744_A _04234_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1486_A net1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_120_3969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout911_A net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16963__X _02642_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15204__B1 _01574_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12709__A net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09418_ obsg2.obstacleCount\[2\] obsg2.obstacleCount\[1\] obsg2.obstacleCount\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04397_ sky130_fd_sc_hd__and3_1
X_10690_ ag2.body\[147\] net1163 vssd1 vssd1 vccd1 vccd1 _05663_ sky130_fd_sc_hd__xor2_1
XFILLER_0_109_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17778__Y _03457_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14558__A2 ag2.body\[70\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12428__B net1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_4_3__f_clk_A clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09349_ _03958_ _04352_ net272 vssd1 vssd1 vccd1 vccd1 _01422_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_8_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_1530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_411 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12360_ _06631_ _07288_ _07296_ _07324_ _07326_ vssd1 vssd1 vccd1 vccd1 _07327_ sky130_fd_sc_hd__a32o_1
XFILLER_0_63_876 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout999_X net999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11311_ ag2.body\[272\] net1232 vssd1 vssd1 vccd1 vccd1 _06284_ sky130_fd_sc_hd__xor2_1
XANTENNA__17794__X _03468_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11792__A2 net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20509_ clknet_leaf_112_clk ag2.goodColl net1424 vssd1 vssd1 vccd1 vccd1 score_detect.N\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_12291_ img_gen.updater.commands.mode\[2\] _07257_ vssd1 vssd1 vccd1 vccd1 _07260_
+ sky130_fd_sc_hd__nand2_1
XANTENNA__10516__X _05489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14030_ _08182_ _08183_ _08189_ _08190_ vssd1 vssd1 vccd1 vccd1 _08191_ sky130_fd_sc_hd__or4b_1
XFILLER_0_47_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11242_ ag2.body\[199\] net1057 vssd1 vssd1 vccd1 vccd1 _06215_ sky130_fd_sc_hd__xor2_1
XFILLER_0_120_447 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1574 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12163__B net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11544__A2 net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12741__A1 net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11173_ net1201 control.body\[777\] vssd1 vssd1 vccd1 vccd1 _06146_ sky130_fd_sc_hd__xor2_1
XFILLER_0_30_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18131__A _03531_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10124_ net1072 control.body\[710\] vssd1 vssd1 vccd1 vccd1 _05097_ sky130_fd_sc_hd__or2_1
X_15981_ _01663_ _01664_ _03964_ vssd1 vssd1 vccd1 vccd1 _01666_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_59_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17720_ _03397_ _03398_ net378 vssd1 vssd1 vccd1 vccd1 _03399_ sky130_fd_sc_hd__mux2_1
X_10055_ ag2.body\[484\] net1138 vssd1 vssd1 vccd1 vccd1 _05028_ sky130_fd_sc_hd__or2_1
X_14932_ net2232 net173 _01544_ net2252 vssd1 vssd1 vccd1 vccd1 _00275_ sky130_fd_sc_hd__a22o_1
X_17651_ ag2.body\[35\] net716 net928 _03986_ _03329_ vssd1 vssd1 vccd1 vccd1 _03330_
+ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_19_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14863_ _08226_ _01524_ _01525_ _01533_ vssd1 vssd1 vccd1 vccd1 _01534_ sky130_fd_sc_hd__and4_1
XANTENNA__14658__X _08819_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14246__B2 net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16602_ obsg2.obstacleArray\[86\] obsg2.obstacleArray\[87\] net447 vssd1 vssd1 vccd1
+ vccd1 _02281_ sky130_fd_sc_hd__mux2_1
X_13814_ control.detect4.Q\[1\] control.detect4.Q\[0\] vssd1 vssd1 vccd1 vccd1 _08111_
+ sky130_fd_sc_hd__nand2b_1
X_17582_ ag2.body\[336\] net741 net878 _04119_ _03260_ vssd1 vssd1 vccd1 vccd1 _03261_
+ sky130_fd_sc_hd__a221o_1
XANTENNA__14797__A2 ag2.body\[291\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14794_ net804 ag2.body\[550\] ag2.body\[551\] net794 _01464_ vssd1 vssd1 vccd1 vccd1
+ _01465_ sky130_fd_sc_hd__a221o_1
XFILLER_0_85_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19321_ clknet_leaf_104_clk _00265_ net1433 vssd1 vssd1 vccd1 vccd1 control.body\[1079\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16533_ _02211_ vssd1 vssd1 vccd1 vccd1 _02212_ sky130_fd_sc_hd__inv_2
XFILLER_0_74_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13745_ net687 _07238_ _08061_ _08062_ vssd1 vssd1 vccd1 vccd1 _08065_ sky130_fd_sc_hd__o211a_1
XANTENNA__13722__B net25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10957_ ag2.body\[174\] net1081 vssd1 vssd1 vccd1 vccd1 _05930_ sky130_fd_sc_hd__nand2_1
XANTENNA__17735__A2 _03251_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12619__A _06639_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19252_ clknet_leaf_75_clk _00196_ net1484 vssd1 vssd1 vccd1 vccd1 ag2.body\[115\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_6_1463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18009__C net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16464_ obsg2.obstacleArray\[58\] obsg2.obstacleArray\[59\] net454 vssd1 vssd1 vccd1
+ vccd1 _02143_ sky130_fd_sc_hd__mux2_1
XANTENNA__15746__A1 ag2.body\[341\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13676_ track.current_collision _07181_ vssd1 vssd1 vccd1 vccd1 _08023_ sky130_fd_sc_hd__nor2_1
X_10888_ net1073 control.body\[654\] vssd1 vssd1 vccd1 vccd1 _05861_ sky130_fd_sc_hd__xor2_1
X_18203_ obsg2.obstacleArray\[98\] _03740_ net521 vssd1 vssd1 vccd1 vccd1 _01349_
+ sky130_fd_sc_hd__o21a_1
XANTENNA__12338__B net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11242__B net1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15415_ control.body\[639\] net81 _01597_ control.body\[631\] vssd1 vssd1 vccd1 vccd1
+ _00705_ sky130_fd_sc_hd__a22o_1
X_12627_ net336 net328 net316 _07515_ vssd1 vssd1 vccd1 vccd1 _07516_ sky130_fd_sc_hd__or4b_1
X_19183_ clknet_leaf_20_clk _00127_ net1331 vssd1 vssd1 vccd1 vccd1 ag2.body\[46\]
+ sky130_fd_sc_hd__dfrtp_4
X_16395_ _02070_ _02072_ _02073_ net364 vssd1 vssd1 vccd1 vccd1 _02074_ sky130_fd_sc_hd__a22o_1
XFILLER_0_112_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10139__A net1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18134_ _03549_ net41 vssd1 vssd1 vccd1 vccd1 _03705_ sky130_fd_sc_hd__nor2_2
X_15346_ net2364 net71 _01591_ control.body\[680\] vssd1 vssd1 vccd1 vccd1 _00642_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__09928__A _04818_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12558_ img_gen.tracker.frame\[38\] net660 _07477_ vssd1 vssd1 vccd1 vccd1 _07478_
+ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_130_Left_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18025__B _01713_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11783__A2 net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18065_ obsg2.obstacleArray\[41\] _03659_ net520 vssd1 vssd1 vccd1 vccd1 _01292_
+ sky130_fd_sc_hd__o21a_1
X_11509_ _06480_ _06481_ vssd1 vssd1 vccd1 vccd1 _06482_ sky130_fd_sc_hd__nand2b_2
XTAP_TAPCELL_ROW_130_4276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15277_ control.body\[755\] net88 _01583_ control.body\[747\] vssd1 vssd1 vccd1 vccd1
+ _00581_ sky130_fd_sc_hd__a22o_1
XFILLER_0_79_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold107 img_gen.tracker.frame\[91\] vssd1 vssd1 vccd1 vccd1 net1669 sky130_fd_sc_hd__dlygate4sd3_1
X_12489_ net594 net469 net561 _07312_ vssd1 vssd1 vccd1 vccd1 _07438_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_130_4287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold118 img_gen.tracker.frame\[177\] vssd1 vssd1 vccd1 vccd1 net1680 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_130_4298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17016_ ag2.body\[332\] net966 vssd1 vssd1 vccd1 vccd1 _02695_ sky130_fd_sc_hd__xor2_1
Xhold129 img_gen.tracker.frame\[206\] vssd1 vssd1 vccd1 vccd1 net1691 sky130_fd_sc_hd__dlygate4sd3_1
X_14228_ net980 net971 net1025 net1019 vssd1 vssd1 vccd1 vccd1 _08389_ sky130_fd_sc_hd__or4_1
XFILLER_0_61_1603 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16260__S net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14159_ net806 ag2.body\[621\] ag2.body\[623\] net790 vssd1 vssd1 vccd1 vccd1 _08320_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__18463__A3 net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18041__A net42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout609 net610 vssd1 vssd1 vccd1 vccd1 net609 sky130_fd_sc_hd__clkbuf_4
XANTENNA__18808__CLK clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09663__A net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_14__f_clk_A clknet_3_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18967_ clknet_leaf_5_clk img_gen.tracker.next_frame\[405\] net1269 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[405\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__12801__B _07444_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15682__B1 _01627_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13185__A net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17918_ _03536_ _03551_ vssd1 vssd1 vccd1 vccd1 _03552_ sky130_fd_sc_hd__nor2_1
X_18898_ clknet_leaf_144_clk img_gen.tracker.next_frame\[336\] net1252 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[336\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__10602__A net1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11838__A3 _06809_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19390__CLK clknet_leaf_102_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1180 net1189 vssd1 vssd1 vccd1 vccd1 net1180 sky130_fd_sc_hd__buf_4
Xfanout1191 net1200 vssd1 vssd1 vccd1 vccd1 net1191 sky130_fd_sc_hd__buf_4
XANTENNA__09900__A2 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17849_ img_gen.updater.commands.rR1.rainbowRNG\[12\] img_gen.updater.commands.rR1.rainbowRNG\[11\]
+ _03504_ vssd1 vssd1 vccd1 vccd1 _03505_ sky130_fd_sc_hd__and3_1
XFILLER_0_59_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14237__A1 net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14237__B2 net980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19519_ clknet_leaf_121_clk _00463_ net1401 vssd1 vssd1 vccd1 vccd1 control.body\[877\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__17879__X _03519_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17104__B net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_957 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout158_A net161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20519__Q control.body_update.curr_length\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15737__B2 ag2.body\[341\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19255__RESET_B net1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09203_ net1192 vssd1 vssd1 vccd1 vccd1 _04228_ sky130_fd_sc_hd__inv_2
XFILLER_0_91_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14744__A net1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09134_ ag2.body\[447\] vssd1 vssd1 vccd1 vccd1 _04159_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout1067_A net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09838__A net1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15559__B net56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12420__B1 net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10991__B net1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11579__S net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12971__A1 net233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09065_ ag2.body\[266\] vssd1 vssd1 vccd1 vccd1 _04090_ sky130_fd_sc_hd__inv_2
XANTENNA__10431__C1 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout113_X net113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_3762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1234_A net1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_113_3773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09719__A2 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_3784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17774__B _03442_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold630 img_gen.updater.commands.rR1.rainbowRNG\[8\] vssd1 vssd1 vccd1 vccd1 net2192
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13079__B net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout694_A net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold641 control.body\[1015\] vssd1 vssd1 vccd1 vccd1 net2203 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11526__A2 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold652 control.body\[995\] vssd1 vssd1 vccd1 vccd1 net2214 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12723__A1 net247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_778 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20225_ clknet_leaf_61_clk _01169_ net1469 vssd1 vssd1 vccd1 vccd1 ag2.body\[175\]
+ sky130_fd_sc_hd__dfrtp_4
Xhold663 control.body\[693\] vssd1 vssd1 vccd1 vccd1 net2225 sky130_fd_sc_hd__dlygate4sd3_1
Xhold674 control.body\[968\] vssd1 vssd1 vccd1 vccd1 net2236 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1022_X net1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold685 control.body\[708\] vssd1 vssd1 vccd1 vccd1 net2247 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_1423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold696 _00576_ vssd1 vssd1 vccd1 vccd1 net2258 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20156_ clknet_leaf_96_clk _01100_ net1441 vssd1 vssd1 vccd1 vccd1 ag2.body\[234\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA_fanout861_A net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09967_ ag2.body\[84\] net1138 vssd1 vssd1 vccd1 vccd1 _04940_ sky130_fd_sc_hd__xor2_1
XANTENNA_fanout482_X net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1367 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout959_A net961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17790__A net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13095__A net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20087_ clknet_leaf_76_clk _01031_ net1492 vssd1 vssd1 vccd1 vccd1 ag2.body\[309\]
+ sky130_fd_sc_hd__dfrtp_4
X_09898_ ag2.body\[74\] net1185 vssd1 vssd1 vccd1 vccd1 _04871_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_107_3577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_107_3588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_107_3599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout747_X net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11860_ img_gen.tracker.frame\[205\] net624 net607 img_gen.tracker.frame\[208\] vssd1
+ vssd1 vccd1 vccd1 _06832_ sky130_fd_sc_hd__o22a_1
X_10811_ net1182 control.body\[1090\] vssd1 vssd1 vccd1 vccd1 _05784_ sky130_fd_sc_hd__or2_1
XFILLER_0_131_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17014__B net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11791_ img_gen.tracker.frame\[374\] net621 net587 img_gen.tracker.frame\[383\] _06762_
+ vssd1 vssd1 vccd1 vccd1 _06763_ sky130_fd_sc_hd__o221a_1
XFILLER_0_95_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19113__CLK clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13530_ net2101 net655 _07923_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[564\]
+ sky130_fd_sc_hd__and3_1
X_10742_ ag2.body\[501\] net1114 vssd1 vssd1 vccd1 vccd1 _05715_ sky130_fd_sc_hd__or2_1
XFILLER_0_32_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17949__B net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_2784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_2795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11062__B net1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10673_ ag2.body\[344\] net1235 vssd1 vssd1 vccd1 vccd1 _05646_ sky130_fd_sc_hd__xor2_1
X_13461_ net682 _07896_ vssd1 vssd1 vccd1 vccd1 _07897_ sky130_fd_sc_hd__nor2_1
XANTENNA__16345__S net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12726__X _07567_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15200_ net890 net904 _04758_ _01548_ vssd1 vssd1 vccd1 vccd1 _01574_ sky130_fd_sc_hd__o31a_4
X_12412_ _07318_ _07337_ _07371_ _07374_ vssd1 vssd1 vccd1 vccd1 _07375_ sky130_fd_sc_hd__a211o_1
X_16180_ obsg2.obstacleArray\[36\] obsg2.obstacleArray\[37\] net423 vssd1 vssd1 vccd1
+ vccd1 _01859_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13392_ net388 net382 _07306_ net312 vssd1 vssd1 vccd1 vccd1 _07870_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_11_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18142__A2 net37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15131_ net2586 net103 _01566_ net2249 vssd1 vssd1 vccd1 vccd1 _00452_ sky130_fd_sc_hd__a22o_1
XANTENNA__11765__A2 net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12962__A1 net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17965__A net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12343_ net438 _07305_ vssd1 vssd1 vccd1 vccd1 _07310_ sky130_fd_sc_hd__nand2_1
XFILLER_0_133_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15062_ net2279 net150 _01559_ net2354 vssd1 vssd1 vccd1 vccd1 _00390_ sky130_fd_sc_hd__a22o_1
X_12274_ _07206_ _07241_ _07231_ img_gen.updater.commands.cmd_num\[2\] vssd1 vssd1
+ vccd1 vccd1 _07244_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_107_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18132__Y _03703_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14013_ net825 ag2.body\[458\] _04162_ net1036 _08172_ vssd1 vssd1 vccd1 vccd1 _08174_
+ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_75_2599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11225_ net1149 control.body\[859\] vssd1 vssd1 vccd1 vccd1 _06198_ sky130_fd_sc_hd__xor2_1
XFILLER_0_121_789 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19870_ clknet_leaf_95_clk _00814_ net1440 vssd1 vssd1 vccd1 vccd1 ag2.body\[524\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_120_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18821_ clknet_leaf_5_clk img_gen.tracker.next_frame\[259\] net1269 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[259\] sky130_fd_sc_hd__dfrtp_1
X_11156_ ag2.body\[607\] net1047 vssd1 vssd1 vccd1 vccd1 _06129_ sky130_fd_sc_hd__nand2_1
XFILLER_0_43_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10107_ net1058 control.body\[943\] vssd1 vssd1 vccd1 vccd1 _05080_ sky130_fd_sc_hd__nand2_1
XFILLER_0_65_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18752_ clknet_leaf_143_clk img_gen.tracker.next_frame\[190\] net1256 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[190\] sky130_fd_sc_hd__dfrtp_1
X_15964_ _05239_ net60 vssd1 vssd1 vccd1 vccd1 _01658_ sky130_fd_sc_hd__nor2_2
X_11087_ net1180 ag2.body\[538\] vssd1 vssd1 vccd1 vccd1 _06060_ sky130_fd_sc_hd__and2b_1
X_17703_ obsg2.obstacleArray\[138\] obsg2.obstacleArray\[139\] net410 vssd1 vssd1
+ vccd1 vccd1 _03382_ sky130_fd_sc_hd__mux2_1
X_10038_ net1083 control.body\[902\] vssd1 vssd1 vccd1 vccd1 _05011_ sky130_fd_sc_hd__xor2_1
X_14915_ control.body\[1074\] net171 _01542_ control.body\[1066\] vssd1 vssd1 vccd1
+ vccd1 _00260_ sky130_fd_sc_hd__a22o_1
X_18683_ clknet_leaf_28_clk img_gen.tracker.next_frame\[121\] net1336 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[121\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__11237__B net1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14219__A1 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15895_ ag2.body\[202\] net133 _01650_ ag2.body\[194\] vssd1 vssd1 vccd1 vccd1 _01132_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_136_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_123_4080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14219__B2 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17634_ ag2.body\[164\] net961 vssd1 vssd1 vccd1 vccd1 _03313_ sky130_fd_sc_hd__nand2_1
XFILLER_0_8_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14846_ _08758_ _08762_ _01456_ _01516_ vssd1 vssd1 vccd1 vccd1 _01517_ sky130_fd_sc_hd__o211a_1
XANTENNA__09930__B _04792_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_1451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17565_ ag2.body\[577\] net730 net848 _04211_ vssd1 vssd1 vccd1 vccd1 _03244_ sky130_fd_sc_hd__a22o_1
XFILLER_0_19_1582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14777_ net983 _04093_ ag2.body\[279\] net795 _01447_ vssd1 vssd1 vccd1 vccd1 _01448_
+ sky130_fd_sc_hd__a221o_1
XANTENNA__17708__A2 net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12349__A net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11989_ img_gen.tracker.frame\[400\] net600 net584 img_gen.tracker.frame\[406\] _06960_
+ vssd1 vssd1 vccd1 vccd1 _06961_ sky130_fd_sc_hd__o221a_1
XFILLER_0_54_1473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19304_ clknet_leaf_98_clk net2324 net1446 vssd1 vssd1 vccd1 vccd1 control.body\[1094\]
+ sky130_fd_sc_hd__dfrtp_1
X_16516_ _02184_ _02185_ net402 vssd1 vssd1 vccd1 vccd1 _02195_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13728_ _04318_ sound_gen.osc1.keepCounting_nxt vssd1 vssd1 vccd1 vccd1 sound_gen.osc1.at_max_nxt
+ sky130_fd_sc_hd__and2b_1
XFILLER_0_128_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17496_ _03169_ _03174_ vssd1 vssd1 vccd1 vccd1 _03175_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_15_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_50_clk_A clknet_4_6__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12068__B net1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_136_4463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19235_ clknet_leaf_84_clk _00179_ net1481 vssd1 vssd1 vccd1 vccd1 ag2.body\[98\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_136_4474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16447_ obsg2.obstacleArray\[68\] obsg2.obstacleArray\[69\] net456 vssd1 vssd1 vccd1
+ vccd1 _02126_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_4485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13659_ net998 net989 vssd1 vssd1 vccd1 vccd1 _08013_ sky130_fd_sc_hd__nand2_1
XANTENNA__16255__S net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18036__A net39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14564__A net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_4338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_4349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19166_ clknet_leaf_21_clk _00110_ net1363 vssd1 vssd1 vccd1 vccd1 ag2.body\[29\]
+ sky130_fd_sc_hd__dfrtp_4
X_16378_ _02055_ _02056_ vssd1 vssd1 vccd1 vccd1 _02057_ sky130_fd_sc_hd__nand2b_4
XFILLER_0_42_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__20253__RESET_B net1499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_515 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_1566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18117_ net44 _03693_ vssd1 vssd1 vccd1 vccd1 _03694_ sky130_fd_sc_hd__nor2_1
XANTENNA__11756__A2 _06476_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_1588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15329_ net2343 net73 _01587_ control.body\[697\] vssd1 vssd1 vccd1 vccd1 _00627_
+ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_65_clk_A clknet_4_13__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16144__A1 net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19097_ clknet_leaf_145_clk img_gen.tracker.next_frame\[535\] net1241 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[535\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__14851__X _01522_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18630__CLK clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16695__A2 net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18048_ obsg2.obstacleArray\[35\] _03648_ net521 vssd1 vssd1 vccd1 vccd1 _01286_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_83_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_767 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10316__B net1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_1467 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_3091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12812__A net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout406 net408 vssd1 vssd1 vccd1 vccd1 net406 sky130_fd_sc_hd__buf_2
X_20010_ clknet_leaf_59_clk _00954_ net1467 vssd1 vssd1 vccd1 vccd1 ag2.body\[376\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_1_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout417 _01899_ vssd1 vssd1 vccd1 vccd1 net417 sky130_fd_sc_hd__buf_4
XFILLER_0_26_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09821_ net750 control.body\[1054\] _04793_ vssd1 vssd1 vccd1 vccd1 _04794_ sky130_fd_sc_hd__a21oi_1
Xfanout428 net429 vssd1 vssd1 vccd1 vccd1 net428 sky130_fd_sc_hd__clkbuf_4
XANTENNA__17881__Y _03521_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout439 net440 vssd1 vssd1 vccd1 vccd1 net439 sky130_fd_sc_hd__buf_2
X_19999_ clknet_leaf_66_clk _00943_ net1475 vssd1 vssd1 vccd1 vccd1 ag2.body\[397\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__14458__B2 net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18780__CLK clknet_leaf_13_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09752_ ag2.body\[211\] net1162 vssd1 vssd1 vccd1 vccd1 _04725_ sky130_fd_sc_hd__nand2_1
XANTENNA_clkbuf_leaf_123_clk_A clknet_4_9__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10332__A _04600_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09683_ ag2.body\[8\] net1223 vssd1 vssd1 vccd1 vccd1 _04656_ sky130_fd_sc_hd__xor2_1
XANTENNA__14739__A net1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10051__B net1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout275_A net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19136__CLK clknet_leaf_132_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10495__A2 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_3430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_102_3441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_138_clk_A clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13362__B _07528_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09637__A1 net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout442_A net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14630__A1 net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09637__B2 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1184_A net1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14630__B2 net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_18_clk_A clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout35 net36 vssd1 vssd1 vccd1 vccd1 net35 sky130_fd_sc_hd__clkbuf_4
XANTENNA__17769__B _02837_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16907__B1 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout46 _03591_ vssd1 vssd1 vccd1 vccd1 net46 sky130_fd_sc_hd__clkbuf_4
Xfanout57 net62 vssd1 vssd1 vccd1 vccd1 net57 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_91_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19286__CLK clknet_leaf_98_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout230_X net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout68 net70 vssd1 vssd1 vccd1 vccd1 net68 sky130_fd_sc_hd__buf_2
XANTENNA_fanout1351_A net1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_119_3960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_575 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout79 net91 vssd1 vssd1 vccd1 vccd1 net79 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_68_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout707_A net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout328_X net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1449_A net1451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14394__B1 ag2.body\[122\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_115_3824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_3835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18124__A2 net38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14193__B ag2.body\[164\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_3_5_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20263__CLK clknet_leaf_43_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12944__A1 net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09117_ ag2.body\[401\] vssd1 vssd1 vccd1 vccd1 _04142_ sky130_fd_sc_hd__inv_2
XANTENNA__10507__A net1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1237_X net1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09048_ ag2.body\[237\] vssd1 vssd1 vccd1 vccd1 _04073_ sky130_fd_sc_hd__inv_2
XFILLER_0_108_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14697__A1 net993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10226__B net1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14697__B2 net1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout697_X net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold460 img_gen.tracker.frame\[507\] vssd1 vssd1 vccd1 vccd1 net2022 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12722__A net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1404_X net1404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold471 img_gen.tracker.frame\[224\] vssd1 vssd1 vccd1 vccd1 net2033 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout90_A net91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold482 img_gen.tracker.frame\[83\] vssd1 vssd1 vccd1 vccd1 net2044 sky130_fd_sc_hd__dlygate4sd3_1
X_11010_ net755 control.body\[1085\] control.body\[1086\] net750 vssd1 vssd1 vccd1
+ vccd1 _05983_ sky130_fd_sc_hd__a22o_1
X_20208_ clknet_leaf_56_clk _01152_ net1457 vssd1 vssd1 vccd1 vccd1 ag2.body\[190\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__09573__B1 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold493 img_gen.tracker.frame\[475\] vssd1 vssd1 vccd1 vccd1 net2055 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_70_2452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17009__B net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_2463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout864_X net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15646__B1 _01623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout940 net941 vssd1 vssd1 vccd1 vccd1 net940 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_109_3639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout951 net952 vssd1 vssd1 vccd1 vccd1 net951 sky130_fd_sc_hd__buf_4
X_20139_ clknet_leaf_97_clk _01083_ net1450 vssd1 vssd1 vccd1 vccd1 ag2.body\[249\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_95_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout962 net963 vssd1 vssd1 vccd1 vccd1 net962 sky130_fd_sc_hd__buf_4
Xfanout973 net974 vssd1 vssd1 vccd1 vccd1 net973 sky130_fd_sc_hd__buf_4
Xfanout984 ag2.randCord\[2\] vssd1 vssd1 vccd1 vccd1 net984 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_5_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09453__D net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout995 ag2.randCord\[1\] vssd1 vssd1 vccd1 vccd1 net995 sky130_fd_sc_hd__buf_4
XANTENNA__16848__B net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11057__B net1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_5_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12961_ net254 _07676_ _07677_ net2072 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[241\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__17399__B1 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11132__B1 net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14700_ _08858_ _08860_ vssd1 vssd1 vccd1 vccd1 _08861_ sky130_fd_sc_hd__nand2_1
XFILLER_0_99_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_87_2971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_2982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11912_ img_gen.tracker.frame\[346\] net580 net542 img_gen.tracker.frame\[343\] _06883_
+ vssd1 vssd1 vccd1 vccd1 _06884_ sky130_fd_sc_hd__o221a_1
X_15680_ ag2.body\[394\] net143 _01627_ ag2.body\[386\] vssd1 vssd1 vccd1 vccd1 _00940_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_73_1326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10486__A2 net1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12892_ net681 _07645_ vssd1 vssd1 vccd1 vccd1 _07646_ sky130_fd_sc_hd__nor2_1
XFILLER_0_115_1614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_83_2846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_2392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14631_ _08785_ _08786_ _08789_ _08791_ vssd1 vssd1 vccd1 vccd1 _08792_ sky130_fd_sc_hd__or4b_1
XTAP_TAPCELL_ROW_83_2857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_83_2868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11843_ img_gen.tracker.frame\[521\] net599 net583 img_gen.tracker.frame\[527\] vssd1
+ vssd1 vccd1 vccd1 _06815_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_64_2267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17350_ _03024_ _03028_ _03009_ vssd1 vssd1 vccd1 vccd1 _03029_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_36_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_64_2278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14562_ net1023 ag2.body\[358\] vssd1 vssd1 vccd1 vccd1 _08723_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_64_2289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11774_ _06743_ _06745_ net564 vssd1 vssd1 vccd1 vccd1 _06746_ sky130_fd_sc_hd__mux2_1
X_16301_ obsg2.obstacleArray\[96\] obsg2.obstacleArray\[97\] net404 vssd1 vssd1 vccd1
+ vccd1 _01980_ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13513_ net288 _07612_ _07806_ _07916_ net1714 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[554\]
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_51_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10725_ net643 _05697_ vssd1 vssd1 vccd1 vccd1 _05698_ sky130_fd_sc_hd__nor2_2
X_17281_ _02952_ _02953_ _02958_ _02959_ vssd1 vssd1 vccd1 vccd1 _02960_ sky130_fd_sc_hd__or4_1
X_14493_ _08648_ _08649_ _08652_ _08653_ vssd1 vssd1 vccd1 vccd1 _08654_ sky130_fd_sc_hd__or4_2
XANTENNA__14384__A net1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13188__A1 net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19020_ clknet_leaf_2_clk img_gen.tracker.next_frame\[458\] net1247 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[458\] sky130_fd_sc_hd__dfrtp_1
X_16232_ net463 _01905_ vssd1 vssd1 vccd1 vccd1 _01911_ sky130_fd_sc_hd__xnor2_2
XANTENNA__18653__CLK clknet_leaf_131_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1108 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13444_ net282 _07888_ _07889_ net1724 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[512\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__19779__CLK clknet_leaf_127_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10656_ ag2.body\[281\] net1212 vssd1 vssd1 vccd1 vccd1 _05629_ sky130_fd_sc_hd__xor2_1
XANTENNA__12175__Y _07147_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11738__A2 net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16163_ obsg2.obstacleArray\[8\] net426 net374 _01841_ vssd1 vssd1 vccd1 vccd1 _01842_
+ sky130_fd_sc_hd__o211a_1
Xclkload16 clknet_leaf_6_clk vssd1 vssd1 vccd1 vccd1 clkload16/Y sky130_fd_sc_hd__bufinv_16
X_10587_ net1051 control.body\[831\] vssd1 vssd1 vccd1 vccd1 _05560_ sky130_fd_sc_hd__nand2_1
Xclkload27 clknet_leaf_132_clk vssd1 vssd1 vccd1 vccd1 clkload27/X sky130_fd_sc_hd__clkbuf_8
X_13375_ net255 _07862_ _07863_ net1683 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[469\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_49_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkload38 clknet_leaf_19_clk vssd1 vssd1 vccd1 vccd1 clkload38/Y sky130_fd_sc_hd__inv_16
Xclkload49 clknet_leaf_31_clk vssd1 vssd1 vccd1 vccd1 clkload49/Y sky130_fd_sc_hd__inv_12
X_15114_ control.body\[899\] net146 _01554_ net2544 vssd1 vssd1 vccd1 vccd1 _00437_
+ sky130_fd_sc_hd__a22o_1
X_12326_ _07255_ _07292_ vssd1 vssd1 vccd1 vccd1 _07293_ sky130_fd_sc_hd__nand2_1
XFILLER_0_49_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16094_ obsg2.obstacleArray\[118\] net425 vssd1 vssd1 vccd1 vccd1 _01773_ sky130_fd_sc_hd__or2_1
XFILLER_0_80_1319 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14688__A1 net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14688__B2 net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19922_ clknet_leaf_51_clk _00866_ net1368 vssd1 vssd1 vccd1 vccd1 ag2.body\[464\]
+ sky130_fd_sc_hd__dfrtp_4
X_15045_ control.body\[965\] net165 _01556_ net2375 vssd1 vssd1 vccd1 vccd1 _00375_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__09925__B net1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12257_ _07195_ _07226_ _07204_ vssd1 vssd1 vccd1 vccd1 _07227_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_76_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12632__A net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13360__A1 net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11208_ _04446_ _05051_ vssd1 vssd1 vccd1 vccd1 _06181_ sky130_fd_sc_hd__nor2_1
X_12188_ net1102 ag2.apple_cord\[5\] vssd1 vssd1 vccd1 vccd1 _07160_ sky130_fd_sc_hd__nand2_1
X_19853_ clknet_leaf_92_clk _00797_ net1413 vssd1 vssd1 vccd1 vccd1 ag2.body\[539\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_43_1185 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_125_4131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11910__A2 net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_4142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18804_ clknet_leaf_3_clk img_gen.tracker.next_frame\[242\] net1259 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[242\] sky130_fd_sc_hd__dfrtp_1
X_11139_ ag2.body\[410\] net1176 vssd1 vssd1 vccd1 vccd1 _06112_ sky130_fd_sc_hd__xor2_1
XFILLER_0_120_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19159__CLK clknet_leaf_52_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16996_ ag2.body\[143\] net934 vssd1 vssd1 vccd1 vccd1 _02675_ sky130_fd_sc_hd__xor2_1
X_19784_ clknet_leaf_127_clk _00728_ net1331 vssd1 vssd1 vccd1 vccd1 ag2.body\[614\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_121_4006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_34_1370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15947_ ag2.body\[152\] net195 _01656_ ag2.body\[144\] vssd1 vssd1 vccd1 vccd1 _01178_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_121_4028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18735_ clknet_leaf_143_clk img_gen.tracker.next_frame\[173\] net1257 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[173\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_1494 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09660__B net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10477__A2 _04446_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18666_ clknet_leaf_11_clk img_gen.tracker.next_frame\[104\] net1282 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[104\] sky130_fd_sc_hd__dfrtp_1
X_15878_ ag2.body\[219\] net188 _01648_ ag2.body\[211\] vssd1 vssd1 vccd1 vccd1 _01117_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__16601__A2 net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14829_ _08650_ _08654_ _01478_ _08635_ _08613_ vssd1 vssd1 vccd1 vccd1 _01500_ sky130_fd_sc_hd__o2111a_1
XANTENNA__13182__B net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17617_ ag2.body\[603\] net715 net698 ag2.body\[606\] vssd1 vssd1 vccd1 vccd1 _03296_
+ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_138_4525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18597_ clknet_leaf_13_clk img_gen.tracker.next_frame\[35\] net1282 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[35\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_138_4536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_1753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17548_ _04111_ net967 net694 ag2.body\[327\] vssd1 vssd1 vccd1 vccd1 _03227_ sky130_fd_sc_hd__a22o_1
XANTENNA__11426__A1 _04556_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_4569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11977__A2 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13910__B net57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17479_ ag2.body\[134\] net944 vssd1 vssd1 vccd1 vccd1 _03158_ sky130_fd_sc_hd__nand2_1
XFILLER_0_73_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12807__A net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13179__A1 net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_15_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19218_ clknet_leaf_67_clk _00162_ net1494 vssd1 vssd1 vccd1 vccd1 ag2.body\[81\]
+ sky130_fd_sc_hd__dfrtp_4
X_20490_ clknet_leaf_38_clk _01377_ net1353 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[126\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_15_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14915__A2 net171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_982 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12526__B net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11729__A2 net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11430__B net1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19149_ clknet_leaf_50_clk _00093_ net1367 vssd1 vssd1 vccd1 vccd1 ag2.body\[13\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_6_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17314__B1 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16713__S net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_3153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_93_3164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16668__A2 net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10614__X _05587_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout203 net204 vssd1 vssd1 vccd1 vccd1 net203 sky130_fd_sc_hd__clkbuf_2
Xfanout214 net218 vssd1 vssd1 vccd1 vccd1 net214 sky130_fd_sc_hd__clkbuf_2
XANTENNA__13357__B _07523_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout392_A net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout225 net227 vssd1 vssd1 vccd1 vccd1 net225 sky130_fd_sc_hd__buf_4
XANTENNA__15628__B1 _01621_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1304 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout236 net247 vssd1 vssd1 vccd1 vccd1 net236 sky130_fd_sc_hd__buf_2
X_09804_ net1181 control.body\[962\] vssd1 vssd1 vccd1 vccd1 _04777_ sky130_fd_sc_hd__nand2_1
XANTENNA__11901__A2 net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout247 _07331_ vssd1 vssd1 vccd1 vccd1 net247 sky130_fd_sc_hd__buf_4
Xfanout258 net259 vssd1 vssd1 vccd1 vccd1 net258 sky130_fd_sc_hd__clkbuf_4
Xfanout269 _07303_ vssd1 vssd1 vccd1 vccd1 net269 sky130_fd_sc_hd__buf_2
XANTENNA__13103__A1 net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_3503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09735_ _04017_ net1210 net1114 _04020_ vssd1 vssd1 vccd1 vccd1 _04708_ sky130_fd_sc_hd__a22o_1
XFILLER_0_39_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14469__A net1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09858__A1 net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11592__S net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout278_X net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13373__A net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09666_ _04425_ _04637_ vssd1 vssd1 vccd1 vccd1 _04639_ sky130_fd_sc_hd__nand2_4
XANTENNA__14188__B ag2.body\[160\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14603__A1 net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout445_X net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout824_A net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09597_ _04540_ _04543_ _04549_ _04569_ vssd1 vssd1 vccd1 vccd1 _04570_ sky130_fd_sc_hd__o31a_1
XANTENNA__14603__B2 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1187_X net1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17499__B net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_510 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11968__A2 net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13820__B _08114_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout612_X net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_143_clk clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_143_clk
+ sky130_fd_sc_hd__clkbuf_8
X_10510_ net769 control.body\[979\] control.body\[981\] net755 vssd1 vssd1 vccd1 vccd1
+ _05483_ sky130_fd_sc_hd__o22a_1
XFILLER_0_64_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11490_ net1222 net1102 vssd1 vssd1 vccd1 vccd1 _06463_ sky130_fd_sc_hd__and2b_2
X_10441_ net1107 control.body\[933\] vssd1 vssd1 vccd1 vccd1 _05414_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_33_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17719__S net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17946__C _03574_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_2650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16203__S1 net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13160_ img_gen.tracker.frame\[346\] net646 vssd1 vssd1 vccd1 vccd1 _07772_ sky130_fd_sc_hd__and2_1
X_10372_ net767 control.body\[763\] _05342_ _05343_ _05344_ vssd1 vssd1 vccd1 vccd1
+ _05345_ sky130_fd_sc_hd__a2111o_1
XANTENNA_fanout981_X net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_72_2514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_2060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_57_2071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12111_ img_gen.tracker.frame\[183\] net610 net563 _07082_ vssd1 vssd1 vccd1 vccd1
+ _07083_ sky130_fd_sc_hd__a211o_1
X_13091_ img_gen.tracker.frame\[310\] net662 vssd1 vssd1 vccd1 vccd1 _07739_ sky130_fd_sc_hd__and2_1
XFILLER_0_32_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09745__B _04421_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1326 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12042_ net470 _07004_ _07007_ vssd1 vssd1 vccd1 vccd1 _07014_ sky130_fd_sc_hd__or3_1
XANTENNA__12145__A2 net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold290 img_gen.tracker.frame\[374\] vssd1 vssd1 vccd1 vccd1 net1852 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_1502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16850_ ag2.body\[168\] net737 net940 _04053_ _02528_ vssd1 vssd1 vccd1 vccd1 _02529_
+ sky130_fd_sc_hd__a221o_1
XANTENNA__17084__A2 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16578__B net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15801_ ag2.body\[294\] net207 _01640_ ag2.body\[286\] vssd1 vssd1 vccd1 vccd1 _01048_
+ sky130_fd_sc_hd__a22o_1
Xfanout770 net771 vssd1 vssd1 vccd1 vccd1 net770 sky130_fd_sc_hd__buf_4
XANTENNA__09761__A ag2.body\[209\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout781 net782 vssd1 vssd1 vccd1 vccd1 net781 sky130_fd_sc_hd__buf_6
Xfanout792 net797 vssd1 vssd1 vccd1 vccd1 net792 sky130_fd_sc_hd__buf_4
X_16781_ net380 _02414_ _02409_ net350 vssd1 vssd1 vccd1 vccd1 _02460_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_85_2908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13993_ ag2.body\[129\] net213 _08160_ ag2.body\[121\] vssd1 vssd1 vccd1 vccd1 _00210_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_85_2919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09849__A1 _04445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18520_ net1 net9 vssd1 vssd1 vccd1 vccd1 _00051_ sky130_fd_sc_hd__or2_1
XANTENNA__13283__A net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15732_ ag2.body\[344\] net212 _01633_ ag2.body\[336\] vssd1 vssd1 vccd1 vccd1 _00986_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_66_2329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12944_ _07669_ net268 _07667_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[232\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_1179 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18451_ _04696_ _04791_ _03825_ _03939_ vssd1 vssd1 vccd1 vccd1 _03940_ sky130_fd_sc_hd__a31o_1
X_15663_ ag2.body\[411\] net143 _01625_ ag2.body\[403\] vssd1 vssd1 vccd1 vccd1 _00925_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_115_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12875_ net342 net316 vssd1 vssd1 vccd1 vccd1 _07638_ sky130_fd_sc_hd__nor2_4
X_17402_ ag2.body\[40\] net879 vssd1 vssd1 vccd1 vccd1 _03081_ sky130_fd_sc_hd__xor2_1
XFILLER_0_115_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14614_ net979 ag2.body\[58\] vssd1 vssd1 vccd1 vccd1 _08775_ sky130_fd_sc_hd__xnor2_1
XANTENNA__12426__A_N _06505_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18382_ _03786_ _03798_ vssd1 vssd1 vccd1 vccd1 _03872_ sky130_fd_sc_hd__nor2_1
X_11826_ img_gen.tracker.frame\[425\] net600 net584 img_gen.tracker.frame\[431\] _06797_
+ vssd1 vssd1 vccd1 vccd1 _06798_ sky130_fd_sc_hd__o221a_1
X_15594_ ag2.body\[477\] net122 _01618_ ag2.body\[469\] vssd1 vssd1 vccd1 vccd1 _00863_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_5_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_1492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_1574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17333_ ag2.body\[7\] net690 vssd1 vssd1 vccd1 vccd1 _03012_ sky130_fd_sc_hd__nor2_1
X_14545_ net983 ag2.body\[242\] vssd1 vssd1 vccd1 vccd1 _08706_ sky130_fd_sc_hd__xor2_1
XFILLER_0_56_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17202__B net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_134_clk clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_134_clk
+ sky130_fd_sc_hd__clkbuf_8
X_11757_ img_gen.tracker.frame\[254\] net615 net543 img_gen.tracker.frame\[260\] _06728_
+ vssd1 vssd1 vccd1 vccd1 _06729_ sky130_fd_sc_hd__o221a_1
XFILLER_0_56_779 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11531__A net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10708_ ag2.body\[19\] net1152 vssd1 vssd1 vccd1 vccd1 _05681_ sky130_fd_sc_hd__xor2_1
X_17264_ _04079_ net885 net873 _04080_ _02942_ vssd1 vssd1 vccd1 vccd1 _02943_ sky130_fd_sc_hd__a221o_1
X_14476_ net1036 ag2.body\[444\] vssd1 vssd1 vccd1 vccd1 _08637_ sky130_fd_sc_hd__xor2_1
XFILLER_0_86_1528 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11688_ _06630_ _06659_ _06658_ vssd1 vssd1 vccd1 vccd1 _06660_ sky130_fd_sc_hd__a21o_2
X_19003_ clknet_leaf_2_clk img_gen.tracker.next_frame\[441\] net1249 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[441\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__12346__B _06638_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16215_ net355 _01893_ vssd1 vssd1 vccd1 vccd1 _01894_ sky130_fd_sc_hd__nor2_1
Xclkload105 clknet_leaf_55_clk vssd1 vssd1 vccd1 vccd1 clkload105/Y sky130_fd_sc_hd__inv_6
X_13427_ net2102 net647 _07882_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[502\]
+ sky130_fd_sc_hd__and3_1
Xclkload116 clknet_leaf_63_clk vssd1 vssd1 vccd1 vccd1 clkload116/Y sky130_fd_sc_hd__clkinv_8
X_17195_ ag2.body\[179\] net852 vssd1 vssd1 vccd1 vccd1 _02874_ sky130_fd_sc_hd__xor2_1
X_10639_ net1218 control.body\[664\] vssd1 vssd1 vccd1 vccd1 _05612_ sky130_fd_sc_hd__xor2_1
Xclkload127 clknet_leaf_68_clk vssd1 vssd1 vccd1 vccd1 clkload127/Y sky130_fd_sc_hd__clkinv_2
XANTENNA__15570__A2 net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10147__A _04640_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16146_ obsg2.obstacleArray\[16\] net427 net374 _01824_ vssd1 vssd1 vccd1 vccd1 _01825_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_122_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13358_ net664 _07856_ vssd1 vssd1 vccd1 vccd1 _07857_ sky130_fd_sc_hd__nor2_1
XANTENNA__18033__B net38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12309_ _07210_ _07263_ _07264_ vssd1 vssd1 vccd1 vccd1 _07276_ sky130_fd_sc_hd__and3_1
XFILLER_0_122_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16077_ obsg2.obstacleArray\[108\] obsg2.obstacleArray\[109\] net421 vssd1 vssd1
+ vccd1 vccd1 _01756_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_127_4204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13289_ net671 _07829_ vssd1 vssd1 vccd1 vccd1 _07830_ sky130_fd_sc_hd__nor2_1
XFILLER_0_126_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_1410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_1421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12136__A2 net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19905_ clknet_leaf_86_clk _00849_ net1464 vssd1 vssd1 vccd1 vccd1 ag2.body\[495\]
+ sky130_fd_sc_hd__dfrtp_4
X_15028_ control.body\[982\] net166 _01555_ net2204 vssd1 vssd1 vccd1 vccd1 _00360_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_36_1432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13177__B net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_18_Right_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18549__CLK clknet_leaf_131_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18272__A1 net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19836_ clknet_leaf_92_clk _00780_ net1414 vssd1 vssd1 vccd1 vccd1 ag2.body\[554\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_97_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19767_ clknet_leaf_19_clk _00711_ net1321 vssd1 vssd1 vccd1 vccd1 control.body\[629\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput3 gpio_in[26] vssd1 vssd1 vccd1 vccd1 net3 sky130_fd_sc_hd__clkbuf_1
X_16979_ ag2.body\[431\] net931 vssd1 vssd1 vccd1 vccd1 _02658_ sky130_fd_sc_hd__xnor2_1
XANTENNA__14289__A net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09520_ net909 net905 vssd1 vssd1 vccd1 vccd1 _04493_ sky130_fd_sc_hd__or2_4
X_18718_ clknet_leaf_142_clk img_gen.tracker.next_frame\[156\] net1258 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[156\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_49_1804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_1212 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10610__A net1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19698_ clknet_leaf_136_clk _00642_ net1300 vssd1 vssd1 vccd1 vccd1 control.body\[688\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_49_1826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09451_ net919 net915 net922 vssd1 vssd1 vccd1 vccd1 _04424_ sky130_fd_sc_hd__and3_1
X_18649_ clknet_leaf_130_clk img_gen.tracker.next_frame\[87\] net1317 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[87\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_56_1387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09382_ _04365_ _04375_ vssd1 vssd1 vccd1 vccd1 _01412_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_27_Right_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15722__A_N _04719_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_3340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_595 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20611_ net1543 vssd1 vssd1 vccd1 vccd1 gpio_oeb[23] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_99_3351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_125_clk clknet_4_9__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_125_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__17112__B net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12537__A net225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17535__B1 net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_3215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11441__A net1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout238_A net247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_3226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16889__A2 net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20542_ clknet_leaf_105_clk _01407_ _00016_ vssd1 vssd1 vccd1 vccd1 sound_gen.osc1.stayCount\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_62_727 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16951__B net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11160__B net1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20473_ clknet_leaf_31_clk _01360_ net1338 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[109\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_85_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14752__A net975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16443__S net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout405_A net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1147_A net1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15200__X _01574_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09846__A net1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19324__CLK clknet_leaf_103_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09776__B1 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13368__A net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09565__B _04445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16510__A1 obsg2.obstacleArray\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1314_A net1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_36_Right_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1009 net1014 vssd1 vssd1 vccd1 vccd1 net1009 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_7_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout774_A _04229_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout395_X net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1102_X net1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout941_A obsg2.randCord\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14199__A net1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout562_X net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14824__A1 net1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14824__B2 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11638__A1 _06511_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09718_ net770 ag2.body\[243\] _04075_ net1231 vssd1 vssd1 vccd1 vccd1 _04691_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_97_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10990_ _05937_ _05938_ _05947_ _05949_ net478 vssd1 vssd1 vccd1 vccd1 _05963_ sky130_fd_sc_hd__a41o_1
XANTENNA_fanout53_A net54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09649_ net1073 control.body\[750\] vssd1 vssd1 vccd1 vccd1 _04622_ sky130_fd_sc_hd__or2_1
XANTENNA__16577__A1 net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout827_X net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_45_Right_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_1498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12660_ net288 _07533_ _07534_ net2044 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[83\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_96_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11611_ _06578_ _06583_ _06497_ vssd1 vssd1 vccd1 vccd1 _06584_ sky130_fd_sc_hd__or3b_1
XFILLER_0_33_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16329__A1 net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12063__A1 net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17526__B1 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12591_ net250 net308 _07495_ _07496_ net1623 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[52\]
+ sky130_fd_sc_hd__a32o_1
Xclkbuf_leaf_116_clk clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_116_clk
+ sky130_fd_sc_hd__clkbuf_8
X_14330_ net827 ag2.body\[426\] _04153_ net1017 vssd1 vssd1 vccd1 vccd1 _08491_ sky130_fd_sc_hd__a22o_1
XFILLER_0_107_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11542_ obsg2.obstacleArray\[104\] obsg2.obstacleArray\[105\] obsg2.obstacleArray\[108\]
+ obsg2.obstacleArray\[109\] net1125 net511 vssd1 vssd1 vccd1 vccd1 _06515_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_78_2701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_2712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_59_2111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_2122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14261_ _08418_ _08419_ _08420_ _08421_ vssd1 vssd1 vccd1 vccd1 _08422_ sky130_fd_sc_hd__or4_1
XANTENNA__15758__A _05212_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11473_ _06442_ _06443_ _06444_ _06445_ vssd1 vssd1 vccd1 vccd1 _06446_ sky130_fd_sc_hd__or4_1
XANTENNA__15552__A2 net191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_2133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14662__A net1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16000_ net871 net939 vssd1 vssd1 vccd1 vccd1 _01679_ sky130_fd_sc_hd__and2_1
XANTENNA__18129__A_N _01691_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13212_ net289 _07794_ _07795_ net1852 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[374\]
+ sky130_fd_sc_hd__a22o_1
Xwire478 _05962_ vssd1 vssd1 vccd1 vccd1 net478 sky130_fd_sc_hd__buf_1
XANTENNA__09767__B1 _04688_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10424_ net769 control.body\[1067\] control.body\[1070\] net750 vssd1 vssd1 vccd1
+ vccd1 _05397_ sky130_fd_sc_hd__a22oi_1
XTAP_TAPCELL_ROW_55_2008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14192_ net1028 ag2.body\[165\] vssd1 vssd1 vccd1 vccd1 _08353_ sky130_fd_sc_hd__xor2_1
XFILLER_0_81_1425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_54_Right_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17973__A net45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13143_ net252 _07762_ _07763_ net1987 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[337\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__19817__CLK clknet_leaf_124_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13278__A net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16501__A1 net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09475__B net1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10355_ ag2.body\[290\] net1187 vssd1 vssd1 vccd1 vccd1 _05328_ sky130_fd_sc_hd__and2b_1
XANTENNA__12182__A net1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12613__C net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10286_ ag2.body\[335\] net1067 vssd1 vssd1 vccd1 vccd1 _05259_ sky130_fd_sc_hd__or2_1
X_17951_ net529 _03578_ vssd1 vssd1 vccd1 vccd1 _01259_ sky130_fd_sc_hd__and2_1
X_13074_ net266 _07729_ _07730_ net1901 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[301\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_57_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1510 net1511 vssd1 vssd1 vccd1 vccd1 net1510 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_20_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16902_ ag2.body\[246\] net943 vssd1 vssd1 vccd1 vccd1 _02581_ sky130_fd_sc_hd__nand2_1
X_12025_ img_gen.tracker.frame\[207\] net612 net557 img_gen.tracker.frame\[210\] _06996_
+ vssd1 vssd1 vccd1 vccd1 _06997_ sky130_fd_sc_hd__a221o_1
X_17882_ _04431_ _04758_ vssd1 vssd1 vccd1 vccd1 _03522_ sky130_fd_sc_hd__nand2_1
XANTENNA__12910__A _07315_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18841__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19621_ clknet_leaf_123_clk _00565_ net1407 vssd1 vssd1 vccd1 vccd1 control.body\[771\]
+ sky130_fd_sc_hd__dfrtp_1
X_16833_ ag2.body\[98\] net864 vssd1 vssd1 vccd1 vccd1 _02512_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_73_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16764_ obsg2.obstacleArray\[3\] net502 net484 obsg2.obstacleArray\[1\] _02442_ vssd1
+ vssd1 vccd1 vccd1 _02443_ sky130_fd_sc_hd__a221o_1
X_19552_ clknet_leaf_116_clk _00496_ net1387 vssd1 vssd1 vccd1 vccd1 control.body\[846\]
+ sky130_fd_sc_hd__dfrtp_1
X_13976_ ag2.body\[114\] net189 _08158_ ag2.body\[106\] vssd1 vssd1 vccd1 vccd1 _00195_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__10430__A net1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_63_Right_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_1543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15715_ ag2.body\[362\] net193 _01630_ ag2.body\[354\] vssd1 vssd1 vccd1 vccd1 _00972_
+ sky130_fd_sc_hd__a22o_1
X_18503_ net1515 net1509 vssd1 vssd1 vccd1 vccd1 _00034_ sky130_fd_sc_hd__or2_1
XANTENNA__11245__B net1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1636 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12927_ _07661_ net265 _07659_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[223\]
+ sky130_fd_sc_hd__mux2_1
X_16695_ obsg2.obstacleArray\[67\] net502 net488 obsg2.obstacleArray\[66\] vssd1 vssd1
+ vccd1 vccd1 _02374_ sky130_fd_sc_hd__a22o_1
X_19483_ clknet_leaf_114_clk _00427_ net1398 vssd1 vssd1 vccd1 vccd1 control.body\[905\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__17765__B1 _03218_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15646_ ag2.body\[428\] net138 _01623_ ag2.body\[420\] vssd1 vssd1 vccd1 vccd1 _00910_
+ sky130_fd_sc_hd__a22o_1
X_18434_ _03921_ _03922_ _03808_ _03918_ vssd1 vssd1 vccd1 vccd1 _03923_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_17_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12858_ net435 net467 _06672_ _07452_ vssd1 vssd1 vccd1 vccd1 _07630_ sky130_fd_sc_hd__or4_2
XFILLER_0_69_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18028__B _01713_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11532__Y _06505_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18365_ net464 track.nextHighScore\[6\] _03785_ _03796_ vssd1 vssd1 vccd1 vccd1 _03859_
+ sky130_fd_sc_hd__or4b_1
X_11809_ net558 _06777_ _06780_ vssd1 vssd1 vccd1 vccd1 _06781_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_127_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15577_ ag2.body\[495\] net135 _01615_ ag2.body\[487\] vssd1 vssd1 vccd1 vccd1 _00849_
+ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_107_clk clknet_4_10__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_107_clk
+ sky130_fd_sc_hd__clkbuf_8
X_12789_ net286 _07596_ _07597_ net2028 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[149\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_113_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17316_ ag2.body\[222\] net943 vssd1 vssd1 vccd1 vccd1 _02995_ sky130_fd_sc_hd__xor2_1
XFILLER_0_44_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11801__A1 net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14528_ net1010 ag2.body\[255\] vssd1 vssd1 vccd1 vccd1 _08689_ sky130_fd_sc_hd__nand2_1
X_18296_ track.nextHighScore\[6\] track.nextHighScore\[7\] vssd1 vssd1 vccd1 vccd1
+ _03792_ sky130_fd_sc_hd__nor2_2
XFILLER_0_56_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15668__A _04472_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17247_ ag2.body\[618\] net722 net937 _04225_ _02925_ vssd1 vssd1 vccd1 vccd1 _02926_
+ sky130_fd_sc_hd__o221a_1
X_14459_ _08618_ _08619_ vssd1 vssd1 vccd1 vccd1 _08620_ sky130_fd_sc_hd__nand2_1
XFILLER_0_71_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18044__A net42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_72_Right_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__20324__CLK clknet_leaf_43_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09666__A _04425_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17178_ ag2.body\[459\] net850 vssd1 vssd1 vccd1 vccd1 _02857_ sky130_fd_sc_hd__xor2_1
XFILLER_0_3_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11565__B1 net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19497__CLK clknet_leaf_113_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16129_ obsg2.obstacleArray\[75\] net430 net376 _01807_ vssd1 vssd1 vccd1 vccd1 _01808_
+ sky130_fd_sc_hd__o211a_1
XANTENNA__19962__RESET_B net1470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10605__A net1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13306__A1 net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08951_ ag2.body\[10\] vssd1 vssd1 vccd1 vccd1 _03976_ sky130_fd_sc_hd__inv_2
XFILLER_0_45_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10324__B net1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17048__A2 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_1543 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19819_ clknet_leaf_124_clk _00763_ net1411 vssd1 vssd1 vccd1 vccd1 ag2.body\[569\]
+ sky130_fd_sc_hd__dfrtp_4
XPHY_EDGE_ROW_16_Left_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_81_Right_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout188_A net192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09503_ ag2.body\[400\] net785 net752 ag2.body\[406\] vssd1 vssd1 vccd1 vccd1 _04476_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__16946__B net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11155__B net1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16438__S net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14747__A net1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1097_A net1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09434_ net1044 net1224 vssd1 vssd1 vccd1 vccd1 _04407_ sky130_fd_sc_hd__xor2_1
XANTENNA__17220__A2 net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10843__A2 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10994__B net1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09365_ sound_gen.osc1.stayCount\[17\] sound_gen.osc1.stayCount\[16\] sound_gen.osc1.stayCount\[15\]
+ _04366_ vssd1 vssd1 vccd1 vccd1 _04367_ sky130_fd_sc_hd__and4_1
XFILLER_0_118_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout522_A net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11171__A net1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_30 _03442_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09296_ _04311_ _04313_ _04315_ sound_gen.osc1.count\[5\] vssd1 vssd1 vccd1 vccd1
+ _04316_ sky130_fd_sc_hd__a211o_1
XFILLER_0_7_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_25_Left_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_1545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_90_Right_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15578__A _04429_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18714__CLK clknet_leaf_144_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20525_ clknet_leaf_112_clk track.nextCurrScore\[7\] net1426 vssd1 vssd1 vccd1 vccd1
+ control.body_update.curr_length\[7\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__16173__S net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12554__X _07476_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout408_X net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1052_X net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20456_ clknet_leaf_38_clk _01343_ net1355 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[92\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_120_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout891_A net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout989_A net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17287__A2 net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20387_ clknet_leaf_40_clk _01274_ net1374 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[23\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_101_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10140_ net637 _05110_ _05111_ _05112_ vssd1 vssd1 vccd1 vccd1 _05113_ sky130_fd_sc_hd__or4_1
XANTENNA__10234__B net1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout777_X net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17039__A2 net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10071_ net1193 control.body\[713\] vssd1 vssd1 vccd1 vccd1 _05044_ sky130_fd_sc_hd__or2_1
XANTENNA__11859__A1 net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_34_Left_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09921__B1 net1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17017__B net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout944_X net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13830_ _08111_ _08112_ _08117_ _08120_ _08123_ vssd1 vssd1 vccd1 vccd1 _08127_ sky130_fd_sc_hd__a41o_1
XANTENNA_fanout56_X net56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16856__B net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_966 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13761_ img_gen.updater.commands.count\[5\] _08075_ vssd1 vssd1 vccd1 vccd1 _08077_
+ sky130_fd_sc_hd__and2_1
XANTENNA__16348__S net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10973_ net1179 control.body\[1002\] vssd1 vssd1 vccd1 vccd1 _05946_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_134_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15500_ ag2.body\[554\] net113 _01607_ ag2.body\[546\] vssd1 vssd1 vccd1 vccd1 _00780_
+ sky130_fd_sc_hd__a22o_1
X_12712_ net260 _07559_ _07560_ net1887 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[109\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_116_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16480_ obsg2.obstacleArray\[39\] _02059_ net397 _02158_ vssd1 vssd1 vccd1 vccd1
+ _02159_ sky130_fd_sc_hd__o211a_1
X_13692_ net639 _04427_ _04554_ vssd1 vssd1 vccd1 vccd1 _08034_ sky130_fd_sc_hd__and3_1
X_15431_ ag2.body\[621\] net84 _01599_ ag2.body\[613\] vssd1 vssd1 vccd1 vccd1 _00719_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__17968__A net43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12643_ net242 _07524_ _07525_ net2138 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[75\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_127_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_1447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10249__X _05222_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_43_Left_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_811 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18150_ net47 _03577_ _03704_ obsg2.obstacleArray\[72\] vssd1 vssd1 vccd1 vccd1 _03714_
+ sky130_fd_sc_hd__a31o_1
XANTENNA__12608__C _07505_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15362_ control.body\[687\] net68 _01592_ net2496 vssd1 vssd1 vccd1 vccd1 _00657_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__17687__B net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12574_ net330 _07486_ vssd1 vssd1 vccd1 vccd1 _07487_ sky130_fd_sc_hd__nor2_1
XFILLER_0_93_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17101_ ag2.body\[8\] net882 vssd1 vssd1 vccd1 vccd1 _02780_ sky130_fd_sc_hd__nand2_1
XFILLER_0_68_1022 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14313_ net996 ag2.body\[48\] vssd1 vssd1 vccd1 vccd1 _08474_ sky130_fd_sc_hd__xor2_1
XFILLER_0_4_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11525_ obsg2.obstacleArray\[120\] obsg2.obstacleArray\[121\] obsg2.obstacleArray\[124\]
+ obsg2.obstacleArray\[125\] net1125 net511 vssd1 vssd1 vccd1 vccd1 _06498_ sky130_fd_sc_hd__mux4_1
XFILLER_0_110_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18081_ _01714_ _03540_ net300 vssd1 vssd1 vccd1 vccd1 _03670_ sky130_fd_sc_hd__and3_1
XFILLER_0_81_866 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16183__C1 _01742_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15293_ control.body\[737\] net77 _01585_ net2240 vssd1 vssd1 vccd1 vccd1 _00595_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_41_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_1629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17032_ _04146_ net945 net693 ag2.body\[407\] _02710_ vssd1 vssd1 vccd1 vccd1 _02711_
+ sky130_fd_sc_hd__a221o_1
X_14244_ net1011 ag2.body\[543\] vssd1 vssd1 vccd1 vccd1 _08405_ sky130_fd_sc_hd__xor2_1
XFILLER_0_68_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11456_ ag2.body\[263\] net1066 vssd1 vssd1 vccd1 vccd1 _06429_ sky130_fd_sc_hd__or2_1
XFILLER_0_40_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20497__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_1218 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10407_ net1205 control.body\[1073\] vssd1 vssd1 vccd1 vccd1 _05380_ sky130_fd_sc_hd__xor2_1
XFILLER_0_46_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14175_ net1007 ag2.body\[199\] vssd1 vssd1 vccd1 vccd1 _08336_ sky130_fd_sc_hd__or2_1
XFILLER_0_46_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11387_ net1073 control.body\[646\] vssd1 vssd1 vccd1 vccd1 _06360_ sky130_fd_sc_hd__or2_1
XFILLER_0_110_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13126_ net291 _07752_ _07753_ net1697 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[329\]
+ sky130_fd_sc_hd__a22o_1
X_10338_ ag2.body\[526\] net1085 vssd1 vssd1 vccd1 vccd1 _05311_ sky130_fd_sc_hd__or2_1
XFILLER_0_81_1299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18983_ clknet_leaf_8_clk img_gen.tracker.next_frame\[421\] net1270 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[421\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_123_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_52_Left_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17934_ obsg2.obstacleArray\[4\] _03565_ net534 vssd1 vssd1 vccd1 vccd1 _01255_ sky130_fd_sc_hd__o21a_1
XANTENNA__09933__B net1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13057_ _07722_ net268 _07720_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[292\]
+ sky130_fd_sc_hd__mux2_1
X_10269_ ag2.body\[140\] net1141 vssd1 vssd1 vccd1 vccd1 _05242_ sky130_fd_sc_hd__xor2_1
XFILLER_0_84_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12640__A _06671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10712__X _05685_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1340 net1341 vssd1 vssd1 vccd1 vccd1 net1340 sky130_fd_sc_hd__clkbuf_4
X_12008_ img_gen.tracker.frame\[460\] net597 net578 img_gen.tracker.frame\[466\] vssd1
+ vssd1 vccd1 vccd1 _06980_ sky130_fd_sc_hd__o22a_1
Xfanout1351 net1357 vssd1 vssd1 vccd1 vccd1 net1351 sky130_fd_sc_hd__clkbuf_4
XANTENNA__16789__A1 _01700_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17865_ net2139 _03501_ vssd1 vssd1 vccd1 vccd1 _01238_ sky130_fd_sc_hd__xor2_1
Xfanout1362 net1370 vssd1 vssd1 vccd1 vccd1 net1362 sky130_fd_sc_hd__buf_2
Xfanout1373 net1374 vssd1 vssd1 vccd1 vccd1 net1373 sky130_fd_sc_hd__buf_2
XFILLER_0_89_900 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1384 net1385 vssd1 vssd1 vccd1 vccd1 net1384 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10522__B2 _05494_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19604_ clknet_leaf_119_clk _00548_ net1390 vssd1 vssd1 vccd1 vccd1 control.body\[786\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11256__A net1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16816_ ag2.body\[83\] net855 vssd1 vssd1 vccd1 vccd1 _02495_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_75_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1395 net1404 vssd1 vssd1 vccd1 vccd1 net1395 sky130_fd_sc_hd__buf_2
XFILLER_0_108_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17796_ net969 net958 vssd1 vssd1 vccd1 vccd1 _01215_ sky130_fd_sc_hd__xor2_1
XANTENNA__17591__A1_N ag2.body\[59\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19535_ clknet_leaf_118_clk _00479_ net1393 vssd1 vssd1 vccd1 vccd1 control.body\[861\]
+ sky130_fd_sc_hd__dfrtp_1
X_16747_ obsg2.obstacleArray\[56\] net491 net482 obsg2.obstacleArray\[57\] vssd1 vssd1
+ vccd1 vccd1 _02426_ sky130_fd_sc_hd__a22o_1
X_13959_ ag2.body\[99\] net189 _08156_ ag2.body\[91\] vssd1 vssd1 vccd1 vccd1 _00180_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_92_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13471__A net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16678_ net357 _02296_ _02300_ _02308_ _02212_ vssd1 vssd1 vccd1 vccd1 _02357_ sky130_fd_sc_hd__a311o_1
X_19466_ clknet_leaf_110_clk _00410_ net1418 vssd1 vssd1 vccd1 vccd1 control.body\[920\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10825__A2 _04758_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18417_ _03821_ _03905_ _03906_ vssd1 vssd1 vccd1 vccd1 _03907_ sky130_fd_sc_hd__or3_1
XANTENNA__12027__A1 net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15629_ ag2.body\[445\] net125 _01621_ ag2.body\[437\] vssd1 vssd1 vccd1 vccd1 _00895_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__18737__CLK clknet_leaf_142_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15764__A2 net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19397_ clknet_leaf_111_clk _00341_ net1425 vssd1 vssd1 vccd1 vccd1 control.body\[995\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09150_ ag2.body\[483\] vssd1 vssd1 vccd1 vccd1 _04175_ sky130_fd_sc_hd__inv_2
XFILLER_0_72_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18348_ _03820_ _03843_ _08036_ vssd1 vssd1 vccd1 vccd1 _03844_ sky130_fd_sc_hd__a21oi_2
XANTENNA__14972__B1 net51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11786__B1 net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10319__B net1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16174__C1 _01742_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09081_ ag2.body\[316\] vssd1 vssd1 vccd1 vccd1 _04106_ sky130_fd_sc_hd__inv_2
X_18279_ net530 _03778_ vssd1 vssd1 vccd1 vccd1 _01387_ sky130_fd_sc_hd__and2_1
X_20310_ clknet_leaf_44_clk _01210_ net1380 vssd1 vssd1 vccd1 vccd1 ag2.randCord\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_wire480_X net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold801 control.body\[833\] vssd1 vssd1 vccd1 vccd1 net2363 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__16006__B net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold812 control.body\[1106\] vssd1 vssd1 vccd1 vccd1 net2374 sky130_fd_sc_hd__dlygate4sd3_1
X_20241_ clknet_leaf_69_clk _01185_ net1496 vssd1 vssd1 vccd1 vccd1 ag2.body\[159\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_9_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold823 _00350_ vssd1 vssd1 vccd1 vccd1 net2385 sky130_fd_sc_hd__dlygate4sd3_1
Xhold834 control.body\[668\] vssd1 vssd1 vccd1 vccd1 net2396 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__17269__A2 net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold845 _00282_ vssd1 vssd1 vccd1 vccd1 net2407 sky130_fd_sc_hd__dlygate4sd3_1
Xhold856 control.body\[723\] vssd1 vssd1 vccd1 vccd1 net2418 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold867 control.body\[874\] vssd1 vssd1 vccd1 vccd1 net2429 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20172_ clknet_leaf_83_clk _01116_ net1480 vssd1 vssd1 vccd1 vccd1 ag2.body\[218\]
+ sky130_fd_sc_hd__dfrtp_4
Xhold878 control.body\[795\] vssd1 vssd1 vccd1 vccd1 net2440 sky130_fd_sc_hd__dlygate4sd3_1
Xhold889 control.body\[992\] vssd1 vssd1 vccd1 vccd1 net2451 sky130_fd_sc_hd__dlygate4sd3_1
X_09983_ net1111 control.body\[1117\] vssd1 vssd1 vccd1 vccd1 _04956_ sky130_fd_sc_hd__or2_1
XANTENNA__10054__B net1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10761__A1 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10761__B2 net1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08934_ sound_gen.osc1.stayCount\[21\] vssd1 vssd1 vccd1 vccd1 _03959_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout1012_A net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09903__B1 _04858_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout472_A _06647_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_1224 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11710__B1 net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11166__A net1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10070__A net1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17729__B1 net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout260_X net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout737_A _04262_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14477__A net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11453__X _06426_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1479_A net1480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_0_Right_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12709__B _07558_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09417_ net969 net663 vssd1 vssd1 vccd1 vccd1 _04396_ sky130_fd_sc_hd__nand2_1
XFILLER_0_82_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10029__B1 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09348_ sound_gen.osc1.stayCount\[22\] _04351_ vssd1 vssd1 vccd1 vccd1 _04352_ sky130_fd_sc_hd__nand2_1
XFILLER_0_35_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14963__B1 _01547_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10229__B net1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16165__C1 net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09279_ sound_gen.osc1.stayCount\[23\] _04287_ sound_gen.osc1.stayCount\[22\] vssd1
+ vssd1 vccd1 vccd1 _04302_ sky130_fd_sc_hd__a21o_1
XFILLER_0_106_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13518__A1 net226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11310_ ag2.body\[278\] net1086 vssd1 vssd1 vccd1 vccd1 _06283_ sky130_fd_sc_hd__xor2_1
XFILLER_0_65_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20508_ clknet_leaf_112_clk net2301 net1424 vssd1 vssd1 vccd1 vccd1 score_detect.N\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_12290_ _07258_ _07259_ vssd1 vssd1 vccd1 vccd1 img_gen.updater.update.next\[0\]
+ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout894_X net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11241_ ag2.body\[198\] net1080 vssd1 vssd1 vccd1 vccd1 _06214_ sky130_fd_sc_hd__or2_1
XANTENNA__11624__S0 net1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20439_ clknet_leaf_26_clk _01326_ net1343 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[75\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_47_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_1586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_459 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11172_ net1099 control.body\[781\] vssd1 vssd1 vccd1 vccd1 _06145_ sky130_fd_sc_hd__xor2_1
XANTENNA__11661__A_N _06612_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19042__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10123_ net1072 control.body\[710\] vssd1 vssd1 vccd1 vccd1 _05096_ sky130_fd_sc_hd__nand2_1
X_15980_ _03964_ _01663_ _01664_ vssd1 vssd1 vccd1 vccd1 _01665_ sky130_fd_sc_hd__or3_1
XANTENNA__17680__A2 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09753__B net1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10054_ ag2.body\[484\] net1138 vssd1 vssd1 vccd1 vccd1 _05027_ sky130_fd_sc_hd__nand2_1
X_14931_ net2195 net173 _01544_ net2285 vssd1 vssd1 vccd1 vccd1 _00274_ sky130_fd_sc_hd__a22o_1
XFILLER_0_76_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17315__X _02994_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17432__A2 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14862_ _01526_ _01527_ _01528_ _01532_ vssd1 vssd1 vccd1 vccd1 _01533_ sky130_fd_sc_hd__and4_1
X_17650_ ag2.body\[38\] net937 vssd1 vssd1 vccd1 vccd1 _03329_ sky130_fd_sc_hd__xor2_1
XANTENNA__19192__CLK clknet_leaf_53_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13813_ control.body_update.direction\[2\] control.body_update.direction\[1\] vssd1
+ vssd1 vccd1 vccd1 _08110_ sky130_fd_sc_hd__or2_1
X_16601_ obsg2.obstacleArray\[85\] net451 _02216_ vssd1 vssd1 vccd1 vccd1 _02280_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_118_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17581_ _04118_ net888 net720 ag2.body\[339\] vssd1 vssd1 vccd1 vccd1 _03260_ sky130_fd_sc_hd__a22o_1
X_14793_ net794 ag2.body\[551\] ag2.body\[549\] net808 vssd1 vssd1 vccd1 vccd1 _01464_
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_138_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_121_Right_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16532_ _02206_ _02210_ vssd1 vssd1 vccd1 vccd1 _02211_ sky130_fd_sc_hd__nor2_4
XFILLER_0_98_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19320_ clknet_leaf_104_clk net2206 net1433 vssd1 vssd1 vccd1 vccd1 control.body\[1078\]
+ sky130_fd_sc_hd__dfrtp_1
X_13744_ _08064_ net320 img_gen.updater.commands.count\[0\] vssd1 vssd1 vccd1 vccd1
+ _00057_ sky130_fd_sc_hd__mux2_1
X_10956_ ag2.body\[172\] net1129 vssd1 vssd1 vccd1 vccd1 _05929_ sky130_fd_sc_hd__nand2_1
XFILLER_0_6_1420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_504 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12619__B net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16463_ net397 _02141_ vssd1 vssd1 vccd1 vccd1 _02142_ sky130_fd_sc_hd__or2_1
X_19251_ clknet_leaf_75_clk _00195_ net1482 vssd1 vssd1 vccd1 vccd1 ag2.body\[114\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__18009__D net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13675_ _04402_ _07181_ vssd1 vssd1 vccd1 vccd1 _08022_ sky130_fd_sc_hd__nor2_2
XFILLER_0_6_1475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10887_ net1118 control.body\[652\] vssd1 vssd1 vccd1 vccd1 _05860_ sky130_fd_sc_hd__xor2_1
X_18202_ _03645_ net40 vssd1 vssd1 vccd1 vccd1 _03740_ sky130_fd_sc_hd__nor2_1
XANTENNA__12338__C net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15414_ net2589 net81 _01597_ control.body\[630\] vssd1 vssd1 vccd1 vccd1 _00704_
+ sky130_fd_sc_hd__a22o_1
X_12626_ net593 _06639_ net440 net569 vssd1 vssd1 vccd1 vccd1 _07515_ sky130_fd_sc_hd__and4_2
X_19182_ clknet_leaf_20_clk _00126_ net1331 vssd1 vssd1 vccd1 vccd1 ag2.body\[45\]
+ sky130_fd_sc_hd__dfrtp_4
X_16394_ obsg2.obstacleArray\[124\] obsg2.obstacleArray\[125\] obsg2.obstacleArray\[126\]
+ obsg2.obstacleArray\[127\] net454 net398 vssd1 vssd1 vccd1 vccd1 _02073_ sky130_fd_sc_hd__mux4_1
XANTENNA__14954__B1 _01546_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11768__B1 net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18133_ _03549_ net296 vssd1 vssd1 vccd1 vccd1 _03704_ sky130_fd_sc_hd__nor2_2
XFILLER_0_87_1442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15345_ _05827_ net52 vssd1 vssd1 vccd1 vccd1 _01591_ sky130_fd_sc_hd__nor2_2
XANTENNA__16156__C1 net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12557_ net2079 net660 _07477_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[37\]
+ sky130_fd_sc_hd__and3_1
XANTENNA__17210__B net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12635__A net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_max_cap368_A _01911_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13509__A1 net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18025__C net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18064_ net42 _03658_ vssd1 vssd1 vccd1 vccd1 _03659_ sky130_fd_sc_hd__nor2_1
X_11508_ _06461_ _06463_ _06460_ vssd1 vssd1 vccd1 vccd1 _06481_ sky130_fd_sc_hd__a21o_1
XFILLER_0_124_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15276_ net2361 net88 _01583_ control.body\[746\] vssd1 vssd1 vccd1 vccd1 _00580_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_125_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12488_ net290 _07436_ _07437_ net1596 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[8\]
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_130_4277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold108 img_gen.tracker.frame\[218\] vssd1 vssd1 vccd1 vccd1 net1670 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_130_4288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17015_ ag2.body\[328\] net888 vssd1 vssd1 vccd1 vccd1 _02694_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_130_4299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14227_ _08385_ _08386_ _08387_ vssd1 vssd1 vccd1 vccd1 _08388_ sky130_fd_sc_hd__or3b_1
Xhold119 img_gen.tracker.frame\[491\] vssd1 vssd1 vccd1 vccd1 net1681 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__15946__A _04832_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11439_ _06404_ _06405_ _06406_ _06411_ vssd1 vssd1 vccd1 vccd1 _06412_ sky130_fd_sc_hd__or4_2
XFILLER_0_112_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_1615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_1172 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09944__A net1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14158_ net979 _04223_ _04225_ net1015 _08316_ vssd1 vssd1 vccd1 vccd1 _08319_ sky130_fd_sc_hd__a221o_1
XANTENNA__11940__B1 net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11685__S net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13466__A net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13109_ _07747_ net258 _07745_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[319\]
+ sky130_fd_sc_hd__mux2_1
XANTENNA__09663__B net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14089_ net1010 ag2.body\[287\] vssd1 vssd1 vccd1 vccd1 _08250_ sky130_fd_sc_hd__xor2_1
X_18966_ clknet_leaf_5_clk img_gen.tracker.next_frame\[404\] net1268 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[404\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__12370__A net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19535__CLK clknet_leaf_118_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12801__C _07505_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17917_ net355 _03535_ vssd1 vssd1 vccd1 vccd1 _03551_ sky130_fd_sc_hd__nor2_1
XANTENNA__13185__B net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18897_ clknet_leaf_12_clk img_gen.tracker.next_frame\[335\] net1285 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[335\] sky130_fd_sc_hd__dfrtp_1
Xfanout1170 net1172 vssd1 vssd1 vccd1 vccd1 net1170 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_52_1899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1181 net1183 vssd1 vssd1 vccd1 vccd1 net1181 sky130_fd_sc_hd__buf_4
X_17848_ img_gen.updater.commands.rR1.rainbowRNG\[10\] _03503_ vssd1 vssd1 vccd1 vccd1
+ _03504_ sky130_fd_sc_hd__and2_1
Xfanout1192 net1194 vssd1 vssd1 vccd1 vccd1 net1192 sky130_fd_sc_hd__clkbuf_4
XANTENNA__20512__CLK clknet_leaf_113_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16631__B1 net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17779_ _04260_ obsg2.obsNeeded\[2\] net530 _04398_ vssd1 vssd1 vccd1 vccd1 _03458_
+ sky130_fd_sc_hd__o211a_2
XANTENNA__14297__A net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_64 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19518_ clknet_leaf_121_clk _00462_ net1402 vssd1 vssd1 vccd1 vccd1 control.body\[876\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11433__B net1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15198__B1 _01573_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19449_ clknet_leaf_109_clk _00393_ net1420 vssd1 vssd1 vccd1 vccd1 control.body\[951\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_100_3380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09202_ net1230 vssd1 vssd1 vccd1 vccd1 _04227_ sky130_fd_sc_hd__inv_2
XFILLER_0_119_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11759__B1 net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18216__B net40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09133_ ag2.body\[444\] vssd1 vssd1 vccd1 vccd1 _04158_ sky130_fd_sc_hd__inv_2
XFILLER_0_115_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12420__A1 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16017__A net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout318_A _01818_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16698__B1 net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09064_ ag2.body\[263\] vssd1 vssd1 vccd1 vccd1 _04089_ sky130_fd_sc_hd__inv_2
XFILLER_0_4_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_113_3763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14173__A1 net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_3774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14173__B2 net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15370__B1 _01593_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15856__A _04740_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16451__S net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11606__S0 net1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10065__A net1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold620 control.body\[809\] vssd1 vssd1 vccd1 vccd1 net2182 sky130_fd_sc_hd__dlygate4sd3_1
Xhold631 img_gen.updater.commands.rR1.rainbowRNG\[3\] vssd1 vssd1 vccd1 vccd1 net2193
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold642 control.body\[974\] vssd1 vssd1 vccd1 vccd1 net2204 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1227_A net1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold653 control.body\[793\] vssd1 vssd1 vccd1 vccd1 net2215 sky130_fd_sc_hd__dlygate4sd3_1
X_20224_ clknet_leaf_60_clk _01168_ net1469 vssd1 vssd1 vccd1 vccd1 ag2.body\[174\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__09854__A net1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13920__B2 ag2.body\[56\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold664 control.body\[650\] vssd1 vssd1 vccd1 vccd1 net2226 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold675 control.body\[1013\] vssd1 vssd1 vccd1 vccd1 net2237 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11931__B1 _06661_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold686 control.body\[628\] vssd1 vssd1 vccd1 vccd1 net2248 sky130_fd_sc_hd__dlygate4sd3_1
Xhold697 control.body\[647\] vssd1 vssd1 vccd1 vccd1 net2259 sky130_fd_sc_hd__dlygate4sd3_1
X_20155_ clknet_leaf_94_clk _01099_ net1442 vssd1 vssd1 vccd1 vccd1 ag2.body\[233\]
+ sky130_fd_sc_hd__dfrtp_4
X_09966_ ag2.body\[82\] net1184 vssd1 vssd1 vccd1 vccd1 _04939_ sky130_fd_sc_hd__xor2_1
XFILLER_0_25_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1015_X net1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20086_ clknet_leaf_77_clk _01030_ net1491 vssd1 vssd1 vccd1 vccd1 ag2.body\[308\]
+ sky130_fd_sc_hd__dfrtp_4
X_09897_ _04865_ _04866_ _04868_ _04869_ vssd1 vssd1 vccd1 vccd1 _04870_ sky130_fd_sc_hd__a22o_1
XFILLER_0_99_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10512__B net1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout854_A net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_96_clk clknet_4_11__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_96_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__17414__A2 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20192__CLK clknet_leaf_88_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_1_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11695__C1 net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_3578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_3589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout642_X net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10810_ net1182 control.body\[1090\] vssd1 vssd1 vccd1 vccd1 _05783_ sky130_fd_sc_hd__nand2_1
X_11790_ img_gen.tracker.frame\[377\] net603 vssd1 vssd1 vccd1 vccd1 _06762_ sky130_fd_sc_hd__or2_1
XFILLER_0_138_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_1299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11343__B net1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10741_ ag2.body\[502\] net1089 vssd1 vssd1 vccd1 vccd1 _05714_ sky130_fd_sc_hd__or2_1
XANTENNA__11462__A2 net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_81_2785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout907_X net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17949__C net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_81_2796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13460_ _07587_ net302 vssd1 vssd1 vccd1 vccd1 _07896_ sky130_fd_sc_hd__nor2_1
X_10672_ ag2.body\[348\] net1141 vssd1 vssd1 vccd1 vccd1 _05645_ sky130_fd_sc_hd__xor2_1
X_12411_ _06472_ _06505_ _07354_ _07373_ _07299_ vssd1 vssd1 vccd1 vccd1 _07374_ sky130_fd_sc_hd__a32o_1
XANTENNA__19408__CLK clknet_leaf_103_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13391_ net275 _07868_ _07869_ net1926 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[479\]
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_11_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_20_clk clknet_4_6__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_20_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__16689__B1 _02211_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15130_ net2640 net103 _01566_ net2326 vssd1 vssd1 vccd1 vccd1 _00451_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_11_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12342_ net383 _07307_ vssd1 vssd1 vccd1 vccd1 _07309_ sky130_fd_sc_hd__xnor2_1
XANTENNA__17965__B _01713_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15061_ control.body\[947\] net150 _01559_ net2474 vssd1 vssd1 vccd1 vccd1 _00389_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__15361__B1 _01592_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12273_ img_gen.updater.commands.cmd_num\[4\] _07232_ _07241_ _07226_ vssd1 vssd1
+ vccd1 vccd1 _07243_ sky130_fd_sc_hd__a22o_1
XANTENNA__14670__A net1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15900__A2 net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14012_ net972 ag2.body\[459\] vssd1 vssd1 vccd1 vccd1 _08173_ sky130_fd_sc_hd__xnor2_1
XANTENNA__19558__CLK clknet_leaf_115_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13911__A1 ag2.body\[56\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09764__A ag2.body\[213\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11224_ net1227 control.body\[856\] vssd1 vssd1 vccd1 vccd1 _06197_ sky130_fd_sc_hd__xor2_1
XANTENNA__12902__B net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11358__X _06331_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15113__B1 _01554_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18820_ clknet_leaf_2_clk img_gen.tracker.next_frame\[258\] net1248 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[258\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__10262__X _05235_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11155_ ag2.body\[607\] net1048 vssd1 vssd1 vccd1 vccd1 _06128_ sky130_fd_sc_hd__or2_1
XANTENNA__12190__A net1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_1557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_1419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16861__B1 net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10106_ net1058 control.body\[943\] vssd1 vssd1 vccd1 vccd1 _05079_ sky130_fd_sc_hd__or2_1
X_18751_ clknet_leaf_143_clk img_gen.tracker.next_frame\[189\] net1255 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[189\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__11518__B net1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15963_ ag2.body\[151\] net199 _01657_ ag2.body\[143\] vssd1 vssd1 vccd1 vccd1 _01193_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_95_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11086_ ag2.body\[536\] net783 net746 ag2.body\[543\] _06058_ vssd1 vssd1 vccd1 vccd1
+ _06059_ sky130_fd_sc_hd__a221o_1
XFILLER_0_65_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_87_clk clknet_4_12__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_87_clk
+ sky130_fd_sc_hd__clkbuf_8
X_17702_ obsg2.obstacleArray\[136\] obsg2.obstacleArray\[137\] net410 vssd1 vssd1
+ vccd1 vccd1 _03381_ sky130_fd_sc_hd__mux2_1
X_14914_ control.body\[1073\] net170 _01542_ net2293 vssd1 vssd1 vccd1 vccd1 _00259_
+ sky130_fd_sc_hd__a22o_1
X_10037_ ag2.body\[507\] net771 _04416_ _04944_ _05007_ vssd1 vssd1 vccd1 vccd1 _05010_
+ sky130_fd_sc_hd__a221o_1
XANTENNA__17405__A2 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18682_ clknet_leaf_28_clk img_gen.tracker.next_frame\[120\] net1336 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[120\] sky130_fd_sc_hd__dfrtp_1
X_15894_ ag2.body\[201\] net133 _01650_ ag2.body\[193\] vssd1 vssd1 vccd1 vccd1 _01131_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_123_4070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16613__B1 net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17633_ ag2.body\[164\] net961 vssd1 vssd1 vccd1 vccd1 _03312_ sky130_fd_sc_hd__or2_1
X_14845_ _08660_ _08663_ _08552_ vssd1 vssd1 vccd1 vccd1 _01516_ sky130_fd_sc_hd__o21a_1
XFILLER_0_81_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17564_ ag2.body\[581\] net950 vssd1 vssd1 vccd1 vccd1 _03243_ sky130_fd_sc_hd__or2_1
X_14776_ net1030 ag2.body\[277\] vssd1 vssd1 vccd1 vccd1 _01447_ sky130_fd_sc_hd__xor2_1
XFILLER_0_98_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11988_ img_gen.tracker.frame\[403\] net545 vssd1 vssd1 vccd1 vccd1 _06960_ sky130_fd_sc_hd__or2_1
XANTENNA__12349__B _07315_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11989__B1 net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19303_ clknet_leaf_100_clk _00247_ net1443 vssd1 vssd1 vccd1 vccd1 control.body\[1093\]
+ sky130_fd_sc_hd__dfrtp_1
X_16515_ net365 _02193_ _02192_ net363 vssd1 vssd1 vccd1 vccd1 _02194_ sky130_fd_sc_hd__o211a_1
X_13727_ net2078 toggle1.nextBlinkToggle\[0\] toggle1.nextBlinkToggle\[1\] net1951
+ vssd1 vssd1 vccd1 vccd1 toggle1.nextDisplayOut\[3\] sky130_fd_sc_hd__a22o_1
XFILLER_0_54_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10939_ ag2.body\[301\] net1115 vssd1 vssd1 vccd1 vccd1 _05912_ sky130_fd_sc_hd__xor2_1
X_17495_ _03170_ _03171_ _03173_ vssd1 vssd1 vccd1 vccd1 _03174_ sky130_fd_sc_hd__and3b_1
XFILLER_0_15_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_4464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19234_ clknet_leaf_84_clk _00178_ net1481 vssd1 vssd1 vccd1 vccd1 ag2.body\[97\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__14927__B1 _01543_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09498__X _04471_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13658_ net2170 _08011_ net221 vssd1 vssd1 vccd1 vccd1 control.divider.next_count\[20\]
+ sky130_fd_sc_hd__o21a_1
X_16446_ obsg2.obstacleArray\[71\] _02059_ net399 _02124_ vssd1 vssd1 vccd1 vccd1
+ _02125_ sky130_fd_sc_hd__o211a_1
XFILLER_0_67_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_136_4475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_136_4486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_45_1681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_45_1692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_132_4339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12609_ net665 _07506_ vssd1 vssd1 vccd1 vccd1 _07507_ sky130_fd_sc_hd__nor2_1
XFILLER_0_137_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16377_ _02053_ _02054_ net433 vssd1 vssd1 vccd1 vccd1 _02056_ sky130_fd_sc_hd__a21o_1
X_19165_ clknet_leaf_52_clk _00109_ net1364 vssd1 vssd1 vccd1 vccd1 ag2.body\[28\]
+ sky130_fd_sc_hd__dfrtp_4
X_13589_ _03960_ control.divider.count\[7\] control.divider.count\[9\] _03961_ control.divider.count\[8\]
+ vssd1 vssd1 vccd1 vccd1 _07964_ sky130_fd_sc_hd__o221a_1
Xclkbuf_leaf_11_clk clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_11_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_121_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_1567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18116_ net300 _03630_ vssd1 vssd1 vccd1 vccd1 _03693_ sky130_fd_sc_hd__nand2_1
XFILLER_0_14_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15328_ net2639 net73 _01587_ control.body\[696\] vssd1 vssd1 vccd1 vccd1 _00626_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_41_1578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_847 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19096_ clknet_leaf_146_clk img_gen.tracker.next_frame\[534\] net1239 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[534\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__10964__A1 net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18047_ net42 _03647_ vssd1 vssd1 vccd1 vccd1 _03648_ sky130_fd_sc_hd__nor2_1
X_15259_ net2629 net108 net50 control.body\[765\] vssd1 vssd1 vccd1 vccd1 _00567_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__16271__S net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12166__B1 net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09674__A net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_91_3092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_1479 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11913__B1 net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12812__B _07607_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout407 net408 vssd1 vssd1 vccd1 vccd1 net407 sky130_fd_sc_hd__clkbuf_4
XANTENNA__13196__A net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09820_ net750 control.body\[1054\] control.body\[1053\] net755 vssd1 vssd1 vccd1
+ vccd1 _04793_ sky130_fd_sc_hd__a2bb2o_1
Xfanout418 net419 vssd1 vssd1 vccd1 vccd1 net418 sky130_fd_sc_hd__buf_4
XANTENNA__17891__A net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10172__X _05145_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19998_ clknet_leaf_64_clk _00942_ net1475 vssd1 vssd1 vccd1 vccd1 ag2.body\[396\]
+ sky130_fd_sc_hd__dfrtp_4
Xfanout429 _01735_ vssd1 vssd1 vccd1 vccd1 net429 sky130_fd_sc_hd__clkbuf_2
XANTENNA__11087__A_N net1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16852__B1 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09751_ ag2.body\[211\] net1162 vssd1 vssd1 vccd1 vccd1 _04724_ sky130_fd_sc_hd__or2_1
XANTENNA__11428__B net1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18949_ clknet_leaf_5_clk img_gen.tracker.next_frame\[387\] net1269 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[387\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__13666__B1 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_78_clk clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_78_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_119_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09682_ _04652_ _04653_ _04654_ vssd1 vssd1 vccd1 vccd1 _04655_ sky130_fd_sc_hd__or3_2
XFILLER_0_59_1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_96_508 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17115__B net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout170_A net171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11692__A2 net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_102_3420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16080__A1 net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_3431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11444__A net1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout268_A net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_3442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16954__B net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17769__C _03446_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout435_A net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14755__A net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout36 _03706_ vssd1 vssd1 vccd1 vccd1 net36 sky130_fd_sc_hd__buf_4
XANTENNA_fanout1177_A net1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout47 net48 vssd1 vssd1 vccd1 vccd1 net47 sky130_fd_sc_hd__buf_2
XFILLER_0_9_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_1152 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout58 net59 vssd1 vssd1 vccd1 vccd1 net58 sky130_fd_sc_hd__buf_8
XTAP_TAPCELL_ROW_119_3950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout69 net70 vssd1 vssd1 vccd1 vccd1 net69 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_119_3961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_315 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14394__A1 net1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout223_X net223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14394__B2 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_115_3825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout602_A _06476_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09568__B net1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_115_3836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1344_A net1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09116_ ag2.body\[390\] vssd1 vssd1 vccd1 vccd1 _04141_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_21_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15343__B1 _01590_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09047_ ag2.body\[235\] vssd1 vssd1 vccd1 vccd1 _04072_ sky130_fd_sc_hd__inv_2
XANTENNA__14490__A net1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16181__S net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1511_A net9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1132_X net1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14921__C net66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13818__B _08114_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold450 img_gen.tracker.frame\[545\] vssd1 vssd1 vccd1 vccd1 net2012 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout971_A net974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold461 img_gen.tracker.frame\[181\] vssd1 vssd1 vccd1 vccd1 net2023 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout592_X net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold472 img_gen.tracker.frame\[142\] vssd1 vssd1 vccd1 vccd1 net2034 sky130_fd_sc_hd__dlygate4sd3_1
X_20207_ clknet_leaf_56_clk _01151_ net1457 vssd1 vssd1 vccd1 vccd1 ag2.body\[189\]
+ sky130_fd_sc_hd__dfrtp_4
Xhold483 img_gen.tracker.frame\[572\] vssd1 vssd1 vccd1 vccd1 net2045 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold494 img_gen.tracker.frame\[11\] vssd1 vssd1 vccd1 vccd1 net2056 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__19850__CLK clknet_leaf_93_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_8_Left_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10523__A _05419_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_2453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout83_A net91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_2464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout930 net931 vssd1 vssd1 vccd1 vccd1 net930 sky130_fd_sc_hd__buf_4
XFILLER_0_99_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout941 obsg2.randCord\[6\] vssd1 vssd1 vccd1 vccd1 net941 sky130_fd_sc_hd__buf_4
Xfanout952 net955 vssd1 vssd1 vccd1 vccd1 net952 sky130_fd_sc_hd__buf_4
X_09949_ _04919_ _04920_ _04921_ _04918_ vssd1 vssd1 vccd1 vccd1 _04922_ sky130_fd_sc_hd__a211o_1
X_20138_ clknet_leaf_97_clk _01082_ net1450 vssd1 vssd1 vccd1 vccd1 ag2.body\[248\]
+ sky130_fd_sc_hd__dfrtp_4
Xfanout963 net968 vssd1 vssd1 vccd1 vccd1 net963 sky130_fd_sc_hd__clkbuf_8
XANTENNA__14489__X _08650_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_69_clk clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_69_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout857_X net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10242__B net1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11117__D1 control.body_update.curr_length\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout974 ag2.randCord\[3\] vssd1 vssd1 vccd1 vccd1 net974 sky130_fd_sc_hd__buf_4
Xfanout985 net986 vssd1 vssd1 vccd1 vccd1 net985 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_5_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20069_ clknet_leaf_73_clk _01013_ net1501 vssd1 vssd1 vccd1 vccd1 ag2.body\[323\]
+ sky130_fd_sc_hd__dfrtp_4
Xfanout996 net1005 vssd1 vssd1 vccd1 vccd1 net996 sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_5_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12960_ net232 _07676_ _07677_ net1910 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[240\]
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_5_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11911_ img_gen.tracker.frame\[337\] net615 net598 img_gen.tracker.frame\[340\] vssd1
+ vssd1 vccd1 vccd1 _06883_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_87_2972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17025__B net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09750__C _04719_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_2983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11683__A2 net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12880__A1 net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12891_ _07443_ _07639_ vssd1 vssd1 vccd1 vccd1 _07645_ sky130_fd_sc_hd__nor2_1
XANTENNA__15949__A2 net195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_68_2382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14630_ net842 ag2.body\[464\] ag2.body\[466\] net825 _08790_ vssd1 vssd1 vccd1 vccd1
+ _08791_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_83_2847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_2393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_2858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11842_ img_gen.tracker.frame\[491\] net583 net547 img_gen.tracker.frame\[488\] _06813_
+ vssd1 vssd1 vccd1 vccd1 _06814_ sky130_fd_sc_hd__o221a_1
XFILLER_0_115_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_2869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12169__B net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_2268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14561_ _08717_ _08719_ _08721_ vssd1 vssd1 vccd1 vccd1 _08722_ sky130_fd_sc_hd__or3_1
XFILLER_0_51_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_2279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16359__C1 _01911_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19230__CLK clknet_leaf_75_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11773_ img_gen.tracker.frame\[83\] net588 net550 img_gen.tracker.frame\[80\] _06744_
+ vssd1 vssd1 vccd1 vccd1 _06745_ sky130_fd_sc_hd__o221a_1
XANTENNA__12093__C1 net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16356__S net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14665__A net1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12737__X _07572_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18137__A net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17020__B1 net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16300_ _01912_ _01970_ _01977_ _01978_ _01918_ vssd1 vssd1 vccd1 vccd1 _01979_ sky130_fd_sc_hd__a221o_1
XANTENNA_clkbuf_leaf_142_clk_X clknet_leaf_142_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13512_ net1685 _07916_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[553\]
+ sky130_fd_sc_hd__and2_1
XANTENNA__09759__A ag2.body\[214\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10724_ net906 net639 net902 vssd1 vssd1 vccd1 vccd1 _05697_ sky130_fd_sc_hd__a21o_1
X_17280_ ag2.body\[554\] net723 net929 _04205_ _02951_ vssd1 vssd1 vccd1 vccd1 _02959_
+ sky130_fd_sc_hd__a221o_1
X_14492_ net1023 _04124_ _04125_ net1013 _08646_ vssd1 vssd1 vccd1 vccd1 _08653_ sky130_fd_sc_hd__a221o_1
XANTENNA__11986__A3 _06951_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16231_ net415 _01909_ net371 _01904_ vssd1 vssd1 vccd1 vccd1 _01910_ sky130_fd_sc_hd__a211o_1
XFILLER_0_10_1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14385__A1 net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_22_clk_X clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13443_ net256 _07888_ _07889_ net1799 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[511\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__09478__B net1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14385__B2 net1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17976__A net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10655_ ag2.body\[282\] net1187 vssd1 vssd1 vccd1 vccd1 _05628_ sky130_fd_sc_hd__xor2_1
XANTENNA__12185__A net1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11199__A1 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_1570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12396__B1 net241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11199__B2 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16162_ obsg2.obstacleArray\[9\] net431 vssd1 vssd1 vccd1 vccd1 _01841_ sky130_fd_sc_hd__or2_1
X_13374_ net234 _07862_ _07863_ net2018 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[468\]
+ sky130_fd_sc_hd__a22o_1
Xclkload17 clknet_leaf_7_clk vssd1 vssd1 vccd1 vccd1 clkload17/Y sky130_fd_sc_hd__inv_8
X_10586_ _04425_ net637 _04494_ vssd1 vssd1 vccd1 vccd1 _05559_ sky130_fd_sc_hd__o21a_1
Xclkload28 clknet_leaf_133_clk vssd1 vssd1 vccd1 vccd1 clkload28/Y sky130_fd_sc_hd__inv_8
XFILLER_0_23_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10417__B net1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_1456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15113_ control.body\[898\] net146 _01554_ control.body\[890\] vssd1 vssd1 vccd1
+ vccd1 _00436_ sky130_fd_sc_hd__a22o_1
Xclkload39 clknet_leaf_126_clk vssd1 vssd1 vccd1 vccd1 clkload39/Y sky130_fd_sc_hd__clkinv_16
X_12325_ _07242_ _07245_ vssd1 vssd1 vccd1 vccd1 _07292_ sky130_fd_sc_hd__and2b_1
XFILLER_0_2_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18948__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16093_ obsg2.obstacleArray\[116\] obsg2.obstacleArray\[117\] net425 vssd1 vssd1
+ vccd1 vccd1 _01772_ sky130_fd_sc_hd__mux2_1
XANTENNA__12148__B1 net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15885__A1 ag2.body\[209\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_37_clk_X clknet_leaf_37_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19921_ clknet_leaf_55_clk _00865_ net1456 vssd1 vssd1 vccd1 vccd1 ag2.body\[479\]
+ sky130_fd_sc_hd__dfrtp_4
X_15044_ net2296 net150 _01556_ net2380 vssd1 vssd1 vccd1 vccd1 _00374_ sky130_fd_sc_hd__a22o_1
X_12256_ img_gen.updater.commands.cmd_num\[4\] _07198_ _07225_ _07197_ vssd1 vssd1
+ vccd1 vccd1 _07226_ sky130_fd_sc_hd__a22o_1
XANTENNA__12699__A1 net237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12632__B net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17087__B1 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11207_ _04555_ _05254_ vssd1 vssd1 vccd1 vccd1 _06180_ sky130_fd_sc_hd__nor2_1
X_19852_ clknet_leaf_92_clk _00796_ net1413 vssd1 vssd1 vccd1 vccd1 ag2.body\[538\]
+ sky130_fd_sc_hd__dfrtp_4
X_12187_ net1102 ag2.apple_cord\[5\] vssd1 vssd1 vccd1 vccd1 _07159_ sky130_fd_sc_hd__or2_1
XANTENNA__10433__A net1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_125_4121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18803_ clknet_leaf_3_clk img_gen.tracker.next_frame\[241\] net1260 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[241\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_43_1197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_1950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11138_ _05152_ _06110_ vssd1 vssd1 vccd1 vccd1 _06111_ sky130_fd_sc_hd__and2_1
XANTENNA__11248__B net1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19783_ clknet_leaf_127_clk _00727_ net1326 vssd1 vssd1 vccd1 vccd1 ag2.body\[613\]
+ sky130_fd_sc_hd__dfrtp_4
X_16995_ ag2.body\[137\] net877 vssd1 vssd1 vccd1 vccd1 _02674_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_34_1360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18734_ clknet_leaf_142_clk img_gen.tracker.next_frame\[172\] net1257 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[172\] sky130_fd_sc_hd__dfrtp_1
X_15946_ _04832_ net61 vssd1 vssd1 vccd1 vccd1 _01656_ sky130_fd_sc_hd__nor2_2
X_11069_ ag2.body\[366\] net1088 vssd1 vssd1 vccd1 vccd1 _06042_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_92_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_0_clk clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_0_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_30_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14876__A_N _04859_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19987__RESET_B net1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18665_ clknet_leaf_11_clk img_gen.tracker.next_frame\[103\] net1281 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[103\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_4_5__f_clk_X clknet_4_5__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16598__C1 net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19204__Q ag2.body\[67\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15877_ ag2.body\[218\] net188 _01648_ ag2.body\[210\] vssd1 vssd1 vccd1 vccd1 _01116_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_118_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17616_ _03292_ _03293_ _03294_ vssd1 vssd1 vccd1 vccd1 _03295_ sky130_fd_sc_hd__or3_1
X_14828_ _01494_ _01495_ _01498_ vssd1 vssd1 vccd1 vccd1 _01499_ sky130_fd_sc_hd__or3_1
XFILLER_0_59_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_138_4526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18596_ clknet_leaf_14_clk img_gen.tracker.next_frame\[34\] net1276 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[34\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_138_4537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_1102 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_4559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17547_ ag2.body\[323\] net856 vssd1 vssd1 vccd1 vccd1 _03226_ sky130_fd_sc_hd__xor2_1
XANTENNA__12623__A1 net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11426__A2 _04982_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14575__A net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_1765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14759_ net817 ag2.body\[43\] _03990_ net1006 _08919_ vssd1 vssd1 vccd1 vccd1 _08920_
+ sky130_fd_sc_hd__o221a_1
XANTENNA__18047__A net42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_1461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17478_ ag2.body\[134\] net944 vssd1 vssd1 vccd1 vccd1 _03157_ sky130_fd_sc_hd__or2_1
XANTENNA__19723__CLK clknet_leaf_132_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_15_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_15_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14376__A1 net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19217_ clknet_leaf_67_clk _00161_ net1494 vssd1 vssd1 vccd1 vccd1 ag2.body\[80\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__14376__B2 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16429_ obsg2.obstacleArray\[74\] obsg2.obstacleArray\[75\] net453 vssd1 vssd1 vccd1
+ vccd1 _02108_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10608__A net1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_994 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_3290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12526__C net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19148_ clknet_leaf_51_clk _00092_ net1367 vssd1 vssd1 vccd1 vccd1 ag2.body\[12\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__15677__Y _01627_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_3154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_3165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14128__A1 net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_1210 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14128__B2 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19079_ clknet_leaf_29_clk img_gen.tracker.next_frame\[517\] net1334 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[517\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__12823__A net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15876__B2 ag2.body\[209\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17078__B1 net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17617__A2 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1530 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout204 net218 vssd1 vssd1 vccd1 vccd1 net204 sky130_fd_sc_hd__clkbuf_2
Xfanout215 net216 vssd1 vssd1 vccd1 vccd1 net215 sky130_fd_sc_hd__buf_2
XANTENNA__19103__CLK clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout226 net227 vssd1 vssd1 vccd1 vccd1 net226 sky130_fd_sc_hd__clkbuf_4
XANTENNA__16949__B net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09803_ net1087 control.body\[966\] vssd1 vssd1 vccd1 vccd1 _04776_ sky130_fd_sc_hd__or2_1
Xfanout237 net238 vssd1 vssd1 vccd1 vccd1 net237 sky130_fd_sc_hd__clkbuf_4
Xfanout248 _07317_ vssd1 vssd1 vccd1 vccd1 net248 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_22_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11158__B net1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout259 net260 vssd1 vssd1 vccd1 vccd1 net259 sky130_fd_sc_hd__clkbuf_4
XANTENNA__14836__C1 _08467_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09734_ _04019_ net1163 net1064 _04022_ vssd1 vssd1 vccd1 vccd1 _04707_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_104_3504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09858__A2 _04470_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09665_ _04425_ _04637_ vssd1 vssd1 vccd1 vccd1 _04638_ sky130_fd_sc_hd__and2_2
XANTENNA__12862__A1 net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout552_A net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11174__A net1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09596_ _04557_ _04564_ _04565_ _04568_ vssd1 vssd1 vccd1 vccd1 _04569_ sky130_fd_sc_hd__or4_2
XFILLER_0_136_1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_96_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__20230__CLK clknet_leaf_66_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout340_X net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16029__X _01708_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14485__A net1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout817_A net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1461_A net1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1082_X net1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17002__B1 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout438_X net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10625__B1 net1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09579__A net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12090__A2 net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14367__A1 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14367__B2 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout605_X net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_808 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10440_ net1133 control.body\[932\] vssd1 vssd1 vccd1 vccd1 _05413_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_45_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10237__B net1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20144__RESET_B net1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_2640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10928__B2 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11050__B1 net1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_2651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16513__C1 net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10371_ net783 control.body\[760\] control.body\[762\] net773 vssd1 vssd1 vccd1 vccd1
+ _05344_ sky130_fd_sc_hd__a22o_1
XFILLER_0_61_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12733__A net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_2504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_2050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12110_ img_gen.tracker.frame\[180\] net628 net555 img_gen.tracker.frame\[186\] _07081_
+ vssd1 vssd1 vccd1 vccd1 _07082_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_57_2061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_2072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_351 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13090_ net243 _07737_ _07738_ net1687 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[309\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout974_X net974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12041_ net576 _07012_ _07010_ net474 vssd1 vssd1 vccd1 vccd1 _07013_ sky130_fd_sc_hd__a211o_1
Xhold280 img_gen.tracker.frame\[402\] vssd1 vssd1 vccd1 vccd1 net1842 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold291 img_gen.tracker.frame\[459\] vssd1 vssd1 vccd1 vccd1 net1853 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17962__C _03586_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout760 net766 vssd1 vssd1 vccd1 vccd1 net760 sky130_fd_sc_hd__clkbuf_4
X_15800_ ag2.body\[293\] net210 _01640_ ag2.body\[285\] vssd1 vssd1 vccd1 vccd1 _01047_
+ sky130_fd_sc_hd__a22o_1
Xfanout771 _04230_ vssd1 vssd1 vccd1 vccd1 net771 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09761__B net1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout782 _04228_ vssd1 vssd1 vccd1 vccd1 net782 sky130_fd_sc_hd__buf_4
X_13992_ ag2.body\[128\] net213 _08160_ ag2.body\[120\] vssd1 vssd1 vccd1 vccd1 _00209_
+ sky130_fd_sc_hd__a22o_1
X_16780_ _02403_ _02458_ net350 vssd1 vssd1 vccd1 vccd1 _02459_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_85_2909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout793 net797 vssd1 vssd1 vccd1 vccd1 net793 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09849__A2 _04607_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15731_ _05657_ net60 vssd1 vssd1 vccd1 vccd1 _01633_ sky130_fd_sc_hd__nor2_2
X_12943_ img_gen.tracker.frame\[232\] net662 vssd1 vssd1 vccd1 vccd1 _07669_ sky130_fd_sc_hd__and2_1
XANTENNA__10700__B net1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1610 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_64_clk_A clknet_4_13__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18450_ _04645_ _03826_ _03938_ _03824_ vssd1 vssd1 vccd1 vccd1 _03939_ sky130_fd_sc_hd__o211a_1
XANTENNA__10864__B1 _05836_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15662_ ag2.body\[410\] net143 _01625_ ag2.body\[402\] vssd1 vssd1 vccd1 vccd1 _00924_
+ sky130_fd_sc_hd__a22o_1
X_12874_ net292 _07636_ _07637_ net1638 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[194\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_62_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17401_ ag2.body\[45\] net946 vssd1 vssd1 vccd1 vccd1 _03080_ sky130_fd_sc_hd__xor2_1
X_14613_ net996 ag2.body\[56\] vssd1 vssd1 vccd1 vccd1 _08774_ sky130_fd_sc_hd__xor2_1
X_11825_ img_gen.tracker.frame\[422\] net616 net545 img_gen.tracker.frame\[428\] vssd1
+ vssd1 vccd1 vccd1 _06797_ sky130_fd_sc_hd__o22a_1
X_15593_ ag2.body\[476\] net122 _01618_ ag2.body\[468\] vssd1 vssd1 vccd1 vccd1 _00862_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_90_1471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12605__A1 net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18381_ _08051_ _03800_ _03869_ vssd1 vssd1 vccd1 vccd1 _03871_ sky130_fd_sc_hd__nand3_1
XANTENNA__16086__S net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_1444 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17332_ _03974_ net930 vssd1 vssd1 vccd1 vccd1 _03011_ sky130_fd_sc_hd__nor2_1
XFILLER_0_95_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14544_ net1030 _04077_ _04078_ net1010 _08704_ vssd1 vssd1 vccd1 vccd1 _08705_ sky130_fd_sc_hd__a221o_2
XFILLER_0_95_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11756_ img_gen.tracker.frame\[257\] _06476_ net581 img_gen.tracker.frame\[263\]
+ vssd1 vssd1 vccd1 vccd1 _06728_ sky130_fd_sc_hd__o22a_1
XANTENNA__09482__B1 net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12081__A2 net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_79_clk_A clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12627__B net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14358__A1 net994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10707_ ag2.body\[17\] net1197 vssd1 vssd1 vccd1 vccd1 _05680_ sky130_fd_sc_hd__xor2_1
XFILLER_0_3_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14358__B2 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14475_ net1016 ag2.body\[446\] vssd1 vssd1 vccd1 vccd1 _08636_ sky130_fd_sc_hd__xor2_1
XANTENNA__18770__CLK clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17263_ ag2.body\[251\] net719 net699 ag2.body\[254\] vssd1 vssd1 vccd1 vccd1 _02942_
+ sky130_fd_sc_hd__a22o_1
X_11687_ net1070 net743 vssd1 vssd1 vccd1 vccd1 _06659_ sky130_fd_sc_hd__nor2_2
XANTENNA__10428__A net1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_122_clk_A clknet_4_9__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19002_ clknet_leaf_2_clk img_gen.tracker.next_frame\[440\] net1249 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[440\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12346__C net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16214_ net354 _01892_ vssd1 vssd1 vccd1 vccd1 _01893_ sky130_fd_sc_hd__nand2_1
X_13426_ net2060 net647 _07882_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[501\]
+ sky130_fd_sc_hd__and3_1
XFILLER_0_3_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10638_ net1145 control.body\[667\] vssd1 vssd1 vccd1 vccd1 _05611_ sky130_fd_sc_hd__xor2_1
XANTENNA__13030__A1 net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17194_ _02864_ _02866_ _02869_ _02872_ vssd1 vssd1 vccd1 vccd1 _02873_ sky130_fd_sc_hd__or4_1
XFILLER_0_125_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload106 clknet_leaf_56_clk vssd1 vssd1 vccd1 vccd1 clkload106/Y sky130_fd_sc_hd__inv_4
Xclkload117 clknet_leaf_64_clk vssd1 vssd1 vccd1 vccd1 clkload117/Y sky130_fd_sc_hd__clkinv_2
XANTENNA__10147__B net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkload128 clknet_leaf_69_clk vssd1 vssd1 vccd1 vccd1 clkload128/Y sky130_fd_sc_hd__inv_6
XANTENNA__14325__A1_N net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_1242 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16145_ obsg2.obstacleArray\[17\] net431 vssd1 vssd1 vccd1 vccd1 _01824_ sky130_fd_sc_hd__or2_1
X_13357_ net384 _07523_ vssd1 vssd1 vccd1 vccd1 _07856_ sky130_fd_sc_hd__nor2_1
XFILLER_0_49_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09936__B net1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10569_ _05535_ _05539_ _05540_ _05541_ vssd1 vssd1 vccd1 vccd1 _05542_ sky130_fd_sc_hd__or4b_1
XFILLER_0_87_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19126__CLK clknet_leaf_131_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12308_ _07222_ _07273_ vssd1 vssd1 vccd1 vccd1 _07275_ sky130_fd_sc_hd__nor2_1
X_16076_ net375 _01752_ _01754_ net348 vssd1 vssd1 vccd1 vccd1 _01755_ sky130_fd_sc_hd__a211o_1
X_13288_ _07472_ net303 vssd1 vssd1 vccd1 vccd1 _07829_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_127_4205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_137_clk_A clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19904_ clknet_leaf_86_clk _00848_ net1464 vssd1 vssd1 vccd1 vccd1 ag2.body\[494\]
+ sky130_fd_sc_hd__dfrtp_4
X_15027_ control.body\[981\] net167 _01555_ control.body\[973\] vssd1 vssd1 vccd1
+ vccd1 _00359_ sky130_fd_sc_hd__a22o_1
XFILLER_0_23_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12239_ _07195_ _07203_ vssd1 vssd1 vccd1 vccd1 _07209_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_36_1422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_1433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_17_clk_A clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16807__B1 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19835_ clknet_leaf_92_clk _00779_ net1414 vssd1 vssd1 vccd1 vccd1 ag2.body\[553\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_97_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_1609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19766_ clknet_leaf_130_clk _00710_ net1326 vssd1 vssd1 vccd1 vccd1 control.body\[628\]
+ sky130_fd_sc_hd__dfrtp_1
X_16978_ ag2.body\[425\] net871 vssd1 vssd1 vccd1 vccd1 _02657_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_36_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput4 gpio_in[27] vssd1 vssd1 vccd1 vccd1 net4 sky130_fd_sc_hd__clkbuf_1
X_18717_ clknet_leaf_144_clk img_gen.tracker.next_frame\[155\] net1252 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[155\] sky130_fd_sc_hd__dfrtp_1
X_15929_ _05922_ net57 vssd1 vssd1 vccd1 vccd1 _01655_ sky130_fd_sc_hd__nor2_2
X_19697_ clknet_leaf_136_clk _00641_ net1300 vssd1 vssd1 vccd1 vccd1 control.body\[703\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_49_1805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16785__A net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11125__A_N net1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17232__B1 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_49_1827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09450_ net920 net916 vssd1 vssd1 vccd1 vccd1 _04423_ sky130_fd_sc_hd__nand2_1
X_18648_ clknet_leaf_130_clk img_gen.tracker.next_frame\[86\] net1315 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[86\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16586__A2 net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14597__A1 net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09381_ sound_gen.osc1.stayCount\[13\] _04357_ net271 vssd1 vssd1 vccd1 vccd1 _04375_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_133_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14597__B2 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18579_ clknet_leaf_4_clk img_gen.tracker.next_frame\[17\] net1278 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[17\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__12818__A net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_3330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20610_ net1542 vssd1 vssd1 vccd1 vccd1 gpio_oeb[22] sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_99_3341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_3352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12072__A2 net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkload72_A clknet_leaf_113_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_95_3216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_3227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20541_ clknet_leaf_105_clk _01406_ _00015_ vssd1 vssd1 vccd1 vccd1 sound_gen.osc1.stayCount\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__16724__S net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout133_A net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20472_ clknet_leaf_33_clk _01359_ net1346 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[108\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_6_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17766__D _03444_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18224__B net40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_89_Left_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout300_A net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12553__A net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09565__C _04519_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10073__A net1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18240__A _03681_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout290_X net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11886__A2 net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout388_X net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout767_A net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19838__RESET_B net1414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18643__CLK clknet_leaf_141_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19769__CLK clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_98_Left_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09717_ _04076_ net1207 net1062 _04078_ _04689_ vssd1 vssd1 vccd1 vccd1 _04690_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout934_A net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout555_X net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09648_ net1172 control.body\[746\] vssd1 vssd1 vccd1 vccd1 _04621_ sky130_fd_sc_hd__xor2_1
XANTENNA__10310__A2 _04640_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14588__A1 net994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14588__B2 net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout722_X net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09579_ net895 _04550_ vssd1 vssd1 vccd1 vccd1 _04552_ sky130_fd_sc_hd__or2_1
XANTENNA__18793__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11054__D _04429_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1464_X net1464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12728__A net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11610_ net508 _06579_ _06582_ vssd1 vssd1 vccd1 vccd1 _06583_ sky130_fd_sc_hd__o21a_1
XFILLER_0_77_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12590_ net230 net308 _07495_ _07496_ net1643 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[51\]
+ sky130_fd_sc_hd__a32o_1
XANTENNA__13260__A1 net236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09464__B1 net1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_330 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1331 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11351__B net1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11541_ _06512_ _06513_ net506 vssd1 vssd1 vccd1 vccd1 _06514_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_2702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_2713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_1584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17957__C _03582_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09596__X _04569_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14260_ net845 ag2.body\[72\] _04007_ net1040 _08415_ vssd1 vssd1 vccd1 vccd1 _08421_
+ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_59_2112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11472_ ag2.body\[494\] net1089 vssd1 vssd1 vccd1 vccd1 _06445_ sky130_fd_sc_hd__xor2_1
XANTENNA__13012__A1 net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_59_2123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08941__A net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15758__B net60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_2134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18134__B net41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13211_ net263 _07794_ _07795_ net1619 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[373\]
+ sky130_fd_sc_hd__a22o_1
Xwire479 _05049_ vssd1 vssd1 vccd1 vccd1 net479 sky130_fd_sc_hd__buf_1
X_10423_ net779 control.body\[1065\] control.body\[1067\] net769 vssd1 vssd1 vccd1
+ vccd1 _05396_ sky130_fd_sc_hd__o2bb2a_1
X_14191_ net974 ag2.body\[163\] vssd1 vssd1 vccd1 vccd1 _08352_ sky130_fd_sc_hd__xor2_1
XANTENNA__09756__B net1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14760__A1 net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_2009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14760__B2 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13142_ net232 _07762_ _07763_ net1863 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[336\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_103_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10354_ ag2.body\[294\] net1091 vssd1 vssd1 vccd1 vccd1 _05327_ sky130_fd_sc_hd__and2b_1
XFILLER_0_131_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17950_ net318 net47 net296 _03577_ obsg2.obstacleArray\[8\] vssd1 vssd1 vccd1 vccd1
+ _03578_ sky130_fd_sc_hd__a41o_1
X_13073_ net243 _07729_ _07730_ net1708 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[300\]
+ sky130_fd_sc_hd__a22o_1
X_10285_ ag2.body\[335\] net1067 vssd1 vssd1 vccd1 vccd1 _05258_ sky130_fd_sc_hd__nand2_1
Xfanout1500 net1502 vssd1 vssd1 vccd1 vccd1 net1500 sky130_fd_sc_hd__clkbuf_4
X_12024_ net1219 net1195 img_gen.tracker.frame\[213\] vssd1 vssd1 vccd1 vccd1 _06996_
+ sky130_fd_sc_hd__and3_1
X_16901_ ag2.body\[244\] net711 net933 _04078_ vssd1 vssd1 vccd1 vccd1 _02580_ sky130_fd_sc_hd__a2bb2o_1
Xfanout1511 net9 vssd1 vssd1 vccd1 vccd1 net1511 sky130_fd_sc_hd__clkbuf_2
X_17881_ _04397_ _03520_ vssd1 vssd1 vccd1 vccd1 _03521_ sky130_fd_sc_hd__nor2_2
XANTENNA__12910__B net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19620_ clknet_leaf_123_clk _00564_ net1406 vssd1 vssd1 vccd1 vccd1 control.body\[770\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13294__A net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09491__B net1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16832_ ag2.body\[96\] net885 vssd1 vssd1 vccd1 vccd1 _02511_ sky130_fd_sc_hd__xnor2_1
XANTENNA__19579__RESET_B net1386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout590 net591 vssd1 vssd1 vccd1 vccd1 net590 sky130_fd_sc_hd__clkbuf_4
X_19551_ clknet_leaf_115_clk _00495_ net1397 vssd1 vssd1 vccd1 vccd1 control.body\[845\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_92_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16763_ obsg2.obstacleArray\[0\] net493 net488 obsg2.obstacleArray\[2\] vssd1 vssd1
+ vccd1 vccd1 _02442_ sky130_fd_sc_hd__a22o_1
XFILLER_0_73_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12826__A1 net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13975_ ag2.body\[113\] net202 _08158_ ag2.body\[105\] vssd1 vssd1 vccd1 vccd1 _00194_
+ sky130_fd_sc_hd__a22o_1
X_18502_ net1513 net1507 vssd1 vssd1 vccd1 vccd1 _00033_ sky130_fd_sc_hd__or2_1
XANTENNA__17214__B1 net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15714_ ag2.body\[361\] net193 _01630_ ag2.body\[353\] vssd1 vssd1 vccd1 vccd1 _00971_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_87_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19482_ clknet_leaf_114_clk _00426_ net1400 vssd1 vssd1 vccd1 vccd1 control.body\[904\]
+ sky130_fd_sc_hd__dfrtp_1
X_12926_ img_gen.tracker.frame\[223\] net652 vssd1 vssd1 vccd1 vccd1 _07661_ sky130_fd_sc_hd__and2_1
X_16694_ net709 net538 vssd1 vssd1 vccd1 vccd1 _02373_ sky130_fd_sc_hd__nor2_2
XFILLER_0_88_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_1648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14579__A1 net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18433_ _03802_ _03805_ _03795_ vssd1 vssd1 vccd1 vccd1 _03922_ sky130_fd_sc_hd__a21oi_1
X_15645_ ag2.body\[427\] net126 _01623_ ag2.body\[419\] vssd1 vssd1 vccd1 vccd1 _00909_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__14579__B2 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17213__B net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12857_ net287 _07628_ _07629_ net1864 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[185\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_115_1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18028__C net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_842 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18364_ net1981 _08024_ _03854_ _03858_ vssd1 vssd1 vccd1 vccd1 _01392_ sky130_fd_sc_hd__o22a_1
X_11808_ img_gen.tracker.frame\[446\] net614 net568 _06779_ vssd1 vssd1 vccd1 vccd1
+ _06780_ sky130_fd_sc_hd__o211a_1
XFILLER_0_115_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15576_ ag2.body\[494\] net135 _01615_ ag2.body\[486\] vssd1 vssd1 vccd1 vccd1 _00848_
+ sky130_fd_sc_hd__a22o_1
X_12788_ net261 _07596_ _07597_ net1818 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[148\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_51_1274 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17315_ _02985_ _02988_ _02992_ _02993_ vssd1 vssd1 vccd1 vccd1 _02994_ sky130_fd_sc_hd__or4b_2
XFILLER_0_138_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11739_ img_gen.tracker.frame\[14\] net623 vssd1 vssd1 vccd1 vccd1 _06711_ sky130_fd_sc_hd__or2_1
X_14527_ _08684_ _08685_ _08686_ _08687_ vssd1 vssd1 vccd1 vccd1 _08688_ sky130_fd_sc_hd__a22o_1
XFILLER_0_71_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18295_ net325 net324 net322 track.nextHighScore\[6\] track.nextHighScore\[7\] vssd1
+ vssd1 vccd1 vccd1 _03791_ sky130_fd_sc_hd__a41o_1
XANTENNA__18190__A1 _01703_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17246_ ag2.body\[617\] net730 net858 _04223_ vssd1 vssd1 vccd1 vccd1 _02925_ sky130_fd_sc_hd__o22a_1
X_14458_ net842 ag2.body\[432\] ag2.body\[436\] net812 vssd1 vssd1 vccd1 vccd1 _08619_
+ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__15668__B net67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_975 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_761 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14751__A1 net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15020__Y _01554_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13409_ net281 _07874_ _07875_ net1681 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[491\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_113_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17177_ _02852_ _02853_ _02854_ _02855_ _02851_ vssd1 vssd1 vccd1 vccd1 _02856_ sky130_fd_sc_hd__a221o_1
XANTENNA__14751__B2 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14389_ net830 ag2.body\[298\] ag2.body\[296\] net844 vssd1 vssd1 vccd1 vccd1 _08550_
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_40_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16128_ obsg2.obstacleArray\[74\] net423 vssd1 vssd1 vccd1 vccd1 _01807_ sky130_fd_sc_hd__or2_1
XANTENNA__17883__B obsg2.obstacleCount\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08950_ ag2.body\[9\] vssd1 vssd1 vccd1 vccd1 _03975_ sky130_fd_sc_hd__inv_2
X_16059_ _01716_ _01725_ net538 vssd1 vssd1 vccd1 vccd1 _01738_ sky130_fd_sc_hd__a21oi_1
XANTENNA__18060__A net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_88_3020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_899 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_135_Right_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_1376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19818_ clknet_leaf_89_clk _00762_ net1411 vssd1 vssd1 vccd1 vccd1 ag2.body\[568\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_100_1555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19249__RESET_B net1482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11436__B net1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19749_ clknet_leaf_129_clk net2310 net1325 vssd1 vssd1 vccd1 vccd1 control.body\[643\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_79_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10340__B net1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09502_ ag2.body\[400\] net784 vssd1 vssd1 vccd1 vccd1 _04475_ sky130_fd_sc_hd__nor2_1
XFILLER_0_2_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09433_ net926 net1103 vssd1 vssd1 vccd1 vccd1 _04406_ sky130_fd_sc_hd__xor2_1
XFILLER_0_91_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17123__B net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout250_A net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09364_ sound_gen.osc1.stayCount\[14\] _04365_ vssd1 vssd1 vccd1 vccd1 _04366_ sky130_fd_sc_hd__and2_1
XFILLER_0_93_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12045__A2 net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09295_ _04314_ vssd1 vssd1 vccd1 vccd1 _04315_ sky130_fd_sc_hd__inv_2
XFILLER_0_30_1347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_503 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_20 _08509_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_31 _03442_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10068__A net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20149__CLK clknet_leaf_98_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1257_A net1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20524_ clknet_leaf_93_clk track.nextCurrScore\[6\] net1413 vssd1 vssd1 vccd1 vccd1
+ control.body_update.curr_length\[6\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_1557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15578__B net64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16731__A2 net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_878 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14742__A1 net1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20455_ clknet_leaf_39_clk _01342_ net1356 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[91\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA_fanout1045_X net1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20386_ clknet_leaf_43_clk _01273_ net1372 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[22\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA_fanout884_A net889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10515__B net1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16495__A1 net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17692__B1 net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1212_X net1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09592__A net1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18236__A2 net37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10070_ net1193 control.body\[713\] vssd1 vssd1 vccd1 vccd1 _05043_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout672_X net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_102_Right_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10531__A net1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14003__A net1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12808__A1 net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout937_X net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13842__A net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13760_ _08065_ _08074_ _08076_ net320 img_gen.updater.commands.count\[4\] vssd1
+ vssd1 vccd1 vccd1 _00061_ sky130_fd_sc_hd__a32o_1
XANTENNA__10819__B1 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10972_ net1083 control.body\[1006\] vssd1 vssd1 vccd1 vccd1 _05945_ sky130_fd_sc_hd__nor2_1
XFILLER_0_98_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12711_ net237 _07559_ _07560_ net1689 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[108\]
+ sky130_fd_sc_hd__a22o_1
X_13691_ net892 _08029_ vssd1 vssd1 vccd1 vccd1 _08033_ sky130_fd_sc_hd__nand2_1
XFILLER_0_35_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11362__A net1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12642_ net676 _07524_ vssd1 vssd1 vccd1 vccd1 _07525_ sky130_fd_sc_hd__nor2_1
X_15430_ ag2.body\[620\] net85 _01599_ ag2.body\[612\] vssd1 vssd1 vccd1 vccd1 _00718_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_17_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13233__A1 net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12036__A2 net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16970__A2 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16872__B net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15361_ net2272 net68 _01592_ control.body\[678\] vssd1 vssd1 vccd1 vccd1 _00656_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11081__B net1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12573_ net581 _06639_ net440 net559 vssd1 vssd1 vccd1 vccd1 _07486_ sky130_fd_sc_hd__or4_4
XANTENNA__14673__A net1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16364__S net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_1381 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17100_ _02774_ _02775_ _02776_ _02778_ vssd1 vssd1 vccd1 vccd1 _02779_ sky130_fd_sc_hd__a211o_1
XANTENNA__11795__A1 net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14312_ net971 ag2.body\[51\] vssd1 vssd1 vccd1 vccd1 _08473_ sky130_fd_sc_hd__xor2_1
X_11524_ _06495_ _06496_ vssd1 vssd1 vccd1 vccd1 _06497_ sky130_fd_sc_hd__and2_4
X_18080_ obsg2.obstacleArray\[46\] _03669_ net520 vssd1 vssd1 vccd1 vccd1 _01297_
+ sky130_fd_sc_hd__o21a_1
X_15292_ control.body\[736\] net77 _01585_ control.body\[728\] vssd1 vssd1 vccd1 vccd1
+ _00594_ sky130_fd_sc_hd__a22o_1
XFILLER_0_68_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15488__B net54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16722__A2 net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17031_ ag2.body\[402\] net865 vssd1 vssd1 vccd1 vccd1 _02710_ sky130_fd_sc_hd__xor2_1
X_14243_ net1031 ag2.body\[541\] vssd1 vssd1 vccd1 vccd1 _08404_ sky130_fd_sc_hd__xor2_1
XANTENNA__13289__A net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17984__A net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14733__A1 net1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09486__B net1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11455_ ag2.body\[261\] net1115 vssd1 vssd1 vccd1 vccd1 _06428_ sky130_fd_sc_hd__xor2_1
XANTENNA__14733__B2 net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11547__A1 _06485_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10406_ net1087 control.body\[1078\] vssd1 vssd1 vccd1 vccd1 _05379_ sky130_fd_sc_hd__xor2_1
XFILLER_0_61_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20183__Q ag2.body\[213\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14174_ net1014 ag2.body\[199\] vssd1 vssd1 vccd1 vccd1 _08335_ sky130_fd_sc_hd__nand2_1
X_11386_ net1073 control.body\[646\] vssd1 vssd1 vccd1 vccd1 _06359_ sky130_fd_sc_hd__nand2_1
X_13125_ _07754_ net265 _07752_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[328\]
+ sky130_fd_sc_hd__mux2_1
XANTENNA__17683__B1 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10337_ ag2.body\[526\] net1085 vssd1 vssd1 vccd1 vccd1 _05310_ sky130_fd_sc_hd__nand2_1
XFILLER_0_108_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18982_ clknet_leaf_8_clk img_gen.tracker.next_frame\[420\] net1270 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[420\] sky130_fd_sc_hd__dfrtp_1
X_17933_ _03549_ _03563_ _03564_ vssd1 vssd1 vccd1 vccd1 _03565_ sky130_fd_sc_hd__and3b_1
X_13056_ img_gen.tracker.frame\[292\] net660 vssd1 vssd1 vccd1 vccd1 _07722_ sky130_fd_sc_hd__and2_1
X_10268_ ag2.body\[139\] net1165 vssd1 vssd1 vccd1 vccd1 _05241_ sky130_fd_sc_hd__nand2_1
XANTENNA__17208__B net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1330 net1332 vssd1 vssd1 vccd1 vccd1 net1330 sky130_fd_sc_hd__clkbuf_2
X_12007_ img_gen.tracker.frame\[472\] net600 net545 img_gen.tracker.frame\[475\] _06978_
+ vssd1 vssd1 vccd1 vccd1 _06979_ sky130_fd_sc_hd__o221a_1
Xfanout1341 net1345 vssd1 vssd1 vccd1 vccd1 net1341 sky130_fd_sc_hd__clkbuf_2
Xfanout1352 net1356 vssd1 vssd1 vccd1 vccd1 net1352 sky130_fd_sc_hd__clkbuf_4
X_17864_ _03501_ _03513_ vssd1 vssd1 vccd1 vccd1 _01237_ sky130_fd_sc_hd__and2b_1
XANTENNA__10441__A net1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10199_ ag2.body\[117\] net1116 vssd1 vssd1 vccd1 vccd1 _05172_ sky130_fd_sc_hd__or2_1
Xfanout1363 net1364 vssd1 vssd1 vccd1 vccd1 net1363 sky130_fd_sc_hd__clkbuf_4
Xfanout1374 net1383 vssd1 vssd1 vccd1 vccd1 net1374 sky130_fd_sc_hd__clkbuf_4
X_19603_ clknet_leaf_119_clk _00547_ net1390 vssd1 vssd1 vccd1 vccd1 control.body\[785\]
+ sky130_fd_sc_hd__dfrtp_1
X_16815_ ag2.body\[84\] net966 vssd1 vssd1 vccd1 vccd1 _02494_ sky130_fd_sc_hd__xor2_1
Xfanout1385 net1386 vssd1 vssd1 vccd1 vccd1 net1385 sky130_fd_sc_hd__clkbuf_4
Xfanout1396 net1397 vssd1 vssd1 vccd1 vccd1 net1396 sky130_fd_sc_hd__clkbuf_4
X_17795_ _04261_ _03468_ vssd1 vssd1 vccd1 vccd1 _01214_ sky130_fd_sc_hd__xnor2_1
X_19534_ clknet_leaf_121_clk net2510 net1394 vssd1 vssd1 vccd1 vccd1 control.body\[860\]
+ sky130_fd_sc_hd__dfrtp_1
X_16746_ _02419_ _02424_ net380 vssd1 vssd1 vccd1 vccd1 _02425_ sky130_fd_sc_hd__mux2_1
XFILLER_0_92_1341 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13958_ ag2.body\[98\] net189 _08156_ ag2.body\[90\] vssd1 vssd1 vccd1 vccd1 _00179_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__17738__A1 _02632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13472__A1 net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19465_ clknet_leaf_109_clk _00409_ net1417 vssd1 vssd1 vccd1 vccd1 control.body\[935\]
+ sky130_fd_sc_hd__dfrtp_1
X_12909_ net2096 net661 _07315_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[214\]
+ sky130_fd_sc_hd__and3_1
XFILLER_0_53_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16677_ net358 _02321_ _02325_ _02317_ _02211_ vssd1 vssd1 vccd1 vccd1 _02356_ sky130_fd_sc_hd__a311o_1
X_13889_ ag2.body\[37\] net115 _08148_ ag2.body\[29\] vssd1 vssd1 vccd1 vccd1 _00118_
+ sky130_fd_sc_hd__a22o_1
X_18416_ _03844_ _03890_ vssd1 vssd1 vccd1 vccd1 _03906_ sky130_fd_sc_hd__nor2_1
X_15628_ ag2.body\[444\] net127 _01621_ ag2.body\[436\] vssd1 vssd1 vccd1 vccd1 _00894_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_31_1601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13224__A1 net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19396_ clknet_leaf_103_clk _00340_ net1428 vssd1 vssd1 vccd1 vccd1 control.body\[994\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__17878__B _03458_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18347_ _04420_ _06173_ _08025_ vssd1 vssd1 vccd1 vccd1 _03843_ sky130_fd_sc_hd__a21o_1
XANTENNA__16274__S net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15559_ _04686_ net56 vssd1 vssd1 vccd1 vccd1 _01613_ sky130_fd_sc_hd__nor2_2
XANTENNA__12655__X _07532_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14583__A net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18055__A net43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09080_ ag2.body\[314\] vssd1 vssd1 vccd1 vccd1 _04105_ sky130_fd_sc_hd__inv_2
XFILLER_0_83_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18278_ net319 net48 _03552_ _03577_ obsg2.obstacleArray\[136\] vssd1 vssd1 vccd1
+ vccd1 _03778_ sky130_fd_sc_hd__a41o_1
XFILLER_0_127_796 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17229_ ag2.body\[446\] net940 vssd1 vssd1 vccd1 vccd1 _02908_ sky130_fd_sc_hd__xor2_1
XFILLER_0_31_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold802 control.body\[688\] vssd1 vssd1 vccd1 vccd1 net2364 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09964__X _04937_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20240_ clknet_leaf_69_clk _01184_ net1496 vssd1 vssd1 vccd1 vccd1 ag2.body\[158\]
+ sky130_fd_sc_hd__dfrtp_4
Xhold813 control.body\[957\] vssd1 vssd1 vccd1 vccd1 net2375 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold824 control.body\[731\] vssd1 vssd1 vccd1 vccd1 net2386 sky130_fd_sc_hd__dlygate4sd3_1
Xhold835 _00670_ vssd1 vssd1 vccd1 vccd1 net2397 sky130_fd_sc_hd__dlygate4sd3_1
Xhold846 control.body\[965\] vssd1 vssd1 vccd1 vccd1 net2408 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkload35_A clknet_leaf_141_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10335__B net1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold857 control.body\[652\] vssd1 vssd1 vccd1 vccd1 net2419 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__17674__B1 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold868 _00460_ vssd1 vssd1 vccd1 vccd1 net2430 sky130_fd_sc_hd__dlygate4sd3_1
X_09982_ net787 control.body\[1112\] control.body\[1115\] net770 _04954_ vssd1 vssd1
+ vccd1 vccd1 _04955_ sky130_fd_sc_hd__a221o_1
X_20171_ clknet_leaf_82_clk _01115_ net1479 vssd1 vssd1 vccd1 vccd1 ag2.body\[217\]
+ sky130_fd_sc_hd__dfrtp_4
Xhold879 control.body\[675\] vssd1 vssd1 vccd1 vccd1 net2441 sky130_fd_sc_hd__dlygate4sd3_1
X_08933_ net2547 vssd1 vssd1 vccd1 vccd1 _03958_ sky130_fd_sc_hd__inv_2
XANTENNA__17118__B net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17426__B1 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09903__A1 _04863_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09903__B2 _04831_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10351__A ag2.body\[295\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_1236 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16449__S net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14758__A net1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13463__A1 net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1374_A net1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19807__CLK clknet_leaf_124_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09416_ _04261_ net686 vssd1 vssd1 vccd1 vccd1 _04395_ sky130_fd_sc_hd__nor2_1
XFILLER_0_137_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13215__A1 net240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09347_ _04346_ _04347_ _04349_ _04350_ vssd1 vssd1 vccd1 vccd1 _04351_ sky130_fd_sc_hd__and4_1
XFILLER_0_35_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout420_X net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16184__S net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09858__Y _04831_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1162_X net1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout518_X net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09587__A net1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09278_ sound_gen.osc1.stayCount\[21\] _04288_ _04299_ _04300_ vssd1 vssd1 vccd1
+ vccd1 _04301_ sky130_fd_sc_hd__o22a_1
XANTENNA__18831__CLK clknet_leaf_142_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17901__A1 _01691_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20507_ clknet_leaf_112_clk net1573 net1424 vssd1 vssd1 vccd1 vccd1 score_detect.sig_out\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__15912__B1 _01652_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10526__A net1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10423__A1_N net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11529__A1 net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11240_ ag2.body\[198\] net1080 vssd1 vssd1 vccd1 vccd1 _06213_ sky130_fd_sc_hd__nand2_1
XFILLER_0_121_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_1543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20438_ clknet_leaf_26_clk _01325_ net1343 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[74\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__10245__B net1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11624__S1 net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout887_X net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18981__CLK clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11171_ net1171 control.body\[778\] vssd1 vssd1 vccd1 vccd1 _06144_ sky130_fd_sc_hd__xor2_1
X_20369_ clknet_leaf_21_clk _01256_ net1360 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[5\]
+ sky130_fd_sc_hd__dfrtp_4
X_10122_ net1046 control.body\[711\] vssd1 vssd1 vccd1 vccd1 _05095_ sky130_fd_sc_hd__or2_1
XANTENNA__17028__B net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11357__A net1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10053_ _04429_ _04718_ _05024_ _05025_ vssd1 vssd1 vccd1 vccd1 _05026_ sky130_fd_sc_hd__nand4_2
X_14930_ _05364_ net59 vssd1 vssd1 vccd1 vccd1 _01544_ sky130_fd_sc_hd__nor2_2
XANTENNA__19337__CLK clknet_leaf_103_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16867__B net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14861_ _08516_ _08521_ _01529_ _01531_ _08181_ vssd1 vssd1 vccd1 vccd1 _01532_ sky130_fd_sc_hd__o2111a_1
XTAP_TAPCELL_ROW_19_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16600_ obsg2.obstacleArray\[84\] net447 vssd1 vssd1 vccd1 vccd1 _02279_ sky130_fd_sc_hd__or2_1
XFILLER_0_138_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13812_ control.divider.fsm.current_mode\[0\] net1649 _08109_ vssd1 vssd1 vccd1 vccd1
+ _00080_ sky130_fd_sc_hd__mux2_1
X_17580_ ag2.body\[343\] net935 vssd1 vssd1 vccd1 vccd1 _03259_ sky130_fd_sc_hd__or2_1
XANTENNA__14020__X _08181_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13454__A1 net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09658__B1 _04618_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14792_ net974 _04201_ _04202_ net1025 _01462_ vssd1 vssd1 vccd1 vccd1 _01463_ sky130_fd_sc_hd__a221o_1
XFILLER_0_86_904 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__20340__RESET_B net1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16531_ net433 _02205_ vssd1 vssd1 vccd1 vccd1 _02210_ sky130_fd_sc_hd__and2_1
X_10955_ ag2.body\[172\] net1127 vssd1 vssd1 vccd1 vccd1 _05928_ sky130_fd_sc_hd__or2_1
X_13743_ _08061_ _08062_ _08063_ vssd1 vssd1 vccd1 vccd1 _08064_ sky130_fd_sc_hd__and3_1
XANTENNA__12188__A net1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19250_ clknet_leaf_75_clk _00194_ net1492 vssd1 vssd1 vccd1 vccd1 ag2.body\[113\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_54_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_516 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16462_ obsg2.obstacleArray\[48\] obsg2.obstacleArray\[49\] net454 vssd1 vssd1 vccd1
+ vccd1 _02141_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13206__A1 net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13674_ _07181_ _08021_ vssd1 vssd1 vccd1 vccd1 track.nextCurrScore\[1\] sky130_fd_sc_hd__nor2_1
X_10886_ net1094 control.body\[653\] vssd1 vssd1 vccd1 vccd1 _05859_ sky130_fd_sc_hd__xor2_1
XFILLER_0_39_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18201_ obsg2.obstacleArray\[97\] _03739_ net520 vssd1 vssd1 vccd1 vccd1 _01348_
+ sky130_fd_sc_hd__o21a_1
X_15413_ net2487 net81 _01597_ control.body\[629\] vssd1 vssd1 vccd1 vccd1 _00703_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_94_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12625_ net277 _07513_ _07514_ net2024 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[68\]
+ sky130_fd_sc_hd__a22o_1
X_19181_ clknet_leaf_20_clk _00125_ net1365 vssd1 vssd1 vccd1 vccd1 ag2.body\[44\]
+ sky130_fd_sc_hd__dfrtp_4
X_16393_ net401 _02071_ net366 vssd1 vssd1 vccd1 vccd1 _02072_ sky130_fd_sc_hd__o21a_1
XFILLER_0_26_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18132_ net41 vssd1 vssd1 vccd1 vccd1 _03703_ sky130_fd_sc_hd__inv_2
XANTENNA__14834__C _08378_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15344_ net2616 net71 _01590_ net2431 vssd1 vssd1 vccd1 vccd1 _00641_ sky130_fd_sc_hd__a22o_1
X_12556_ net2070 net660 _07477_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[36\]
+ sky130_fd_sc_hd__and3_1
XFILLER_0_26_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09928__C _04876_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11507_ net1054 _06478_ vssd1 vssd1 vccd1 vccd1 _06480_ sky130_fd_sc_hd__xnor2_2
X_18063_ net300 _03579_ vssd1 vssd1 vccd1 vccd1 _03658_ sky130_fd_sc_hd__nand2_1
XANTENNA__15011__B net58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10436__A net1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15275_ net2061 net88 _01583_ control.body\[745\] vssd1 vssd1 vccd1 vccd1 _00579_
+ sky130_fd_sc_hd__a22o_1
X_12487_ net1666 _07437_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[7\] sky130_fd_sc_hd__and2_1
XFILLER_0_53_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_130_4278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17014_ ag2.body\[328\] net889 vssd1 vssd1 vccd1 vccd1 _02693_ sky130_fd_sc_hd__nand2_1
Xhold109 img_gen.tracker.frame\[461\] vssd1 vssd1 vccd1 vccd1 net1671 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_130_4289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11438_ _06407_ _06408_ _06409_ _06410_ vssd1 vssd1 vccd1 vccd1 _06411_ sky130_fd_sc_hd__or4_1
X_14226_ net833 ag2.body\[393\] ag2.body\[398\] net800 vssd1 vssd1 vccd1 vccd1 _08387_
+ sky130_fd_sc_hd__o22a_1
XANTENNA__15946__B net61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1031 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14157_ net824 ag2.body\[618\] ag2.body\[622\] net798 _08317_ vssd1 vssd1 vccd1 vccd1
+ _08318_ sky130_fd_sc_hd__a221o_1
X_11369_ _06331_ _06334_ _06341_ _06327_ _06314_ vssd1 vssd1 vccd1 vccd1 _06342_ sky130_fd_sc_hd__o32a_1
XFILLER_0_46_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10723__X _05696_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13108_ img_gen.tracker.frame\[319\] net652 vssd1 vssd1 vccd1 vccd1 _07747_ sky130_fd_sc_hd__and2_1
XANTENNA__11538__Y _06511_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14088_ net1022 ag2.body\[286\] vssd1 vssd1 vccd1 vccd1 _08249_ sky130_fd_sc_hd__xor2_1
X_18965_ clknet_leaf_5_clk img_gen.tracker.next_frame\[403\] net1268 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[403\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__19207__Q ag2.body\[70\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17408__B1 net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11267__A net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17916_ _04258_ _03550_ net517 vssd1 vssd1 vccd1 vccd1 _01252_ sky130_fd_sc_hd__a21oi_1
X_13039_ net233 _07713_ _07714_ net1999 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[282\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_28_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10171__A _05133_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18896_ clknet_leaf_12_clk img_gen.tracker.next_frame\[334\] net1285 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[334\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_101_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__20428__RESET_B net1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1160 net1161 vssd1 vssd1 vccd1 vccd1 net1160 sky130_fd_sc_hd__buf_2
XFILLER_0_94_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1171 net1172 vssd1 vssd1 vccd1 vccd1 net1171 sky130_fd_sc_hd__buf_4
X_17847_ img_gen.updater.commands.rR1.rainbowRNG\[9\] img_gen.updater.commands.rR1.rainbowRNG\[8\]
+ img_gen.updater.commands.rR1.rainbowRNG\[7\] _03501_ vssd1 vssd1 vccd1 vccd1 _03503_
+ sky130_fd_sc_hd__and4_1
Xfanout1182 net1183 vssd1 vssd1 vccd1 vccd1 net1182 sky130_fd_sc_hd__buf_4
XANTENNA__16269__S net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1193 net1194 vssd1 vssd1 vccd1 vccd1 net1193 sky130_fd_sc_hd__buf_4
XANTENNA__16092__C1 net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17778_ _01819_ _01887_ _02051_ _03456_ vssd1 vssd1 vccd1 vccd1 _03457_ sky130_fd_sc_hd__a211oi_4
XANTENNA__12369__Y _07335_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10259__A1 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19517_ clknet_leaf_121_clk _00461_ net1402 vssd1 vssd1 vccd1 vccd1 control.body\[875\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_135_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16729_ obsg2.obstacleArray\[113\] net482 _02407_ net499 vssd1 vssd1 vccd1 vccd1
+ _02408_ sky130_fd_sc_hd__a211o_1
XANTENNA__10259__B2 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_425 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1155 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19448_ clknet_leaf_109_clk _00392_ net1420 vssd1 vssd1 vccd1 vccd1 control.body\[950\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_76_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_100_3370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09201_ ag2.body\[623\] vssd1 vssd1 vccd1 vccd1 _04226_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_100_3381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_406 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19379_ clknet_leaf_112_clk _00323_ net1426 vssd1 vssd1 vccd1 vccd1 control.body\[1009\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__17401__B net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18136__A1 _03542_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09132_ ag2.body\[443\] vssd1 vssd1 vccd1 vccd1 _04157_ sky130_fd_sc_hd__inv_2
XFILLER_0_72_631 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_582 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10431__A1 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09063_ ag2.body\[259\] vssd1 vssd1 vccd1 vccd1 _04088_ sky130_fd_sc_hd__inv_2
XFILLER_0_72_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout213_A net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_3764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold610 sound_gen.osc1.stayCount\[4\] vssd1 vssd1 vccd1 vccd1 net2172 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__15856__B net59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11606__S1 net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_3775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold621 control.body\[1067\] vssd1 vssd1 vccd1 vccd1 net2183 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18232__B net41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold632 control.body\[910\] vssd1 vssd1 vccd1 vccd1 net2194 sky130_fd_sc_hd__dlygate4sd3_1
X_20223_ clknet_leaf_61_clk _01167_ net1469 vssd1 vssd1 vccd1 vccd1 ag2.body\[173\]
+ sky130_fd_sc_hd__dfrtp_4
Xhold643 control.body\[1070\] vssd1 vssd1 vccd1 vccd1 net2205 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13920__A2 net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold654 control.body\[789\] vssd1 vssd1 vccd1 vccd1 net2216 sky130_fd_sc_hd__dlygate4sd3_1
Xhold665 _00676_ vssd1 vssd1 vccd1 vccd1 net2227 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1122_A ag2.x\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold676 control.body\[759\] vssd1 vssd1 vccd1 vccd1 net2238 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11931__A1 net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10734__A2 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold687 control.body\[874\] vssd1 vssd1 vccd1 vccd1 net2249 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__19264__RESET_B net1504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold698 control.body\[1032\] vssd1 vssd1 vccd1 vccd1 net2260 sky130_fd_sc_hd__dlygate4sd3_1
X_20154_ clknet_leaf_94_clk _01098_ net1439 vssd1 vssd1 vccd1 vccd1 ag2.body\[232\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_60_1159 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09965_ ag2.body\[85\] net1117 vssd1 vssd1 vccd1 vccd1 _04938_ sky130_fd_sc_hd__xor2_1
XANTENNA_fanout582_A net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10081__A net1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20085_ clknet_leaf_77_clk _01029_ net1491 vssd1 vssd1 vccd1 vccd1 ag2.body\[307\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__20337__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09896_ ag2.body\[78\] net1088 vssd1 vssd1 vccd1 vccd1 _04869_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout1008_X net1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout370_X net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14488__A net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1491_A net1492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_3579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout468_X net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13392__A net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__20487__CLK clknet_leaf_37_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11542__S0 net1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1377_X net1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11998__A1 net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10740_ ag2.body\[502\] net1089 vssd1 vssd1 vccd1 vccd1 _05713_ sky130_fd_sc_hd__nand2_1
XFILLER_0_67_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17949__D net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_929 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_2786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_2797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout802_X net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10671_ _04418_ _04984_ _05632_ _05634_ _05643_ vssd1 vssd1 vccd1 vccd1 _05644_ sky130_fd_sc_hd__o32a_1
XANTENNA__10808__X _05781_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12410_ net1118 _06721_ _07372_ _06625_ vssd1 vssd1 vccd1 vccd1 _07373_ sky130_fd_sc_hd__a31o_1
XANTENNA__18126__C net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13390_ net251 _07868_ _07869_ net1800 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[478\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_10_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12411__A2 _06505_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09812__B1 net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12341_ _06821_ _07307_ vssd1 vssd1 vccd1 vccd1 _07308_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10256__A net1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17965__C net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15060_ net2663 net149 _01559_ control.body\[938\] vssd1 vssd1 vccd1 vccd1 _00388_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_133_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12272_ _07200_ _07241_ _07231_ img_gen.updater.commands.cmd_num\[3\] vssd1 vssd1
+ vccd1 vccd1 _07242_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_65_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14011_ net989 ag2.body\[457\] vssd1 vssd1 vccd1 vccd1 _08172_ sky130_fd_sc_hd__xor2_1
XANTENNA__11639__X _06612_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11223_ net1130 control.body\[860\] vssd1 vssd1 vccd1 vccd1 _06196_ sky130_fd_sc_hd__or2_1
XFILLER_0_82_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09764__B net1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12471__A _06724_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12902__C net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11922__B2 net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1514 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11154_ ag2.body\[605\] net1097 vssd1 vssd1 vccd1 vccd1 _06127_ sky130_fd_sc_hd__or2_1
XFILLER_0_101_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18727__CLK clknet_leaf_144_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10105_ net1107 control.body\[941\] vssd1 vssd1 vccd1 vccd1 _05078_ sky130_fd_sc_hd__nand2_1
X_18750_ clknet_leaf_143_clk img_gen.tracker.next_frame\[188\] net1255 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[188\] sky130_fd_sc_hd__dfrtp_1
X_15962_ ag2.body\[150\] net198 _01657_ ag2.body\[142\] vssd1 vssd1 vccd1 vccd1 _01192_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_41_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11085_ ag2.body\[537\] net1203 vssd1 vssd1 vccd1 vccd1 _06058_ sky130_fd_sc_hd__xor2_1
X_17701_ net420 _03377_ _03379_ _01911_ vssd1 vssd1 vccd1 vccd1 _03380_ sky130_fd_sc_hd__o211a_1
XANTENNA__09780__A net1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10036_ ag2.body\[504\] net788 _05005_ _05006_ _05004_ vssd1 vssd1 vccd1 vccd1 _05009_
+ sky130_fd_sc_hd__a221o_1
X_14913_ net2553 net171 _01542_ control.body\[1064\] vssd1 vssd1 vccd1 vccd1 _00258_
+ sky130_fd_sc_hd__a22o_1
X_18681_ clknet_leaf_27_clk img_gen.tracker.next_frame\[119\] net1340 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[119\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__10930__A1_N net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_4060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16089__S net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15893_ ag2.body\[200\] net133 _01650_ ag2.body\[192\] vssd1 vssd1 vccd1 vccd1 _01130_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_56_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_123_4071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17632_ ag2.body\[161\] net733 net941 _04051_ _03310_ vssd1 vssd1 vccd1 vccd1 _03311_
+ sky130_fd_sc_hd__a221o_1
X_14844_ _08705_ _08712_ _08783_ _01489_ _01499_ vssd1 vssd1 vccd1 vccd1 _01515_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_54_1420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17563_ ag2.body\[581\] net950 vssd1 vssd1 vccd1 vccd1 _03242_ sky130_fd_sc_hd__nand2_1
XFILLER_0_58_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14775_ net1038 ag2.body\[276\] vssd1 vssd1 vccd1 vccd1 _01446_ sky130_fd_sc_hd__xor2_1
XFILLER_0_114_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11987_ img_gen.tracker.frame\[397\] net616 net571 vssd1 vssd1 vccd1 vccd1 _06959_
+ sky130_fd_sc_hd__o21a_1
X_19302_ clknet_leaf_99_clk _00246_ net1448 vssd1 vssd1 vccd1 vccd1 control.body\[1092\]
+ sky130_fd_sc_hd__dfrtp_1
X_16514_ _02182_ _02183_ net402 vssd1 vssd1 vccd1 vccd1 _02193_ sky130_fd_sc_hd__mux2_1
X_13726_ net2058 toggle1.nextBlinkToggle\[0\] toggle1.nextBlinkToggle\[1\] net1923
+ vssd1 vssd1 vccd1 vccd1 toggle1.nextDisplayOut\[2\] sky130_fd_sc_hd__a22o_1
X_17494_ ag2.body\[364\] net713 net706 ag2.body\[365\] _03172_ vssd1 vssd1 vccd1 vccd1
+ _03173_ sky130_fd_sc_hd__o221a_1
XFILLER_0_105_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10938_ ag2.body\[297\] net1210 vssd1 vssd1 vccd1 vccd1 _05911_ sky130_fd_sc_hd__xor2_1
XFILLER_0_15_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19233_ clknet_leaf_84_clk _00177_ net1481 vssd1 vssd1 vccd1 vccd1 ag2.body\[96\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__17221__B net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16445_ obsg2.obstacleArray\[70\] net456 vssd1 vssd1 vccd1 vccd1 _02124_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_136_4465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13657_ _08011_ _08012_ vssd1 vssd1 vccd1 vccd1 control.divider.next_count\[19\]
+ sky130_fd_sc_hd__nor2_1
X_10869_ ag2.body\[534\] net1084 vssd1 vssd1 vccd1 vccd1 _05842_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_136_4476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12646__A net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11550__A net1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16129__B1 net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19164_ clknet_leaf_52_clk _00108_ net1368 vssd1 vssd1 vccd1 vccd1 ag2.body\[27\]
+ sky130_fd_sc_hd__dfrtp_4
X_12608_ net333 _07444_ _07505_ vssd1 vssd1 vccd1 vccd1 _07506_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_45_1693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16376_ net433 _02053_ _02054_ vssd1 vssd1 vccd1 vccd1 _02055_ sky130_fd_sc_hd__and3_1
XFILLER_0_13_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13588_ control.divider.count\[6\] _07949_ _07956_ _07962_ vssd1 vssd1 vccd1 vccd1
+ _07963_ sky130_fd_sc_hd__a22o_1
X_18115_ obsg2.obstacleArray\[58\] _03692_ net525 vssd1 vssd1 vccd1 vccd1 _01309_
+ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_41_1568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_472 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15327_ net2607 net74 _01589_ control.body\[711\] vssd1 vssd1 vccd1 vccd1 _00625_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_41_1579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19095_ clknet_leaf_146_clk img_gen.tracker.next_frame\[533\] net1239 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[533\] sky130_fd_sc_hd__dfrtp_1
X_12539_ net439 net469 net572 net546 vssd1 vssd1 vccd1 vccd1 _07467_ sky130_fd_sc_hd__or4_1
XFILLER_0_129_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18046_ net301 _03558_ vssd1 vssd1 vccd1 vccd1 _03647_ sky130_fd_sc_hd__nand2_1
XANTENNA__19502__CLK clknet_leaf_115_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15258_ net2103 net109 net50 control.body\[764\] vssd1 vssd1 vccd1 vccd1 _00566_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_41_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14209_ net1037 ag2.body\[412\] vssd1 vssd1 vccd1 vccd1 _08370_ sky130_fd_sc_hd__xor2_1
XANTENNA__17629__B1 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09674__B _04646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_3093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15189_ net2608 net101 _01572_ net2251 vssd1 vssd1 vccd1 vccd1 _00504_ sky130_fd_sc_hd__a22o_1
XANTENNA__17724__S0 net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20371__Q obsg2.obstacleArray\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout408 _01902_ vssd1 vssd1 vccd1 vccd1 net408 sky130_fd_sc_hd__buf_2
XFILLER_0_22_1419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19997_ clknet_leaf_66_clk _00941_ net1475 vssd1 vssd1 vccd1 vccd1 ag2.body\[395\]
+ sky130_fd_sc_hd__dfrtp_4
Xfanout419 _01898_ vssd1 vssd1 vccd1 vccd1 net419 sky130_fd_sc_hd__buf_4
XANTENNA__15655__A2 net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09750_ _04712_ _04713_ _04719_ _04722_ vssd1 vssd1 vccd1 vccd1 _04723_ sky130_fd_sc_hd__or4_2
XANTENNA__13666__A1 net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18948_ clknet_leaf_5_clk img_gen.tracker.next_frame\[386\] net1277 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[386\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__09690__A ag2.body\[68\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09681_ _03979_ net1078 net744 ag2.body\[15\] vssd1 vssd1 vccd1 vccd1 _04654_ sky130_fd_sc_hd__a22o_1
X_18879_ clknet_leaf_12_clk img_gen.tracker.next_frame\[317\] net1281 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[317\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_55_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14101__A net1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13418__A1 net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_102_3421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_3432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_1407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_102_3443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16907__A2 net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout37 _03705_ vssd1 vssd1 vccd1 vccd1 net37 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_58_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout48 _03534_ vssd1 vssd1 vccd1 vccd1 net48 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_119_3940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout330_A net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout59 net62 vssd1 vssd1 vccd1 vccd1 net59 sky130_fd_sc_hd__buf_8
XFILLER_0_130_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16028__A net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout428_A net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_119_3951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1072_A net1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_119_3962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_115_3826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09115_ ag2.body\[387\] vssd1 vssd1 vccd1 vccd1 _04140_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_115_3837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_1302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_70_Left_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_21_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16462__S net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1337_A net1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_645 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19182__CLK clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09046_ ag2.body\[230\] vssd1 vssd1 vccd1 vccd1 _04071_ sky130_fd_sc_hd__inv_2
XFILLER_0_5_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16034__Y _01713_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13387__A _07546_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15894__A2 net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold440 img_gen.tracker.frame\[539\] vssd1 vssd1 vccd1 vccd1 net2002 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_83_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13818__C _08113_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1504_A net1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1125_X net1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold451 img_gen.tracker.frame\[31\] vssd1 vssd1 vccd1 vccd1 net2013 sky130_fd_sc_hd__dlygate4sd3_1
Xhold462 img_gen.tracker.frame\[68\] vssd1 vssd1 vccd1 vccd1 net2024 sky130_fd_sc_hd__dlygate4sd3_1
X_20206_ clknet_leaf_56_clk _01150_ net1456 vssd1 vssd1 vccd1 vccd1 ag2.body\[188\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_74_2590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold473 img_gen.tracker.frame\[250\] vssd1 vssd1 vccd1 vccd1 net2035 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09573__A2 net1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold484 img_gen.tracker.frame\[199\] vssd1 vssd1 vccd1 vccd1 net2046 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11619__B net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold495 img_gen.tracker.frame\[144\] vssd1 vssd1 vccd1 vccd1 net2057 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_70_2443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout964_A net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout585_X net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_2454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout920 control.body_update.curr_length\[1\] vssd1 vssd1 vccd1 vccd1 net920 sky130_fd_sc_hd__clkbuf_4
XANTENNA__15646__A2 net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout931 obsg2.randCord\[7\] vssd1 vssd1 vccd1 vccd1 net931 sky130_fd_sc_hd__buf_4
XANTENNA__11380__A2 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_2465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20137_ clknet_leaf_96_clk _01081_ net1449 vssd1 vssd1 vccd1 vccd1 ag2.body\[263\]
+ sky130_fd_sc_hd__dfrtp_4
Xfanout942 net943 vssd1 vssd1 vccd1 vccd1 net942 sky130_fd_sc_hd__buf_4
X_09948_ net1097 control.body\[741\] vssd1 vssd1 vccd1 vccd1 _04921_ sky130_fd_sc_hd__xor2_1
Xfanout953 net955 vssd1 vssd1 vccd1 vccd1 net953 sky130_fd_sc_hd__buf_4
XFILLER_0_99_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14854__B1 _08862_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout964 net967 vssd1 vssd1 vccd1 vccd1 net964 sky130_fd_sc_hd__buf_4
Xfanout975 net976 vssd1 vssd1 vccd1 vccd1 net975 sky130_fd_sc_hd__buf_4
XANTENNA__18045__B1 net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout986 ag2.randCord\[2\] vssd1 vssd1 vccd1 vccd1 net986 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_5_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17306__B net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20068_ clknet_leaf_73_clk _01012_ net1500 vssd1 vssd1 vccd1 vccd1 ag2.body\[322\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_137_1318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09879_ ag2.body\[166\] net1081 vssd1 vssd1 vccd1 vccd1 _04852_ sky130_fd_sc_hd__nand2_1
Xfanout997 net1005 vssd1 vssd1 vccd1 vccd1 net997 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_5_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout752_X net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17399__A2 net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_2962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11910_ img_gen.tracker.frame\[382\] net588 net575 _06881_ vssd1 vssd1 vccd1 vccd1
+ _06882_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_87_2973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13409__A1 net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14011__A net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_2984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12890_ net292 _07643_ _07644_ net1841 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[203\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12880__A2 _07425_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1620 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_2383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_2848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11841_ img_gen.tracker.frame\[482\] net616 net601 img_gen.tracker.frame\[485\] vssd1
+ vssd1 vccd1 vccd1 _06813_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_68_2394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_2859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14082__A1 net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14082__B2 net1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_734 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14560_ net809 ag2.body\[69\] _04002_ net1013 _08720_ vssd1 vssd1 vccd1 vccd1 _08721_
+ sky130_fd_sc_hd__a221o_1
X_11772_ img_gen.tracker.frame\[74\] net625 net608 img_gen.tracker.frame\[77\] vssd1
+ vssd1 vccd1 vccd1 _06744_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_64_2269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08944__A net1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13511_ net1768 _07916_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[552\]
+ sky130_fd_sc_hd__and2_1
X_10723_ _05686_ _05693_ _05695_ _05684_ _05671_ vssd1 vssd1 vccd1 vccd1 _05696_ sky130_fd_sc_hd__o32a_2
XFILLER_0_71_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11840__B1 net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14491_ net977 _04122_ ag2.body\[350\] net802 _08651_ vssd1 vssd1 vccd1 vccd1 _08652_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_82_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09759__B net1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12466__A net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_109_Left_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11370__A _06267_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16230_ obsg2.obstacleArray\[38\] obsg2.obstacleArray\[39\] net405 vssd1 vssd1 vccd1
+ vccd1 _01909_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10654_ ag2.body\[284\] net1140 vssd1 vssd1 vccd1 vccd1 _05627_ sky130_fd_sc_hd__xor2_1
X_13442_ net235 _07888_ _07889_ net1644 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[510\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__16880__B net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16161_ _01838_ _01839_ net374 vssd1 vssd1 vccd1 vccd1 _01840_ sky130_fd_sc_hd__mux2_1
X_13373_ net670 _07862_ vssd1 vssd1 vccd1 vccd1 _07863_ sky130_fd_sc_hd__nor2_1
X_10585_ _05532_ _05542_ _05544_ _05557_ vssd1 vssd1 vccd1 vccd1 _05558_ sky130_fd_sc_hd__o22a_1
XFILLER_0_134_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18153__A net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload18 clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 clkload18/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_126_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkload29 clknet_leaf_134_clk vssd1 vssd1 vccd1 vccd1 clkload29/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_134_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__20502__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15112_ control.body\[897\] net146 _01554_ control.body\[889\] vssd1 vssd1 vccd1
+ vccd1 _00435_ sky130_fd_sc_hd__a22o_1
X_12324_ _07251_ _07290_ vssd1 vssd1 vccd1 vccd1 _07291_ sky130_fd_sc_hd__nand2_1
X_16092_ net373 _01768_ _01770_ net346 vssd1 vssd1 vccd1 vccd1 _01771_ sky130_fd_sc_hd__a211o_1
XFILLER_0_133_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17992__A net38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09494__B net1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19920_ clknet_leaf_53_clk _00864_ net1368 vssd1 vssd1 vccd1 vccd1 ag2.body\[478\]
+ sky130_fd_sc_hd__dfrtp_4
X_15043_ control.body\[963\] net163 _01556_ net2459 vssd1 vssd1 vccd1 vccd1 _00373_
+ sky130_fd_sc_hd__a22o_1
X_12255_ img_gen.updater.commands.cmd_num\[4\] img_gen.updater.commands.cmd_num\[3\]
+ vssd1 vssd1 vccd1 vccd1 _07225_ sky130_fd_sc_hd__and2b_1
XFILLER_0_122_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12699__A2 net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12632__C net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11206_ _06160_ _06163_ _06168_ _06178_ vssd1 vssd1 vccd1 vccd1 _06179_ sky130_fd_sc_hd__o22a_1
X_19851_ clknet_leaf_93_clk _00795_ net1412 vssd1 vssd1 vccd1 vccd1 ag2.body\[537\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_102_780 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12186_ net1152 ag2.apple_cord\[3\] vssd1 vssd1 vccd1 vccd1 _07158_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_118_Left_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_125_4122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18802_ clknet_leaf_3_clk img_gen.tracker.next_frame\[240\] net1260 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[240\] sky130_fd_sc_hd__dfrtp_1
X_11137_ net642 _04420_ _04428_ _04470_ vssd1 vssd1 vccd1 vccd1 _06110_ sky130_fd_sc_hd__or4_2
XTAP_TAPCELL_ROW_125_4133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19782_ clknet_leaf_127_clk _00726_ net1331 vssd1 vssd1 vccd1 vccd1 ag2.body\[612\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_53_1951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16994_ _02666_ _02667_ _02670_ _02672_ vssd1 vssd1 vccd1 vccd1 _02673_ sky130_fd_sc_hd__a211o_1
XFILLER_0_78_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_1350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_121_4008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18733_ clknet_leaf_143_clk img_gen.tracker.next_frame\[171\] net1257 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[171\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_34_1372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15945_ ag2.body\[167\] net195 _01653_ ag2.body\[159\] vssd1 vssd1 vccd1 vccd1 _01177_
+ sky130_fd_sc_hd__a22o_1
X_11068_ _04981_ _05346_ _04434_ vssd1 vssd1 vccd1 vccd1 _06041_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_121_4019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10019_ ag2.body\[269\] net1115 vssd1 vssd1 vccd1 vccd1 _04992_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_30_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18664_ clknet_leaf_11_clk img_gen.tracker.next_frame\[102\] net1281 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[102\] sky130_fd_sc_hd__dfrtp_1
X_15876_ ag2.body\[217\] net188 _01648_ ag2.body\[209\] vssd1 vssd1 vccd1 vccd1 _01115_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_133_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17615_ ag2.body\[601\] net868 vssd1 vssd1 vccd1 vccd1 _03294_ sky130_fd_sc_hd__xor2_1
X_14827_ _01496_ _01497_ vssd1 vssd1 vccd1 vccd1 _01498_ sky130_fd_sc_hd__nand2_1
XANTENNA__19055__CLK clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18595_ clknet_leaf_13_clk img_gen.tracker.next_frame\[33\] net1282 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[33\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_118_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_138_4527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17546_ ag2.body\[321\] net876 vssd1 vssd1 vccd1 vccd1 _03225_ sky130_fd_sc_hd__or2_1
XFILLER_0_86_542 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_1744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12084__B1 net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_138_4549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14758_ net1026 ag2.body\[45\] vssd1 vssd1 vccd1 vccd1 _08919_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_127_Left_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_47_1755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_1766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20032__CLK clknet_leaf_66_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13709_ track.highScore\[7\] _08035_ _08049_ _04402_ vssd1 vssd1 vccd1 vccd1 _08050_
+ sky130_fd_sc_hd__a211oi_2
XTAP_TAPCELL_ROW_28_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17477_ ag2.body\[130\] net728 net720 ag2.body\[131\] _03155_ vssd1 vssd1 vccd1 vccd1
+ _03156_ sky130_fd_sc_hd__o221a_1
XANTENNA__11831__B1 net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09669__B _04640_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14689_ net1002 _04016_ ag2.body\[90\] net828 _08844_ vssd1 vssd1 vccd1 vccd1 _08850_
+ sky130_fd_sc_hd__o221a_1
XANTENNA__15022__B1 _01555_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19216_ clknet_leaf_57_clk _00160_ net1462 vssd1 vssd1 vccd1 vccd1 ag2.body\[79\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_15_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_940 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16428_ _02105_ _02106_ vssd1 vssd1 vccd1 vccd1 _02107_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_15_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_15_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16770__B1 net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1600 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_3280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19147_ clknet_leaf_51_clk _00091_ net1377 vssd1 vssd1 vccd1 vccd1 ag2.body\[11\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_97_3291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12526__D net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16282__S net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16359_ net369 _02037_ _02034_ _01911_ vssd1 vssd1 vccd1 vccd1 _02038_ sky130_fd_sc_hd__o211a_1
XFILLER_0_15_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18063__A net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17314__A2 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11595__C1 net1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_93_3155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_3166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19078_ clknet_leaf_29_clk img_gen.tracker.next_frame\[516\] net1334 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[516\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_112_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13919__B net61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12823__B net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12139__A1 net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18029_ net351 _03635_ vssd1 vssd1 vccd1 vccd1 _03636_ sky130_fd_sc_hd__nand2_1
XFILLER_0_26_1330 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_136_Left_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11898__B1 net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout205 net210 vssd1 vssd1 vccd1 vccd1 net205 sky130_fd_sc_hd__buf_2
Xfanout216 net217 vssd1 vssd1 vccd1 vccd1 net216 sky130_fd_sc_hd__buf_2
XFILLER_0_103_1542 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15628__A2 net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09802_ net1087 control.body\[966\] vssd1 vssd1 vccd1 vccd1 _04775_ sky130_fd_sc_hd__nand2_1
Xfanout227 _07336_ vssd1 vssd1 vccd1 vccd1 net227 sky130_fd_sc_hd__buf_2
XFILLER_0_61_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout238 net247 vssd1 vssd1 vccd1 vccd1 net238 sky130_fd_sc_hd__clkbuf_4
Xfanout249 net251 vssd1 vssd1 vccd1 vccd1 net249 sky130_fd_sc_hd__clkbuf_4
XANTENNA__14836__B1 _08884_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_3630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18027__B1 net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1339 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09733_ ag2.body\[88\] net1235 vssd1 vssd1 vccd1 vccd1 _04706_ sky130_fd_sc_hd__or2_1
XANTENNA__17126__B net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout280_A net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_3505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout378_A net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16589__B1 net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09664_ net918 net921 net913 vssd1 vssd1 vccd1 vccd1 _04637_ sky130_fd_sc_hd__a21o_2
XFILLER_0_96_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16965__B net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17250__B2 net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09595_ _04560_ _04561_ _04567_ _04558_ vssd1 vssd1 vccd1 vccd1 _04568_ sky130_fd_sc_hd__a211o_1
XANTENNA__14766__A net992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18238__A _03679_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15261__B1 net50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout545_A net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13670__A _04239_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1287_A net1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15800__A2 net210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12075__B1 net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19548__CLK clknet_leaf_115_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout712_A net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout333_X net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1075_X net1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15013__B1 _01553_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1454_A net1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11190__A _05921_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17796__B net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16761__B1 net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15597__A _04447_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18572__CLK clknet_leaf_15_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout500_X net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16192__S net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12573__X _07486_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_76_2630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_2641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10370_ net783 control.body\[760\] vssd1 vssd1 vccd1 vccd1 _05343_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_76_2652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17710__C1 net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_72_2505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_2051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09029_ ag2.body\[176\] vssd1 vssd1 vccd1 vccd1 _04054_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_72_2516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_2062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10534__A net1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_2073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14006__A net1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_1490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12040_ img_gen.tracker.frame\[15\] net611 net594 img_gen.tracker.frame\[21\] _07011_
+ vssd1 vssd1 vccd1 vccd1 _07012_ sky130_fd_sc_hd__a221oi_1
Xhold270 img_gen.tracker.frame\[60\] vssd1 vssd1 vccd1 vccd1 net1832 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11349__B net1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11889__B1 net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold281 img_gen.tracker.frame\[549\] vssd1 vssd1 vccd1 vccd1 net1843 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10253__B net1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout967_X net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold292 img_gen.tracker.frame\[195\] vssd1 vssd1 vccd1 vccd1 net1854 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16221__A net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout750 net751 vssd1 vssd1 vccd1 vccd1 net750 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_102_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout761 net762 vssd1 vssd1 vccd1 vccd1 net761 sky130_fd_sc_hd__clkbuf_4
XANTENNA__17036__B net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout772 _04230_ vssd1 vssd1 vccd1 vccd1 net772 sky130_fd_sc_hd__buf_4
X_13991_ _04697_ net67 vssd1 vssd1 vccd1 vccd1 _08160_ sky130_fd_sc_hd__and2_2
Xfanout783 net785 vssd1 vssd1 vccd1 vccd1 net783 sky130_fd_sc_hd__buf_4
XFILLER_0_99_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout794 net796 vssd1 vssd1 vccd1 vccd1 net794 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11365__A net1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15730_ ag2.body\[359\] net194 _01632_ ag2.body\[351\] vssd1 vssd1 vccd1 vccd1 _00985_
+ sky130_fd_sc_hd__a22o_1
X_12942_ net246 _07667_ _07668_ net1881 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[231\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_87_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20055__CLK clknet_leaf_73_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10864__A1 _05813_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15661_ ag2.body\[409\] net142 _01625_ ag2.body\[401\] vssd1 vssd1 vccd1 vccd1 _00923_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_119_1582 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12873_ net267 _07636_ _07637_ net1616 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[193\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__14676__A net1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17400_ _03071_ _03073_ _03077_ _03078_ vssd1 vssd1 vccd1 vccd1 _03079_ sky130_fd_sc_hd__or4_1
X_14612_ _08770_ _08772_ vssd1 vssd1 vccd1 vccd1 _08773_ sky130_fd_sc_hd__nand2_1
XFILLER_0_115_1446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18380_ _03800_ _03869_ _08051_ vssd1 vssd1 vccd1 vccd1 _03870_ sky130_fd_sc_hd__a21o_1
X_11824_ img_gen.tracker.frame\[419\] net584 net560 _06795_ vssd1 vssd1 vccd1 vccd1
+ _06796_ sky130_fd_sc_hd__o211a_1
XFILLER_0_115_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15592_ ag2.body\[475\] net131 _01618_ ag2.body\[467\] vssd1 vssd1 vccd1 vccd1 _00861_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_90_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17331_ net924 net696 vssd1 vssd1 vccd1 vccd1 _03010_ sky130_fd_sc_hd__nor2_1
X_14543_ net991 ag2.body\[241\] vssd1 vssd1 vccd1 vccd1 _08704_ sky130_fd_sc_hd__xor2_1
XFILLER_0_68_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09489__B net1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11755_ img_gen.tracker.frame\[248\] net542 _06725_ _06726_ vssd1 vssd1 vccd1 vccd1
+ _06727_ sky130_fd_sc_hd__o211a_1
XANTENNA__15004__B1 _01552_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12627__C net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10706_ ag2.body\[18\] net1175 vssd1 vssd1 vccd1 vccd1 _05679_ sky130_fd_sc_hd__xor2_1
X_17262_ ag2.body\[255\] net936 vssd1 vssd1 vccd1 vccd1 _02941_ sky130_fd_sc_hd__xor2_1
X_14474_ _08631_ _08632_ _08634_ vssd1 vssd1 vccd1 vccd1 _08635_ sky130_fd_sc_hd__or3_1
XFILLER_0_125_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16752__B1 net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11686_ net1095 net1070 net743 vssd1 vssd1 vccd1 vccd1 _06658_ sky130_fd_sc_hd__and3_1
X_19001_ clknet_leaf_2_clk img_gen.tracker.next_frame\[439\] net1247 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[439\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_71_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16213_ net433 _01891_ vssd1 vssd1 vccd1 vccd1 _01892_ sky130_fd_sc_hd__and2_1
XANTENNA__12346__D net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13425_ _07567_ net302 vssd1 vssd1 vccd1 vccd1 _07882_ sky130_fd_sc_hd__or2_1
XFILLER_0_10_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10637_ _05606_ _05607_ _05608_ _05609_ _05605_ vssd1 vssd1 vccd1 vccd1 _05610_ sky130_fd_sc_hd__a221o_1
XFILLER_0_36_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17193_ _02862_ _02863_ _02870_ _02871_ vssd1 vssd1 vccd1 vccd1 _02872_ sky130_fd_sc_hd__a22o_1
Xclkload107 clknet_leaf_57_clk vssd1 vssd1 vccd1 vccd1 clkload107/Y sky130_fd_sc_hd__inv_6
XANTENNA__12924__A net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload118 clknet_leaf_65_clk vssd1 vssd1 vccd1 vccd1 clkload118/Y sky130_fd_sc_hd__clkinv_8
Xclkload129 clknet_leaf_70_clk vssd1 vssd1 vccd1 vccd1 clkload129/Y sky130_fd_sc_hd__inv_4
X_16144_ net374 _01820_ _01822_ net347 vssd1 vssd1 vccd1 vccd1 _01823_ sky130_fd_sc_hd__a211o_1
XANTENNA__11041__A1 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_116_Right_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13356_ net274 _07854_ _07855_ net1772 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[458\]
+ sky130_fd_sc_hd__a22o_1
X_10568_ ag2.body\[515\] net771 net751 ag2.body\[518\] vssd1 vssd1 vccd1 vccd1 _05541_
+ sky130_fd_sc_hd__o22a_1
XANTENNA__17701__C1 _01911_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12307_ _07273_ vssd1 vssd1 vccd1 vccd1 _07274_ sky130_fd_sc_hd__inv_2
X_16075_ obsg2.obstacleArray\[127\] net430 net376 _01753_ vssd1 vssd1 vccd1 vccd1
+ _01754_ sky130_fd_sc_hd__o211a_1
XANTENNA__10444__A net1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10499_ _05467_ _05468_ _05470_ _05471_ vssd1 vssd1 vccd1 vccd1 _05472_ sky130_fd_sc_hd__and4b_1
X_13287_ net280 _07827_ _07828_ net1976 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[416\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_62_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_127_4206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19903_ clknet_leaf_86_clk _00847_ net1464 vssd1 vssd1 vccd1 vccd1 ag2.body\[493\]
+ sky130_fd_sc_hd__dfrtp_4
X_15026_ control.body\[980\] net152 _01555_ net2239 vssd1 vssd1 vccd1 vccd1 _00358_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_36_1412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12238_ _07196_ _07207_ _07206_ vssd1 vssd1 vccd1 vccd1 _07208_ sky130_fd_sc_hd__o21bai_1
XTAP_TAPCELL_ROW_36_1423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_36_1434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10163__B net1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16807__B2 ag2.body\[70\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09952__B net1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19834_ clknet_leaf_122_clk _00778_ net1414 vssd1 vssd1 vccd1 vccd1 ag2.body\[552\]
+ sky130_fd_sc_hd__dfrtp_4
X_12169_ img_gen.tracker.frame\[423\] net599 vssd1 vssd1 vccd1 vccd1 _07141_ sky130_fd_sc_hd__or2_1
XFILLER_0_23_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16977_ ag2.body\[428\] net960 vssd1 vssd1 vccd1 vccd1 _02656_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_120_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19765_ clknet_leaf_127_clk _00709_ net1326 vssd1 vssd1 vccd1 vccd1 control.body\[627\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_120_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14294__A1 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14294__B2 net1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput5 gpio_in[28] vssd1 vssd1 vccd1 vccd1 net5 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_127_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17514__X _03193_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15928_ ag2.body\[183\] net136 _01654_ ag2.body\[175\] vssd1 vssd1 vccd1 vccd1 _01161_
+ sky130_fd_sc_hd__a22o_1
X_18716_ clknet_leaf_144_clk img_gen.tracker.next_frame\[154\] net1252 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[154\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_36_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19696_ clknet_leaf_136_clk net2231 net1301 vssd1 vssd1 vccd1 vccd1 control.body\[702\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_49_1806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18647_ clknet_leaf_130_clk img_gen.tracker.next_frame\[85\] net1316 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[85\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_49_1828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15859_ ag2.body\[234\] net175 _01646_ ag2.body\[226\] vssd1 vssd1 vccd1 vccd1 _01100_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_133_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18058__A net43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15243__B1 _01578_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13490__A net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09380_ _04366_ _04374_ vssd1 vssd1 vccd1 vccd1 _01413_ sky130_fd_sc_hd__nor2_1
XANTENNA__20548__CLK clknet_leaf_105_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12057__B1 net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18578_ clknet_leaf_15_clk img_gen.tracker.next_frame\[16\] net1279 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[16\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__16991__B1 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_99_3331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18595__CLK clknet_leaf_13_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17529_ ag2.body\[277\] net951 vssd1 vssd1 vccd1 vccd1 _03208_ sky130_fd_sc_hd__or2_1
XANTENNA__11722__B net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10178__X _05151_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_3342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11804__B1 net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_3353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_3206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20540_ clknet_leaf_106_clk _01405_ _00014_ vssd1 vssd1 vccd1 vccd1 sound_gen.osc1.stayCount\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_95_3217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_3228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16743__B1 net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10338__B net1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20471_ clknet_leaf_33_clk _01358_ net1346 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[107\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__12834__A _06671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout126_A net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_83_clk_X clknet_leaf_83_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11568__C1 _06497_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09776__A2 net1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12553__B net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16740__S net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1035_A net1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_98_clk_X clknet_leaf_98_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1040 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16259__C1 _01912_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18240__B net35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout495_A net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19220__CLK clknet_leaf_75_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09862__B net1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_141_clk_X clknet_leaf_141_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1202_A net1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout662_A net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout283_X net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_21_clk_X clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10801__B net1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15482__B1 _01605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09716_ ag2.body\[244\] net765 net745 ag2.body\[247\] vssd1 vssd1 vccd1 vccd1 _04689_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_78_1570 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19370__CLK clknet_leaf_102_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_626 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18420__B1 net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout450_X net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09647_ net1196 control.body\[745\] vssd1 vssd1 vccd1 vccd1 _04620_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_65_2320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14037__A1 net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14496__A net1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14037__B2 net1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1192_X net1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout548_X net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12048__B1 net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09578_ net899 net902 net908 net892 vssd1 vssd1 vccd1 vccd1 _04551_ sky130_fd_sc_hd__a31oi_4
XANTENNA__12599__A1 net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout715_X net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17526__A2 net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10529__A net1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_342 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11540_ obsg2.obstacleArray\[98\] obsg2.obstacleArray\[99\] obsg2.obstacleArray\[102\]
+ obsg2.obstacleArray\[103\] net1123 net510 vssd1 vssd1 vccd1 vccd1 _06513_ sky130_fd_sc_hd__mux4_1
XFILLER_0_110_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16734__B1 net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_2703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_2714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11471_ ag2.body\[495\] net1064 vssd1 vssd1 vccd1 vccd1 _06444_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_59_2113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_1387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16216__A net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12744__A net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_2124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_1484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_59_2135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13210_ net241 _07794_ _07795_ net1874 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[372\]
+ sky130_fd_sc_hd__a22o_1
X_10422_ _05393_ _05394_ _05392_ vssd1 vssd1 vccd1 vccd1 _05395_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09767__A2 _04599_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14190_ _08347_ _08348_ _08349_ _08350_ vssd1 vssd1 vccd1 vccd1 _08351_ sky130_fd_sc_hd__a22o_1
XFILLER_0_60_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12771__A1 net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10353_ ag2.body\[288\] net1237 vssd1 vssd1 vccd1 vccd1 _05326_ sky130_fd_sc_hd__and2b_1
X_13141_ net667 _07762_ vssd1 vssd1 vccd1 vccd1 _07763_ sky130_fd_sc_hd__nor2_1
XFILLER_0_81_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13072_ net685 _07729_ vssd1 vssd1 vccd1 vccd1 _07730_ sky130_fd_sc_hd__nor2_1
X_10284_ ag2.body\[329\] net1211 vssd1 vssd1 vccd1 vccd1 _05257_ sky130_fd_sc_hd__nand2_1
XFILLER_0_40_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12023_ img_gen.tracker.frame\[192\] net630 net557 img_gen.tracker.frame\[198\] _06994_
+ vssd1 vssd1 vccd1 vccd1 _06995_ sky130_fd_sc_hd__a221o_1
X_16900_ ag2.body\[242\] net726 net735 ag2.body\[241\] vssd1 vssd1 vccd1 vccd1 _02579_
+ sky130_fd_sc_hd__a2bb2o_1
Xfanout1501 net1502 vssd1 vssd1 vccd1 vccd1 net1501 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_20_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09772__B net1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17880_ obsg2.obstacleCount\[1\] obsg2.obstacleCount\[0\] obsg2.obstacleCount\[2\]
+ vssd1 vssd1 vccd1 vccd1 _03520_ sky130_fd_sc_hd__a21oi_1
XANTENNA__18254__A3 net37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1512 net1514 vssd1 vssd1 vccd1 vccd1 net1512 sky130_fd_sc_hd__clkbuf_2
XANTENNA__16265__A2 net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16831_ _02504_ _02505_ _02507_ _02509_ vssd1 vssd1 vccd1 vccd1 _02510_ sky130_fd_sc_hd__or4b_1
Xfanout580 net582 vssd1 vssd1 vccd1 vccd1 net580 sky130_fd_sc_hd__clkbuf_4
XANTENNA__16670__C1 net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19550_ clknet_leaf_115_clk _00494_ net1388 vssd1 vssd1 vccd1 vccd1 control.body\[844\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout591 net592 vssd1 vssd1 vccd1 vccd1 net591 sky130_fd_sc_hd__clkbuf_4
X_16762_ _02438_ _02440_ net498 vssd1 vssd1 vccd1 vccd1 _02441_ sky130_fd_sc_hd__mux2_1
X_13974_ ag2.body\[112\] net202 _08158_ ag2.body\[104\] vssd1 vssd1 vccd1 vccd1 _00193_
+ sky130_fd_sc_hd__a22o_1
X_18501_ net1512 net1506 vssd1 vssd1 vccd1 vccd1 _00032_ sky130_fd_sc_hd__or2_1
X_15713_ ag2.body\[360\] net193 _01630_ ag2.body\[352\] vssd1 vssd1 vccd1 vccd1 _00970_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_18_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19481_ clknet_leaf_109_clk net2111 net1416 vssd1 vssd1 vccd1 vccd1 control.body\[919\]
+ sky130_fd_sc_hd__dfrtp_1
X_12925_ net244 _07659_ _07660_ net1809 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[222\]
+ sky130_fd_sc_hd__a22o_1
X_16693_ net709 net538 vssd1 vssd1 vccd1 vccd1 _02372_ sky130_fd_sc_hd__and2_1
XFILLER_0_87_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18432_ _03917_ _03920_ _03875_ vssd1 vssd1 vccd1 vccd1 _03921_ sky130_fd_sc_hd__o21ai_1
X_15644_ ag2.body\[426\] net138 _01623_ ag2.body\[418\] vssd1 vssd1 vccd1 vccd1 _00908_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_17_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12039__B1 net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12856_ net261 _07628_ _07629_ net1891 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[184\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_69_862 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12197__Y _07169_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11807_ img_gen.tracker.frame\[455\] net578 net540 img_gen.tracker.frame\[452\] _06778_
+ vssd1 vssd1 vccd1 vccd1 _06779_ sky130_fd_sc_hd__o221a_1
X_18363_ _03856_ _03857_ net434 vssd1 vssd1 vccd1 vccd1 _03858_ sky130_fd_sc_hd__a21o_1
X_15575_ ag2.body\[493\] net135 _01615_ ag2.body\[485\] vssd1 vssd1 vccd1 vccd1 _00847_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__10439__A net1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12787_ net239 _07596_ _07597_ net1678 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[147\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_84_854 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11798__C1 net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17314_ ag2.body\[392\] net738 net733 ag2.body\[393\] _02984_ vssd1 vssd1 vccd1 vccd1
+ _02993_ sky130_fd_sc_hd__o221a_1
XFILLER_0_127_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11262__A1 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14526_ net992 ag2.body\[249\] vssd1 vssd1 vccd1 vccd1 _08687_ sky130_fd_sc_hd__or2_1
XFILLER_0_113_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18294_ net325 net323 vssd1 vssd1 vccd1 vccd1 _03790_ sky130_fd_sc_hd__nand2_1
XANTENNA__11262__B2 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11738_ img_gen.tracker.frame\[41\] net607 net577 _06709_ vssd1 vssd1 vccd1 vccd1
+ _06710_ sky130_fd_sc_hd__o211a_1
XANTENNA__16725__B1 net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17245_ ag2.body\[619\] net715 net704 ag2.body\[621\] _02923_ vssd1 vssd1 vccd1 vccd1
+ _02924_ sky130_fd_sc_hd__o221a_1
XFILLER_0_127_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14457_ net842 ag2.body\[432\] ag2.body\[438\] net800 vssd1 vssd1 vccd1 vccd1 _08618_
+ sky130_fd_sc_hd__o22a_1
XANTENNA__14200__A1 net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12654__A net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11669_ _06639_ _06640_ _06637_ vssd1 vssd1 vccd1 vccd1 _06641_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_126_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14200__B2 net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15030__A _04772_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13408_ net255 _07874_ _07875_ net1878 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[490\]
+ sky130_fd_sc_hd__a22o_1
X_17176_ ag2.body\[463\] net930 vssd1 vssd1 vccd1 vccd1 _02855_ sky130_fd_sc_hd__or2_1
X_14388_ _08547_ _08548_ vssd1 vssd1 vccd1 vccd1 _08549_ sky130_fd_sc_hd__or2_1
XFILLER_0_12_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_773 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20035__RESET_B net1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16489__C1 net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19243__CLK clknet_leaf_75_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11565__A2 net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16127_ net378 _01805_ _01804_ net348 vssd1 vssd1 vccd1 vccd1 _01806_ sky130_fd_sc_hd__a211o_1
XFILLER_0_24_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13339_ net228 _07848_ _07849_ net2047 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[447\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_110_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16560__S net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_672 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16058_ net956 net538 vssd1 vssd1 vccd1 vccd1 _01737_ sky130_fd_sc_hd__or2_2
XFILLER_0_62_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18060__B _03577_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15009_ control.body\[998\] net153 _01552_ control.body\[990\] vssd1 vssd1 vccd1
+ vccd1 _00344_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_88_3010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_3021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19393__CLK clknet_leaf_102_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19817_ clknet_leaf_124_clk _00761_ net1405 vssd1 vssd1 vccd1 vccd1 ag2.body\[583\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_23_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11717__B net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16796__A net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10621__B net1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15464__B1 _01603_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__20370__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19748_ clknet_leaf_129_clk _00692_ net1325 vssd1 vssd1 vccd1 vccd1 control.body\[642\]
+ sky130_fd_sc_hd__dfrtp_1
X_09501_ ag2.body\[402\] net1185 vssd1 vssd1 vccd1 vccd1 _04474_ sky130_fd_sc_hd__or2_1
XANTENNA__19971__RESET_B net1470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14019__A1 net999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17404__B net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14019__B2 net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19679_ clknet_leaf_135_clk _00623_ net1301 vssd1 vssd1 vccd1 vccd1 control.body\[717\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12829__A _07431_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09432_ ag2.body\[2\] net1178 vssd1 vssd1 vccd1 vccd1 _04405_ sky130_fd_sc_hd__xor2_1
XANTENNA__19900__RESET_B net1464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12548__B _07472_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09203__A net1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09363_ sound_gen.osc1.stayCount\[13\] sound_gen.osc1.stayCount\[12\] _04364_ vssd1
+ vssd1 vccd1 vccd1 _04365_ sky130_fd_sc_hd__and3_1
XANTENNA__16735__S net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13242__A2 _07807_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09294_ sound_gen.osc1.freq\[1\] sound_gen.osc1.freq\[2\] _04284_ _04285_ vssd1 vssd1
+ vccd1 vccd1 _04314_ sky130_fd_sc_hd__or4_1
XANTENNA__12450__B1 net1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16716__B1 net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_10 _03446_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_21 _08509_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_515 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_32 _03442_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20523_ clknet_leaf_93_clk track.nextCurrScore\[5\] net1413 vssd1 vssd1 vccd1 vccd1
+ control.body_update.curr_length\[5\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_28_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout410_A net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16036__A net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1152_A net1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11005__A1 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18469__B1 net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20454_ clknet_leaf_39_clk _01341_ net1356 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[90\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_28_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11005__B2 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12753__A1 net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17419__X _03098_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_63_clk_A clknet_4_13__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20385_ clknet_leaf_43_clk _01272_ net1372 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[21\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA_fanout1038_X net1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19736__CLK clknet_leaf_132_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_856 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout877_A net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout498_X net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11467__X _06440_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11908__A net1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10516__B1 net1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1205_X net1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10812__A net1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20638__1555 vssd1 vssd1 vccd1 vccd1 _20638__1555/HI net1555 sky130_fd_sc_hd__conb_1
XANTENNA_clkbuf_leaf_78_clk_A clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09921__A2 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14258__A1 net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14258__B2 net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18760__CLK clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15455__B1 _01602_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_121_clk_A clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10819__A1 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13842__B net223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10971_ net1083 control.body\[1006\] vssd1 vssd1 vccd1 vccd1 _05944_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout832_X net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12739__A net683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15207__B1 _01574_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12710_ net683 _07559_ vssd1 vssd1 vccd1 vccd1 _07560_ sky130_fd_sc_hd__nor2_1
XFILLER_0_116_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18129__C net39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19116__CLK clknet_leaf_141_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13690_ net639 _04550_ net742 vssd1 vssd1 vccd1 vccd1 _08032_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_97_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_136_clk_A clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12641_ net307 _07523_ vssd1 vssd1 vccd1 vccd1 _07524_ sky130_fd_sc_hd__nor2_1
XFILLER_0_84_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14430__A1 net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14430__B2 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15360_ control.body\[685\] net68 _01592_ net2490 vssd1 vssd1 vccd1 vccd1 _00655_
+ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_16_clk_A clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16707__B1 net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12572_ net292 _07484_ _07485_ net1850 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[44\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_108_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18172__A2 _03705_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14311_ net1034 ag2.body\[52\] vssd1 vssd1 vccd1 vccd1 _08472_ sky130_fd_sc_hd__or2_1
X_11523_ _06479_ _06482_ _06494_ vssd1 vssd1 vccd1 vccd1 _06496_ sky130_fd_sc_hd__nand3_1
XFILLER_0_4_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16183__A1 net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15291_ _04930_ net52 vssd1 vssd1 vccd1 vccd1 _01585_ sky130_fd_sc_hd__nor2_2
XFILLER_0_108_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17030_ _04144_ net855 net935 _04147_ _02704_ vssd1 vssd1 vccd1 vccd1 _02709_ sky130_fd_sc_hd__a221o_1
XANTENNA__14194__B1 ag2.body\[162\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14242_ _08397_ _08402_ vssd1 vssd1 vccd1 vccd1 _08403_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_29_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_1068 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11454_ _06399_ _06412_ _06413_ _06426_ vssd1 vssd1 vccd1 vccd1 _06427_ sky130_fd_sc_hd__o22a_1
XANTENNA__15930__B2 ag2.body\[160\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10265__Y _05238_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10706__B net1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15785__A _05909_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10405_ net1062 control.body\[1079\] vssd1 vssd1 vccd1 vccd1 _05378_ sky130_fd_sc_hd__xor2_1
X_14173_ net841 ag2.body\[192\] _04061_ net971 vssd1 vssd1 vccd1 vccd1 _08334_ sky130_fd_sc_hd__a22o_1
X_11385_ _06354_ _06355_ _06356_ _06357_ vssd1 vssd1 vccd1 vccd1 _06358_ sky130_fd_sc_hd__a22o_1
XFILLER_0_81_1235 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13124_ img_gen.tracker.frame\[328\] net663 vssd1 vssd1 vccd1 vccd1 _07754_ sky130_fd_sc_hd__and2_1
XANTENNA__09783__A net1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_480 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10336_ ag2.body\[524\] net1136 vssd1 vssd1 vccd1 vccd1 _05309_ sky130_fd_sc_hd__or2_1
X_18981_ clknet_leaf_8_clk img_gen.tracker.next_frame\[419\] net1265 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[419\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__14497__A1 net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14497__B2 net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10267_ ag2.body\[139\] net1165 vssd1 vssd1 vccd1 vccd1 _05240_ sky130_fd_sc_hd__or2_1
X_17932_ _01700_ _03531_ vssd1 vssd1 vccd1 vccd1 _03564_ sky130_fd_sc_hd__nor2_1
XFILLER_0_24_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10281__X _05254_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13055_ net246 _07720_ _07721_ net1674 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[291\]
+ sky130_fd_sc_hd__a22o_1
Xfanout1320 net1324 vssd1 vssd1 vccd1 vccd1 net1320 sky130_fd_sc_hd__buf_2
X_12006_ img_gen.tracker.frame\[469\] net616 vssd1 vssd1 vccd1 vccd1 _06978_ sky130_fd_sc_hd__or2_1
X_17863_ _04277_ _03500_ vssd1 vssd1 vccd1 vccd1 _03513_ sky130_fd_sc_hd__nand2_1
Xfanout1331 net1332 vssd1 vssd1 vccd1 vccd1 net1331 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_59_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10198_ ag2.body\[117\] net1116 vssd1 vssd1 vccd1 vccd1 _05171_ sky130_fd_sc_hd__nand2_1
XFILLER_0_20_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14249__A1 net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1342 net1344 vssd1 vssd1 vccd1 vccd1 net1342 sky130_fd_sc_hd__clkbuf_4
Xfanout1353 net1355 vssd1 vssd1 vccd1 vccd1 net1353 sky130_fd_sc_hd__clkbuf_4
XANTENNA__15446__B1 _01601_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14249__B2 net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1364 net1370 vssd1 vssd1 vccd1 vccd1 net1364 sky130_fd_sc_hd__clkbuf_4
Xfanout1375 net1377 vssd1 vssd1 vccd1 vccd1 net1375 sky130_fd_sc_hd__clkbuf_4
X_19602_ clknet_leaf_120_clk net2508 net1393 vssd1 vssd1 vccd1 vccd1 control.body\[784\]
+ sky130_fd_sc_hd__dfrtp_1
X_16814_ _04014_ net944 net694 ag2.body\[87\] vssd1 vssd1 vccd1 vccd1 _02493_ sky130_fd_sc_hd__o22a_1
X_17794_ obsmode.sOBSMODE.pb_2 obsmode.sOBSMODE.pb_1 vssd1 vssd1 vccd1 vccd1 _03468_
+ sky130_fd_sc_hd__and2b_2
Xfanout1386 net1404 vssd1 vssd1 vccd1 vccd1 net1386 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_17_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1397 net1404 vssd1 vssd1 vccd1 vccd1 net1397 sky130_fd_sc_hd__clkbuf_4
X_16745_ _02422_ _02423_ net499 vssd1 vssd1 vccd1 vccd1 _02424_ sky130_fd_sc_hd__mux2_1
X_19533_ clknet_leaf_120_clk _00477_ net1393 vssd1 vssd1 vccd1 vccd1 control.body\[859\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__17199__B1 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13957_ ag2.body\[97\] net189 _08156_ ag2.body\[89\] vssd1 vssd1 vccd1 vccd1 _00178_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12649__A net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17738__A2 _02633_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19464_ clknet_leaf_109_clk _00408_ net1416 vssd1 vssd1 vccd1 vccd1 control.body\[934\]
+ sky130_fd_sc_hd__dfrtp_1
X_12908_ net1986 net661 _07315_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[213\]
+ sky130_fd_sc_hd__and3_1
X_16676_ obsg2.obstacleArray\[27\] net451 net392 vssd1 vssd1 vccd1 vccd1 _02355_ sky130_fd_sc_hd__o21a_1
X_13888_ ag2.body\[36\] net117 _08148_ ag2.body\[28\] vssd1 vssd1 vccd1 vccd1 _00117_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_115_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10691__C1 _05237_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15627_ ag2.body\[443\] net127 _01621_ ag2.body\[435\] vssd1 vssd1 vccd1 vccd1 _00893_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11272__B net1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18415_ _04639_ _08145_ _03844_ _03904_ vssd1 vssd1 vccd1 vccd1 _03905_ sky130_fd_sc_hd__o211a_1
X_12839_ net286 _07619_ _07620_ net1660 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[176\]
+ sky130_fd_sc_hd__a22o_1
X_19395_ clknet_leaf_103_clk _00339_ net1428 vssd1 vssd1 vccd1 vccd1 control.body\[993\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_31_1613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14421__A1 net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14421__B2 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17878__C _04688_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18346_ _03840_ _03841_ _08145_ vssd1 vssd1 vccd1 vccd1 _03842_ sky130_fd_sc_hd__o21ai_1
X_15558_ ag2.body\[511\] net188 _01612_ ag2.body\[503\] vssd1 vssd1 vccd1 vccd1 _00833_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_90_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11786__A2 net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_904 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14509_ net990 _04055_ _04059_ net1008 _08666_ vssd1 vssd1 vccd1 vccd1 _08670_ sky130_fd_sc_hd__a221o_1
XFILLER_0_31_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12983__A1 net254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16174__A1 net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09677__B net1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18277_ net517 _03777_ vssd1 vssd1 vccd1 vccd1 _01386_ sky130_fd_sc_hd__nor2_1
X_15489_ ag2.body\[560\] net113 _01606_ ag2.body\[552\] vssd1 vssd1 vccd1 vccd1 _00770_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_66_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_1423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17228_ _02904_ _02906_ vssd1 vssd1 vccd1 vccd1 _02907_ sky130_fd_sc_hd__nand2_1
XANTENNA__18633__CLK clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10616__B net1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12735__A1 net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold803 control.body\[850\] vssd1 vssd1 vccd1 vccd1 net2365 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold814 _00375_ vssd1 vssd1 vccd1 vccd1 net2376 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_155 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17159_ ag2.body\[598\] net937 vssd1 vssd1 vccd1 vccd1 _02838_ sky130_fd_sc_hd__xor2_1
XANTENNA__16290__S net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold825 ag2.body\[590\] vssd1 vssd1 vccd1 vccd1 net2387 sky130_fd_sc_hd__dlygate4sd3_1
Xhold836 track.highScore\[0\] vssd1 vssd1 vccd1 vccd1 net2398 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09693__A ag2.body\[65\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold847 control.body\[934\] vssd1 vssd1 vccd1 vccd1 net2409 sky130_fd_sc_hd__dlygate4sd3_1
X_20170_ clknet_leaf_82_clk _01114_ net1479 vssd1 vssd1 vccd1 vccd1 ag2.body\[216\]
+ sky130_fd_sc_hd__dfrtp_4
Xhold858 control.body\[1046\] vssd1 vssd1 vccd1 vccd1 net2420 sky130_fd_sc_hd__dlygate4sd3_1
Xhold869 control.body\[695\] vssd1 vssd1 vccd1 vccd1 net2431 sky130_fd_sc_hd__dlygate4sd3_1
X_09981_ net1207 control.body\[1113\] vssd1 vssd1 vccd1 vccd1 _04954_ sky130_fd_sc_hd__xor2_1
XANTENNA__15685__B1 _01627_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_wire633_X net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10351__B net1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11710__A2 net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19139__CLK clknet_leaf_132_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_1248 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17134__B net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17729__A2 net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout458_A net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09204__Y _04229_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09415_ img_gen.control.current\[1\] img_gen.control.current\[0\] vssd1 vssd1 vccd1
+ vccd1 _04394_ sky130_fd_sc_hd__nand2_4
XANTENNA__19289__CLK clknet_leaf_98_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16465__S net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14412__A1 net1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout246_X net246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout625_A net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17695__A2_N net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1367_A net1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11750__X _06722_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10029__A2 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11226__A1 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09346_ sound_gen.osc1.stayCount\[21\] sound_gen.osc1.stayCount\[20\] sound_gen.osc1.stayCount\[15\]
+ sound_gen.osc1.stayCount\[13\] vssd1 vssd1 vccd1 vccd1 _04350_ sky130_fd_sc_hd__and4_1
XANTENNA__11226__B2 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18154__A2 _03582_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12974__A1 net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16165__A1 net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout413_X net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09277_ sound_gen.osc1.stayCount\[20\] _04287_ _04288_ sound_gen.osc1.stayCount\[21\]
+ vssd1 vssd1 vccd1 vccd1 _04300_ sky130_fd_sc_hd__a22o_1
XANTENNA__17901__A2 _03533_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1155_X net1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20506_ clknet_leaf_112_clk net1581 net1424 vssd1 vssd1 vccd1 vccd1 score_detect.sig_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout994_A net995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20437_ clknet_leaf_25_clk _01324_ net1343 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[73\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_107_1529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11170_ _06139_ _06140_ _06141_ _06142_ vssd1 vssd1 vccd1 vccd1 _06143_ sky130_fd_sc_hd__a22o_1
X_20368_ clknet_leaf_24_clk _01255_ net1360 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[4\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__17309__B net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout782_X net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10121_ net1046 control.body\[711\] vssd1 vssd1 vccd1 vccd1 _05094_ sky130_fd_sc_hd__nand2_1
XFILLER_0_100_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20299_ clknet_leaf_36_clk control.divider.next_count\[20\] net1351 vssd1 vssd1 vccd1
+ vccd1 control.divider.count\[20\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_105_1275 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14014__A net1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10052_ ag2.body\[485\] net1104 vssd1 vssd1 vccd1 vccd1 _05025_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_41_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14860_ _08796_ _08801_ _01530_ _08542_ vssd1 vssd1 vccd1 vccd1 _01531_ sky130_fd_sc_hd__o211a_1
XFILLER_0_76_1326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout61_X net61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08947__A net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13811_ net1649 control.divider.fsm.current_mode\[2\] _08109_ vssd1 vssd1 vccd1 vccd1
+ _00079_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17044__B net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14791_ net980 ag2.body\[546\] vssd1 vssd1 vccd1 vccd1 _01462_ sky130_fd_sc_hd__xor2_1
XFILLER_0_98_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16530_ net318 _02208_ vssd1 vssd1 vccd1 vccd1 _02209_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_93_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13742_ _04390_ _07240_ vssd1 vssd1 vccd1 vccd1 _08063_ sky130_fd_sc_hd__or2_1
XFILLER_0_54_1635 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10954_ _05923_ _05924_ _05925_ _05926_ vssd1 vssd1 vccd1 vccd1 _05927_ sky130_fd_sc_hd__or4_1
XANTENNA__16928__B1 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16461_ obsg2.obstacleArray\[50\] obsg2.obstacleArray\[51\] net454 vssd1 vssd1 vccd1
+ vccd1 _02140_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12619__D net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13673_ net919 _08020_ vssd1 vssd1 vccd1 vccd1 _08021_ sky130_fd_sc_hd__xor2_1
XFILLER_0_35_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10885_ net1220 control.body\[648\] vssd1 vssd1 vccd1 vccd1 _05858_ sky130_fd_sc_hd__xor2_1
XFILLER_0_128_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15600__B1 _01619_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18200_ _03643_ net40 vssd1 vssd1 vccd1 vccd1 _03739_ sky130_fd_sc_hd__nor2_1
XANTENNA__20380__RESET_B net1374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15412_ net2598 net81 _01597_ net2248 vssd1 vssd1 vccd1 vccd1 _00702_ sky130_fd_sc_hd__a22o_1
X_12624_ net252 _07513_ _07514_ net1876 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[67\]
+ sky130_fd_sc_hd__a22o_1
X_19180_ clknet_leaf_20_clk _00124_ net1365 vssd1 vssd1 vccd1 vccd1 ag2.body\[43\]
+ sky130_fd_sc_hd__dfrtp_4
X_16392_ obsg2.obstacleArray\[122\] obsg2.obstacleArray\[123\] net455 vssd1 vssd1
+ vccd1 vccd1 _02071_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18131_ _03531_ net296 vssd1 vssd1 vccd1 vccd1 _03702_ sky130_fd_sc_hd__or2_1
XANTENNA__11768__A2 net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12965__A1 net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17995__A net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15343_ control.body\[702\] net71 _01590_ net2230 vssd1 vssd1 vccd1 vccd1 _00640_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__16156__A1 net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12555_ net306 _07476_ vssd1 vssd1 vccd1 vccd1 _07477_ sky130_fd_sc_hd__or2_1
XFILLER_0_65_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09928__D _04900_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18062_ obsg2.obstacleArray\[40\] _03657_ net520 vssd1 vssd1 vccd1 vccd1 _01291_
+ sky130_fd_sc_hd__o21a_1
X_11506_ net1054 _06478_ vssd1 vssd1 vccd1 vccd1 _06479_ sky130_fd_sc_hd__nand2_1
XFILLER_0_41_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15274_ control.body\[752\] net88 _01583_ control.body\[744\] vssd1 vssd1 vccd1 vccd1
+ _00578_ sky130_fd_sc_hd__a22o_1
XFILLER_0_79_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12486_ net1630 _07437_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[6\] sky130_fd_sc_hd__and2_1
XFILLER_0_123_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17013_ _02685_ _02687_ _02689_ _02691_ vssd1 vssd1 vccd1 vccd1 _02692_ sky130_fd_sc_hd__or4_1
XANTENNA__12717__A1 net237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_130_4279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14225_ net843 ag2.body\[392\] ag2.body\[398\] net802 vssd1 vssd1 vccd1 vccd1 _08386_
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_124_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11437_ ag2.body\[393\] net1209 vssd1 vssd1 vccd1 vccd1 _06410_ sky130_fd_sc_hd__xor2_1
XANTENNA__17105__B1 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1190 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14156_ net970 ag2.body\[619\] vssd1 vssd1 vccd1 vccd1 _08317_ sky130_fd_sc_hd__xor2_1
X_11368_ _06328_ _06335_ _06337_ _06340_ vssd1 vssd1 vccd1 vccd1 _06341_ sky130_fd_sc_hd__or4_1
XFILLER_0_95_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11940__A2 net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13107_ net237 _07745_ _07746_ net1949 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[318\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10319_ ag2.body\[610\] net1169 vssd1 vssd1 vccd1 vccd1 _05292_ sky130_fd_sc_hd__nand2_1
X_14087_ net983 ag2.body\[282\] vssd1 vssd1 vccd1 vccd1 _08248_ sky130_fd_sc_hd__nand2_1
X_18964_ clknet_leaf_5_clk img_gen.tracker.next_frame\[402\] net1268 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[402\] sky130_fd_sc_hd__dfrtp_1
X_11299_ net1218 control.body\[680\] vssd1 vssd1 vccd1 vccd1 _06272_ sky130_fd_sc_hd__xor2_1
XANTENNA__13142__A1 net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17915_ _03549_ _03531_ _03547_ vssd1 vssd1 vccd1 vccd1 _03550_ sky130_fd_sc_hd__or3b_1
X_13038_ net673 _07713_ vssd1 vssd1 vccd1 vccd1 _07714_ sky130_fd_sc_hd__nor2_1
XANTENNA__11267__B net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_1494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18895_ clknet_leaf_12_clk img_gen.tracker.next_frame\[333\] net1285 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[333\] sky130_fd_sc_hd__dfrtp_1
Xfanout1150 net1151 vssd1 vssd1 vccd1 vccd1 net1150 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_59_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11835__X _06807_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1161 net1166 vssd1 vssd1 vccd1 vccd1 net1161 sky130_fd_sc_hd__buf_4
XFILLER_0_98_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17846_ img_gen.updater.commands.rR1.rainbowRNG\[7\] _03501_ vssd1 vssd1 vccd1 vccd1
+ _03502_ sky130_fd_sc_hd__nand2_1
Xfanout1172 net1173 vssd1 vssd1 vccd1 vccd1 net1172 sky130_fd_sc_hd__buf_4
Xfanout1183 net1189 vssd1 vssd1 vccd1 vccd1 net1183 sky130_fd_sc_hd__clkbuf_4
Xfanout1194 net1200 vssd1 vssd1 vccd1 vccd1 net1194 sky130_fd_sc_hd__clkbuf_4
XANTENNA__16631__A2 net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17777_ _02202_ _02371_ _03435_ _03455_ vssd1 vssd1 vccd1 vccd1 _03456_ sky130_fd_sc_hd__or4_1
X_14989_ net2645 net151 _01549_ control.body\[1004\] vssd1 vssd1 vccd1 vccd1 _00326_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_135_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11283__A net1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19516_ clknet_leaf_121_clk net2430 net1401 vssd1 vssd1 vccd1 vccd1 control.body\[874\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_44_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16728_ obsg2.obstacleArray\[112\] net491 net489 obsg2.obstacleArray\[114\] _02406_
+ vssd1 vssd1 vccd1 vccd1 _02407_ sky130_fd_sc_hd__a221o_1
XFILLER_0_88_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16919__B1 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_798 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1471 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16659_ obsg2.obstacleArray\[14\] obsg2.obstacleArray\[15\] net443 vssd1 vssd1 vccd1
+ vccd1 _02338_ sky130_fd_sc_hd__mux2_1
X_19447_ clknet_leaf_110_clk _00391_ net1422 vssd1 vssd1 vccd1 vccd1 control.body\[949\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_48_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16285__S net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16395__B2 net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18066__A net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_100_3360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17592__B1 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_100_3371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09200_ ag2.body\[622\] vssd1 vssd1 vccd1 vccd1 _04225_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_100_3382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12405__B1 net241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19378_ clknet_leaf_112_clk _00322_ net1425 vssd1 vssd1 vccd1 vccd1 control.body\[1008\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__18136__A2 net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__20050__RESET_B net1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11759__A2 net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12956__A1 net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09131_ ag2.body\[440\] vssd1 vssd1 vccd1 vccd1 _04156_ sky130_fd_sc_hd__inv_2
X_18329_ net902 _04519_ _04638_ _08140_ vssd1 vssd1 vccd1 vccd1 _03825_ sky130_fd_sc_hd__a31o_1
X_20637__1554 vssd1 vssd1 vccd1 vccd1 _20637__1554/HI net1554 sky130_fd_sc_hd__conb_1
XFILLER_0_72_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09821__A1 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09062_ ag2.body\[258\] vssd1 vssd1 vccd1 vccd1 _04087_ sky130_fd_sc_hd__inv_2
XANTENNA__13003__A _07519_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16698__A2 net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17895__B2 _03521_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_117_3890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_266 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_113_3765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold600 control.body\[767\] vssd1 vssd1 vccd1 vccd1 net2162 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold611 sound_gen.dac1.dacCount\[2\] vssd1 vssd1 vccd1 vccd1 net2173 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12842__A net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10719__B1 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_113_3776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold622 control.body\[1062\] vssd1 vssd1 vccd1 vccd1 net2184 sky130_fd_sc_hd__dlygate4sd3_1
X_20222_ clknet_leaf_60_clk _01166_ net1468 vssd1 vssd1 vccd1 vccd1 ag2.body\[172\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_25_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold633 control.body\[1056\] vssd1 vssd1 vccd1 vccd1 net2195 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold644 _00264_ vssd1 vssd1 vccd1 vccd1 net2206 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap363 _02076_ vssd1 vssd1 vccd1 vccd1 net363 sky130_fd_sc_hd__buf_4
XFILLER_0_60_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold655 control.body\[1043\] vssd1 vssd1 vccd1 vccd1 net2217 sky130_fd_sc_hd__dlygate4sd3_1
Xhold666 sound_gen.osc1.count\[5\] vssd1 vssd1 vccd1 vccd1 net2228 sky130_fd_sc_hd__dlygate4sd3_1
Xhold677 control.body\[972\] vssd1 vssd1 vccd1 vccd1 net2239 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold688 control.body\[921\] vssd1 vssd1 vccd1 vccd1 net2250 sky130_fd_sc_hd__dlygate4sd3_1
X_20153_ clknet_leaf_96_clk _01097_ net1449 vssd1 vssd1 vccd1 vccd1 ag2.body\[247\]
+ sky130_fd_sc_hd__dfrtp_2
X_09964_ _04934_ _04935_ _04936_ _04933_ vssd1 vssd1 vccd1 vccd1 _04937_ sky130_fd_sc_hd__a211o_1
Xhold699 _00290_ vssd1 vssd1 vccd1 vccd1 net2261 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1115_A net1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16968__B net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20084_ clknet_leaf_77_clk _01028_ net1490 vssd1 vssd1 vccd1 vccd1 ag2.body\[306\]
+ sky130_fd_sc_hd__dfrtp_4
X_09895_ ag2.body\[78\] net1092 vssd1 vssd1 vccd1 vccd1 _04868_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout196_X net196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14769__A net1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout575_A _06649_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16607__C1 net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13673__A net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09870__B net1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16083__B1 net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11193__A net1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1484_A net1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19924__CLK clknet_leaf_52_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout530_X net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout628_X net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_81_2787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_1630 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_81_2798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10670_ _05639_ _05640_ _05641_ _05642_ vssd1 vssd1 vccd1 vccd1 _05643_ sky130_fd_sc_hd__or4_2
XFILLER_0_36_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09329_ net2118 _04336_ vssd1 vssd1 vccd1 vccd1 _01432_ sky130_fd_sc_hd__xor2_1
XFILLER_0_63_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09812__A1 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09885__X _04858_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_11_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12340_ net385 _07306_ vssd1 vssd1 vccd1 vccd1 _07307_ sky130_fd_sc_hd__and2_2
XFILLER_0_84_1628 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout997_X net997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12271_ _07231_ _07240_ vssd1 vssd1 vccd1 vccd1 _07241_ sky130_fd_sc_hd__and2_1
XFILLER_0_120_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14010_ _08167_ _08168_ _08170_ _08166_ vssd1 vssd1 vccd1 vccd1 _08171_ sky130_fd_sc_hd__a211o_1
XANTENNA__19304__CLK clknet_leaf_98_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11222_ net1130 control.body\[860\] vssd1 vssd1 vccd1 vccd1 _06195_ sky130_fd_sc_hd__nand2_1
XANTENNA__15649__B1 _01623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_1347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17607__X _03286_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11153_ ag2.body\[605\] net1097 vssd1 vssd1 vccd1 vccd1 _06126_ sky130_fd_sc_hd__nand2_1
XFILLER_0_120_1526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16878__B net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10104_ net1107 control.body\[941\] vssd1 vssd1 vccd1 vccd1 _05077_ sky130_fd_sc_hd__or2_1
XFILLER_0_21_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15961_ ag2.body\[149\] net198 _01657_ ag2.body\[141\] vssd1 vssd1 vccd1 vccd1 _01191_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__16861__A2 net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11084_ _06053_ _06054_ _06055_ _06056_ vssd1 vssd1 vccd1 vccd1 _06057_ sky130_fd_sc_hd__a22o_1
XANTENNA__14679__A net1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17700_ net416 _03378_ vssd1 vssd1 vccd1 vccd1 _03379_ sky130_fd_sc_hd__or2_1
X_14912_ _05375_ net51 vssd1 vssd1 vccd1 vccd1 _01542_ sky130_fd_sc_hd__and2b_2
X_10035_ _05001_ _05002_ _05003_ vssd1 vssd1 vccd1 vccd1 _05008_ sky130_fd_sc_hd__or3b_1
X_18680_ clknet_leaf_27_clk img_gen.tracker.next_frame\[118\] net1339 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[118\] sky130_fd_sc_hd__dfrtp_1
X_15892_ _04540_ net56 vssd1 vssd1 vccd1 vccd1 _01650_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_123_4061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17631_ ag2.body\[165\] net949 vssd1 vssd1 vccd1 vccd1 _03310_ sky130_fd_sc_hd__xor2_1
XANTENNA__16613__A2 net450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14843_ _08258_ _08562_ _08924_ vssd1 vssd1 vccd1 vccd1 _01514_ sky130_fd_sc_hd__and3_1
XANTENNA__16894__A ag2.body\[209\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12199__A net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1444 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17562_ ag2.body\[580\] net959 vssd1 vssd1 vccd1 vccd1 _03241_ sky130_fd_sc_hd__or2_1
XFILLER_0_86_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14774_ _08927_ _08928_ _01443_ _01444_ vssd1 vssd1 vccd1 vccd1 _01445_ sky130_fd_sc_hd__or4_1
X_11986_ _06938_ _06945_ _06957_ _06951_ net471 net440 vssd1 vssd1 vccd1 vccd1 _06958_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_93_1492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16513_ net399 _02189_ _02191_ net367 vssd1 vssd1 vccd1 vccd1 _02192_ sky130_fd_sc_hd__a211o_1
XANTENNA__11989__A2 net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19301_ clknet_leaf_99_clk _00245_ net1445 vssd1 vssd1 vccd1 vccd1 control.body\[1091\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13725_ net2246 toggle1.nextBlinkToggle\[0\] toggle1.nextBlinkToggle\[1\] net1981
+ vssd1 vssd1 vccd1 vccd1 toggle1.nextDisplayOut\[1\] sky130_fd_sc_hd__a22o_1
X_17493_ ag2.body\[364\] net713 net734 ag2.body\[361\] vssd1 vssd1 vccd1 vccd1 _03172_
+ sky130_fd_sc_hd__o2bb2a_1
X_10937_ ag2.body\[303\] net1066 vssd1 vssd1 vccd1 vccd1 _05910_ sky130_fd_sc_hd__xor2_1
XFILLER_0_86_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17574__B1 net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19232_ clknet_leaf_75_clk _00176_ net1483 vssd1 vssd1 vccd1 vccd1 ag2.body\[95\]
+ sky130_fd_sc_hd__dfrtp_4
X_16444_ _02121_ _02122_ net402 vssd1 vssd1 vccd1 vccd1 _02123_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_267 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13656_ control.divider.count\[19\] _08009_ net221 vssd1 vssd1 vccd1 vccd1 _08012_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_128_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10868_ ag2.body\[532\] net1132 vssd1 vssd1 vccd1 vccd1 _05841_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_136_4466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12646__B net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_136_4477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12938__A1 net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19163_ clknet_leaf_52_clk _00107_ net1363 vssd1 vssd1 vccd1 vccd1 ag2.body\[26\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__11550__B net1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12607_ net627 net438 net468 net569 vssd1 vssd1 vccd1 vccd1 _07505_ sky130_fd_sc_hd__and4_2
XTAP_TAPCELL_ROW_45_1683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16375_ _01709_ net498 _01737_ vssd1 vssd1 vccd1 vccd1 _02054_ sky130_fd_sc_hd__or3_4
XTAP_TAPCELL_ROW_45_1694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13587_ control.divider.count\[5\] _07950_ _07960_ _07961_ vssd1 vssd1 vccd1 vccd1
+ _07962_ sky130_fd_sc_hd__a22o_1
XFILLER_0_87_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10799_ ag2.body\[34\] net1175 vssd1 vssd1 vccd1 vccd1 _05772_ sky130_fd_sc_hd__nand2_1
X_18114_ net44 _03691_ vssd1 vssd1 vccd1 vccd1 _03692_ sky130_fd_sc_hd__nor2_1
XFILLER_0_124_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15326_ control.body\[718\] net73 _01589_ net2349 vssd1 vssd1 vccd1 vccd1 _00624_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11610__A1 net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19094_ clknet_leaf_146_clk img_gen.tracker.next_frame\[532\] net1239 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[532\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_41_1569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12538_ net1936 net651 _07465_ _07466_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[29\]
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_87_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10166__B net1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18045_ obsg2.obstacleArray\[34\] _03646_ net521 vssd1 vssd1 vccd1 vccd1 _01285_
+ sky130_fd_sc_hd__o21a_1
XANTENNA__10964__A3 _04599_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15257_ net2135 net109 net50 net2458 vssd1 vssd1 vccd1 vccd1 _00565_ sky130_fd_sc_hd__a22o_1
XFILLER_0_41_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12469_ _07307_ _07422_ vssd1 vssd1 vccd1 vccd1 _07424_ sky130_fd_sc_hd__or2_1
XANTENNA__12662__A net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14208_ net990 ag2.body\[409\] vssd1 vssd1 vccd1 vccd1 _08369_ sky130_fd_sc_hd__xor2_1
XFILLER_0_111_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12166__A2 net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15188_ net2331 net101 _01572_ control.body\[829\] vssd1 vssd1 vccd1 vccd1 _00503_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_91_3094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11374__B1 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1556 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17724__S1 net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11913__A2 net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14139_ _08296_ _08297_ _08298_ _08299_ vssd1 vssd1 vccd1 vccd1 _08300_ sky130_fd_sc_hd__a22o_1
Xfanout409 net412 vssd1 vssd1 vccd1 vccd1 net409 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19996_ clknet_leaf_63_clk _00940_ net1475 vssd1 vssd1 vccd1 vccd1 ag2.body\[394\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_39_1498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13115__A1 net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18947_ clknet_leaf_5_clk img_gen.tracker.next_frame\[385\] net1269 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[385\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__13666__A2 net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09690__B net1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09680_ ag2.body\[14\] net749 net1054 _03980_ vssd1 vssd1 vccd1 vccd1 _04653_ sky130_fd_sc_hd__a22o_1
XFILLER_0_59_1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18878_ clknet_leaf_27_clk img_gen.tracker.next_frame\[316\] net1281 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[316\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_94_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18821__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17829_ net662 _03491_ vssd1 vssd1 vccd1 vccd1 _01224_ sky130_fd_sc_hd__and2_1
XFILLER_0_136_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_102_3422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_102_3433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_3444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17565__B1 net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout156_A net162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout38 net39 vssd1 vssd1 vccd1 vccd1 net38 sky130_fd_sc_hd__clkbuf_4
Xfanout49 _01631_ vssd1 vssd1 vccd1 vccd1 net49 sky130_fd_sc_hd__buf_2
XFILLER_0_119_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18626__RESET_B net1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16028__B net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_119_3941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12556__B net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_119_3952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_3963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_115_3816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_3827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1065_A net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09114_ ag2.body\[385\] vssd1 vssd1 vccd1 vccd1 _04139_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_21_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_3838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09045_ ag2.body\[223\] vssd1 vssd1 vccd1 vccd1 _04070_ sky130_fd_sc_hd__inv_2
XFILLER_0_44_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09865__B net1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1232_A net1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20304__CLK clknet_leaf_37_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12157__A2 net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13387__B net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold430 img_gen.tracker.frame\[398\] vssd1 vssd1 vccd1 vccd1 net1992 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold441 img_gen.tracker.frame\[141\] vssd1 vssd1 vccd1 vccd1 net2003 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout692_A net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold452 img_gen.tracker.frame\[365\] vssd1 vssd1 vccd1 vccd1 net2014 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10804__B net1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_2580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold463 img_gen.tracker.frame\[395\] vssd1 vssd1 vccd1 vccd1 net2025 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20205_ clknet_leaf_56_clk _01149_ net1456 vssd1 vssd1 vccd1 vccd1 ag2.body\[187\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__15883__A _04539_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_2591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10092__A net1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold474 img_gen.tracker.frame\[96\] vssd1 vssd1 vccd1 vccd1 net2036 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1020_X net1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold485 img_gen.tracker.frame\[447\] vssd1 vssd1 vccd1 vccd1 net2047 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold496 toggle1.bcd_ones\[2\] vssd1 vssd1 vccd1 vccd1 net2058 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1118_X net1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_70_2444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout910 net911 vssd1 vssd1 vccd1 vccd1 net910 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_70_2455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09881__A ag2.body\[162\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20136_ clknet_leaf_80_clk _01080_ net1485 vssd1 vssd1 vccd1 vccd1 ag2.body\[262\]
+ sky130_fd_sc_hd__dfrtp_4
Xfanout921 net922 vssd1 vssd1 vccd1 vccd1 net921 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_70_2466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout932 net933 vssd1 vssd1 vccd1 vccd1 net932 sky130_fd_sc_hd__buf_4
X_09947_ net1146 control.body\[739\] vssd1 vssd1 vccd1 vccd1 _04920_ sky130_fd_sc_hd__or2_1
Xfanout943 obsg2.randCord\[6\] vssd1 vssd1 vccd1 vccd1 net943 sky130_fd_sc_hd__buf_4
XANTENNA__11117__B1 _04861_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout954 net955 vssd1 vssd1 vccd1 vccd1 net954 sky130_fd_sc_hd__buf_2
XANTENNA__16050__Y _01729_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout957_A net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout965 net967 vssd1 vssd1 vccd1 vccd1 net965 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11916__A net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20067_ clknet_leaf_73_clk _01011_ net1501 vssd1 vssd1 vccd1 vccd1 ag2.body\[321\]
+ sky130_fd_sc_hd__dfrtp_2
Xfanout976 ag2.randCord\[3\] vssd1 vssd1 vccd1 vccd1 net976 sky130_fd_sc_hd__buf_4
X_09878_ ag2.body\[166\] net1081 vssd1 vssd1 vccd1 vccd1 _04851_ sky130_fd_sc_hd__or2_1
Xfanout987 net988 vssd1 vssd1 vccd1 vccd1 net987 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_5_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout998 net999 vssd1 vssd1 vccd1 vccd1 net998 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_5_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_5_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_87_2963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_2974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout745_X net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_2985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12880__A3 _07638_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11840_ img_gen.tracker.frame\[503\] net586 net544 img_gen.tracker.frame\[500\] _06811_
+ vssd1 vssd1 vccd1 vccd1 _06812_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_68_2384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_83_2849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_2395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_1632 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12093__A1 _06661_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16359__A1 net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_146_clk clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_146_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_36_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11771_ img_gen.tracker.frame\[95\] net592 net550 img_gen.tracker.frame\[92\] _06742_
+ vssd1 vssd1 vccd1 vccd1 _06743_ sky130_fd_sc_hd__o221a_1
XANTENNA_fanout912_X net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_95_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11651__A net1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13510_ _07612_ _07806_ net676 vssd1 vssd1 vccd1 vccd1 _07916_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_51_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17020__A2 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10722_ _05690_ _05691_ _05692_ _05694_ vssd1 vssd1 vccd1 vccd1 _05695_ sky130_fd_sc_hd__or4_1
X_14490_ net1032 ag2.body\[349\] vssd1 vssd1 vccd1 vccd1 _08651_ sky130_fd_sc_hd__xor2_1
XANTENNA__15031__A1 _04445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13441_ net682 _07888_ vssd1 vssd1 vccd1 vccd1 _07889_ sky130_fd_sc_hd__nor2_1
X_10653_ ag2.body\[286\] net1091 vssd1 vssd1 vccd1 vccd1 _05626_ sky130_fd_sc_hd__xor2_1
XFILLER_0_125_339 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_131_4330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16160_ obsg2.obstacleArray\[24\] obsg2.obstacleArray\[25\] net428 vssd1 vssd1 vccd1
+ vccd1 _01839_ sky130_fd_sc_hd__mux2_1
XFILLER_0_91_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1160 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13372_ net385 _07535_ _07813_ vssd1 vssd1 vccd1 vccd1 _07862_ sky130_fd_sc_hd__and3_1
XFILLER_0_64_996 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10584_ _05545_ _05546_ _05551_ _05556_ vssd1 vssd1 vccd1 vccd1 _05557_ sky130_fd_sc_hd__or4_2
Xclkload19 clknet_leaf_9_clk vssd1 vssd1 vccd1 vccd1 clkload19/Y sky130_fd_sc_hd__inv_6
X_15111_ control.body\[896\] net146 _01554_ net2457 vssd1 vssd1 vccd1 vccd1 _00434_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_49_1556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12323_ _07242_ _07286_ vssd1 vssd1 vccd1 vccd1 _07290_ sky130_fd_sc_hd__and2b_1
XFILLER_0_23_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16091_ obsg2.obstacleArray\[103\] net430 net376 _01769_ vssd1 vssd1 vccd1 vccd1
+ _01770_ sky130_fd_sc_hd__o211a_1
XFILLER_0_50_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09775__B net1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09549__B1 _04520_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13345__A1 net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15042_ net2218 net164 _01556_ control.body\[954\] vssd1 vssd1 vccd1 vccd1 _00372_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_121_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12254_ _07202_ _07223_ vssd1 vssd1 vccd1 vccd1 _07224_ sky130_fd_sc_hd__nor2_1
XANTENNA__10714__B net1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11205_ _06169_ _06170_ _06172_ _06177_ vssd1 vssd1 vccd1 vccd1 _06178_ sky130_fd_sc_hd__or4b_1
XFILLER_0_121_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18284__A1 net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17087__A2 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12632__D net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19850_ clknet_leaf_93_clk _00794_ net1412 vssd1 vssd1 vccd1 vccd1 ag2.body\[536\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_76_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12185_ net1152 ag2.apple_cord\[3\] vssd1 vssd1 vccd1 vccd1 _07157_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_129_4270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18844__CLK clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09791__A net1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18801_ clknet_leaf_18_clk img_gen.tracker.next_frame\[239\] net1358 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[239\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_125_4123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11136_ _06097_ _06102_ _06105_ _06108_ vssd1 vssd1 vccd1 vccd1 _06109_ sky130_fd_sc_hd__or4b_4
XTAP_TAPCELL_ROW_53_1941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19781_ clknet_leaf_127_clk _00725_ net1331 vssd1 vssd1 vccd1 vccd1 ag2.body\[611\]
+ sky130_fd_sc_hd__dfrtp_4
X_16993_ _04017_ net876 net707 ag2.body\[93\] _02669_ vssd1 vssd1 vccd1 vccd1 _02672_
+ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_125_4145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18732_ clknet_leaf_141_clk img_gen.tracker.next_frame\[170\] net1261 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[170\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_34_1362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15944_ ag2.body\[166\] net195 _01653_ ag2.body\[158\] vssd1 vssd1 vccd1 vccd1 _01176_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_121_4009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11067_ _06023_ _06024_ _06027_ _06039_ vssd1 vssd1 vccd1 vccd1 _06040_ sky130_fd_sc_hd__a31o_1
XFILLER_0_95_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_1373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20636__1553 vssd1 vssd1 vccd1 vccd1 _20636__1553/HI net1553 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_30_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09721__B1 _04693_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10018_ _04090_ net1187 net747 ag2.body\[271\] _04987_ vssd1 vssd1 vccd1 vccd1 _04991_
+ sky130_fd_sc_hd__a221o_1
XANTENNA__09638__A1_N net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16598__A1 net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15875_ ag2.body\[216\] net188 _01648_ ag2.body\[208\] vssd1 vssd1 vccd1 vccd1 _01114_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_30_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18663_ clknet_leaf_13_clk img_gen.tracker.next_frame\[101\] net1282 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[101\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__10331__A1 net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18994__CLK clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14826_ net829 ag2.body\[154\] _04046_ net977 _01492_ vssd1 vssd1 vccd1 vccd1 _01497_
+ sky130_fd_sc_hd__o221a_1
X_17614_ _04219_ net858 net688 ag2.body\[607\] _03291_ vssd1 vssd1 vccd1 vccd1 _03293_
+ sky130_fd_sc_hd__a221o_1
X_18594_ clknet_leaf_13_clk img_gen.tracker.next_frame\[32\] net1282 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[32\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_4517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_138_4528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1285 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_138_4539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17545_ ag2.body\[321\] net876 vssd1 vssd1 vccd1 vccd1 _03224_ sky130_fd_sc_hd__nand2_1
X_14757_ net840 ag2.body\[40\] ag2.body\[46\] net798 _08917_ vssd1 vssd1 vccd1 vccd1
+ _08918_ sky130_fd_sc_hd__a221o_1
XFILLER_0_8_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_137_clk clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_137_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__12657__A net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11969_ img_gen.tracker.frame\[511\] net544 _06940_ net560 vssd1 vssd1 vccd1 vccd1
+ _06941_ sky130_fd_sc_hd__o211a_1
XFILLER_0_86_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_47_1756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1273 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_47_1767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13708_ track.highScore\[6\] _08031_ _08046_ _08047_ _08048_ vssd1 vssd1 vccd1 vccd1
+ _08049_ sky130_fd_sc_hd__o221a_1
X_17476_ ag2.body\[129\] net876 vssd1 vssd1 vccd1 vccd1 _03155_ sky130_fd_sc_hd__xnor2_1
X_14688_ net991 _04017_ ag2.body\[91\] net820 _08848_ vssd1 vssd1 vccd1 vccd1 _08849_
+ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_28_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_28_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19215_ clknet_leaf_57_clk _00159_ net1463 vssd1 vssd1 vccd1 vccd1 ag2.body\[78\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_15_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13639_ control.divider.count\[13\] control.divider.count\[12\] _07995_ control.divider.count\[14\]
+ vssd1 vssd1 vccd1 vccd1 _08000_ sky130_fd_sc_hd__a31o_1
X_16427_ net355 _02084_ vssd1 vssd1 vccd1 vccd1 _02106_ sky130_fd_sc_hd__and2_1
XANTENNA__15573__A2 net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_15_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_97_3270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20327__CLK clknet_leaf_105_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1612 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19146_ clknet_leaf_51_clk _00090_ net1367 vssd1 vssd1 vccd1 vccd1 ag2.body\[10\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_97_3281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16358_ _02035_ _02036_ net416 vssd1 vssd1 vccd1 vccd1 _02037_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_97_3292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18063__B _03579_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_3145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11595__B1 net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_3156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13488__A net225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15309_ _04520_ net53 vssd1 vssd1 vccd1 vccd1 _01587_ sky130_fd_sc_hd__nor2_2
XFILLER_0_48_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16289_ obsg2.obstacleArray\[122\] obsg2.obstacleArray\[123\] net407 vssd1 vssd1
+ vccd1 vccd1 _01968_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_93_3167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09685__B net1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19077_ clknet_leaf_29_clk img_gen.tracker.next_frame\[515\] net1335 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[515\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19925__RESET_B net1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10905__A net1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18028_ net432 _01713_ net482 vssd1 vssd1 vccd1 vccd1 _03635_ sky130_fd_sc_hd__and3_1
XFILLER_0_125_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_1380 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10624__B net1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17078__A2 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout206 net207 vssd1 vssd1 vccd1 vccd1 net206 sky130_fd_sc_hd__buf_2
Xfanout217 net218 vssd1 vssd1 vccd1 vccd1 net217 sky130_fd_sc_hd__dlymetal6s2s_1
X_09801_ net1229 control.body\[960\] vssd1 vssd1 vccd1 vccd1 _04774_ sky130_fd_sc_hd__xor2_1
XANTENNA__09960__B1 net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout228 net233 vssd1 vssd1 vccd1 vccd1 net228 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_103_1554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19979_ clknet_leaf_64_clk _00923_ net1474 vssd1 vssd1 vccd1 vccd1 ag2.body\[409\]
+ sky130_fd_sc_hd__dfrtp_4
Xfanout239 net240 vssd1 vssd1 vccd1 vccd1 net239 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_108_3620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_3631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09732_ ag2.body\[88\] net1235 vssd1 vssd1 vccd1 vccd1 _04705_ sky130_fd_sc_hd__nand2_1
XANTENNA__10640__A net1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14112__A net1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10373__A_N net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_3506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09206__A net1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11455__B net1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09663_ net919 net922 vssd1 vssd1 vccd1 vccd1 _04636_ sky130_fd_sc_hd__xor2_4
X_09594_ _04559_ _04562_ _04563_ _04566_ vssd1 vssd1 vccd1 vccd1 _04567_ sky130_fd_sc_hd__or4_1
XANTENNA__18238__B net35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17142__B net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_128_clk clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_128_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout1182_A net1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12567__A net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17538__B1 net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout538_A _01707_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17002__A2 net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10625__A2 net1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_320 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18717__CLK clknet_leaf_144_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10087__A net1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout705_A _04267_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1068_X net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09876__A ag2.body\[163\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15597__B net57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_76_2631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11050__A2 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16513__A1 net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_2642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10374__X _05347_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10815__A net1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1235_X net1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_2653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09028_ ag2.body\[174\] vssd1 vssd1 vccd1 vccd1 _04053_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_72_2506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_2052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_2063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_2074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout695_X net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18266__A1 net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold260 img_gen.tracker.frame\[74\] vssd1 vssd1 vccd1 vccd1 net1822 sky130_fd_sc_hd__dlygate4sd3_1
Xhold271 img_gen.tracker.frame\[356\] vssd1 vssd1 vccd1 vccd1 net1833 sky130_fd_sc_hd__dlygate4sd3_1
Xhold282 img_gen.tracker.frame\[246\] vssd1 vssd1 vccd1 vccd1 net1844 sky130_fd_sc_hd__dlygate4sd3_1
Xhold293 img_gen.tracker.frame\[481\] vssd1 vssd1 vccd1 vccd1 net1855 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout862_X net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17317__B net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout740 net741 vssd1 vssd1 vccd1 vccd1 net740 sky130_fd_sc_hd__buf_4
Xfanout751 net752 vssd1 vssd1 vccd1 vccd1 net751 sky130_fd_sc_hd__buf_4
X_20119_ clknet_leaf_79_clk _01063_ net1488 vssd1 vssd1 vccd1 vccd1 ag2.body\[277\]
+ sky130_fd_sc_hd__dfrtp_4
Xfanout762 net765 vssd1 vssd1 vccd1 vccd1 net762 sky130_fd_sc_hd__buf_4
X_13990_ ag2.body\[127\] net211 _08159_ ag2.body\[119\] vssd1 vssd1 vccd1 vccd1 _00208_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__14022__A net1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout773 net774 vssd1 vssd1 vccd1 vccd1 net773 sky130_fd_sc_hd__buf_4
Xfanout784 net785 vssd1 vssd1 vccd1 vccd1 net784 sky130_fd_sc_hd__buf_4
XFILLER_0_102_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout795 net796 vssd1 vssd1 vccd1 vccd1 net795 sky130_fd_sc_hd__buf_4
XANTENNA__20153__RESET_B net1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12941_ net685 _07667_ vssd1 vssd1 vccd1 vccd1 _07668_ sky130_fd_sc_hd__nor2_1
XANTENNA__16648__S net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15660_ ag2.body\[408\] net144 _01625_ ag2.body\[400\] vssd1 vssd1 vccd1 vccd1 _00922_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_99_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12872_ net245 _07636_ _07637_ net2065 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[192\]
+ sky130_fd_sc_hd__a22o_1
X_14611_ net846 ag2.body\[128\] ag2.body\[133\] net810 _08771_ vssd1 vssd1 vccd1 vccd1
+ _08772_ sky130_fd_sc_hd__o221a_1
XFILLER_0_119_1594 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11823_ img_gen.tracker.frame\[410\] net616 net545 img_gen.tracker.frame\[416\] _06794_
+ vssd1 vssd1 vccd1 vccd1 _06795_ sky130_fd_sc_hd__o221a_1
X_15591_ ag2.body\[474\] net122 _01618_ ag2.body\[466\] vssd1 vssd1 vccd1 vccd1 _00860_
+ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_119_clk clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_119_clk
+ sky130_fd_sc_hd__clkbuf_8
X_17330_ _03005_ _03006_ _03007_ _03008_ vssd1 vssd1 vccd1 vccd1 _03009_ sky130_fd_sc_hd__or4_1
XANTENNA__11381__A net1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10077__B1 _05026_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17620__X _03299_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14542_ net1038 ag2.body\[244\] vssd1 vssd1 vccd1 vccd1 _08703_ sky130_fd_sc_hd__or2_1
XANTENNA__12908__C _07315_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_431 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11754_ img_gen.tracker.frame\[242\] net615 net581 img_gen.tracker.frame\[251\] vssd1
+ vssd1 vccd1 vccd1 _06726_ sky130_fd_sc_hd__o22a_1
XFILLER_0_51_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09482__A2 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16891__B net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10709__B net1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10705_ ag2.body\[16\] net1222 vssd1 vssd1 vccd1 vccd1 _05678_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_12_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17261_ ag2.body\[252\] net964 vssd1 vssd1 vccd1 vccd1 _02940_ sky130_fd_sc_hd__or2_1
X_14473_ _08625_ _08626_ _08629_ _08630_ _08633_ vssd1 vssd1 vccd1 vccd1 _08634_ sky130_fd_sc_hd__a221o_1
X_11685_ _06654_ _06656_ net561 vssd1 vssd1 vccd1 vccd1 _06657_ sky130_fd_sc_hd__mux2_1
X_16212_ net502 _01890_ _01889_ vssd1 vssd1 vccd1 vccd1 _01891_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_102_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19000_ clknet_leaf_2_clk img_gen.tracker.next_frame\[438\] net1249 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[438\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_64_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13424_ net281 _07880_ _07881_ net1761 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[500\]
+ sky130_fd_sc_hd__a22o_1
X_10636_ net1095 control.body\[669\] vssd1 vssd1 vccd1 vccd1 _05609_ sky130_fd_sc_hd__nand2_1
X_17192_ ag2.body\[575\] net929 vssd1 vssd1 vccd1 vccd1 _02871_ sky130_fd_sc_hd__nand2_1
XFILLER_0_52_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkload108 clknet_leaf_85_clk vssd1 vssd1 vccd1 vccd1 clkload108/Y sky130_fd_sc_hd__clkinv_2
XFILLER_0_36_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16143_ obsg2.obstacleArray\[3\] net431 net378 _01821_ vssd1 vssd1 vccd1 vccd1 _01822_
+ sky130_fd_sc_hd__o211a_1
Xclkload119 clknet_leaf_76_clk vssd1 vssd1 vccd1 vccd1 clkload119/Y sky130_fd_sc_hd__inv_8
XFILLER_0_11_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13355_ net249 _07854_ _07855_ net1973 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[457\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__15300__B _01581_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10725__A net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10567_ ag2.body\[515\] net771 net751 ag2.body\[518\] vssd1 vssd1 vccd1 vccd1 _05540_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_126_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12306_ _07210_ _07272_ vssd1 vssd1 vccd1 vccd1 _07273_ sky130_fd_sc_hd__or2_1
XFILLER_0_133_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16074_ obsg2.obstacleArray\[126\] net424 vssd1 vssd1 vccd1 vccd1 _01753_ sky130_fd_sc_hd__or2_1
XANTENNA__19792__CLK clknet_leaf_127_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13286_ net255 _07827_ _07828_ net1794 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[415\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_126_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10498_ _05463_ _05464_ _05466_ _05469_ vssd1 vssd1 vccd1 vccd1 _05471_ sky130_fd_sc_hd__and4_1
XFILLER_0_121_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19902_ clknet_leaf_57_clk _00846_ net1464 vssd1 vssd1 vccd1 vccd1 ag2.body\[492\]
+ sky130_fd_sc_hd__dfrtp_4
X_15025_ control.body\[979\] net167 _01555_ net2535 vssd1 vssd1 vccd1 vccd1 _00357_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_127_4207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12237_ img_gen.updater.commands.cmd_num\[3\] img_gen.updater.commands.cmd_num\[2\]
+ img_gen.updater.commands.cmd_num\[4\] vssd1 vssd1 vccd1 vccd1 _07207_ sky130_fd_sc_hd__or3b_1
XFILLER_0_27_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_36_1413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12940__A net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16807__A2 net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19833_ clknet_leaf_122_clk _00777_ net1407 vssd1 vssd1 vccd1 vccd1 ag2.body\[567\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_62_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12168_ img_gen.tracker.frame\[429\] net584 net571 vssd1 vssd1 vccd1 vccd1 _07140_
+ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_9_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11119_ net1227 control.body\[864\] vssd1 vssd1 vccd1 vccd1 _06092_ sky130_fd_sc_hd__xor2_1
XFILLER_0_78_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19764_ clknet_leaf_127_clk _00708_ net1326 vssd1 vssd1 vccd1 vccd1 control.body\[626\]
+ sky130_fd_sc_hd__dfrtp_1
X_16976_ ag2.body\[424\] net883 vssd1 vssd1 vccd1 vccd1 _02655_ sky130_fd_sc_hd__xnor2_1
X_12099_ net570 _07070_ _07068_ net468 vssd1 vssd1 vccd1 vccd1 _07071_ sky130_fd_sc_hd__o211a_1
XANTENNA__09026__A ag2.body\[166\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11275__B net1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18715_ clknet_leaf_144_clk img_gen.tracker.next_frame\[153\] net1252 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[153\] sky130_fd_sc_hd__dfrtp_1
Xinput6 gpio_in[29] vssd1 vssd1 vccd1 vccd1 net6 sky130_fd_sc_hd__clkbuf_1
X_15927_ ag2.body\[182\] net136 _01654_ ag2.body\[174\] vssd1 vssd1 vccd1 vccd1 _01160_
+ sky130_fd_sc_hd__a22o_1
X_19695_ clknet_leaf_136_clk _00639_ net1302 vssd1 vssd1 vccd1 vccd1 control.body\[701\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_49_1807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_1818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19172__CLK clknet_leaf_53_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18646_ clknet_leaf_130_clk img_gen.tracker.next_frame\[84\] net1315 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[84\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_49_1829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15858_ ag2.body\[233\] net172 _01646_ ag2.body\[225\] vssd1 vssd1 vccd1 vccd1 _01099_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_133_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13490__B _07505_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14809_ net818 ag2.body\[379\] _04138_ net1009 vssd1 vssd1 vccd1 vccd1 _01480_ sky130_fd_sc_hd__a2bb2o_1
X_18577_ clknet_leaf_15_clk img_gen.tracker.next_frame\[15\] net1278 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[15\] sky130_fd_sc_hd__dfrtp_1
X_15789_ ag2.body\[299\] net208 _01639_ ag2.body\[291\] vssd1 vssd1 vccd1 vccd1 _01037_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_34_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11291__A net1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17528_ ag2.body\[277\] net951 vssd1 vssd1 vccd1 vccd1 _03207_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_99_3332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_99_3343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_3354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10619__B net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_95_3207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17459_ ag2.body\[432\] net737 net732 ag2.body\[433\] vssd1 vssd1 vccd1 vccd1 _03138_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_131_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16293__S net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_3218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12674__X _07542_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_3229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09696__A net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20470_ clknet_leaf_33_clk _01357_ net1346 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[106\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_104_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkload58_A clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19129_ clknet_leaf_132_clk img_gen.tracker.next_frame\[567\] net1297 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[567\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10635__A net1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10354__B net1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1028_A net1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout390_A net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17137__B net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout488_A net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14809__B2 net1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11466__A _04419_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1384 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09207__Y _04232_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10370__A net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16976__B net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09715_ net641 _04602_ vssd1 vssd1 vccd1 vccd1 _04688_ sky130_fd_sc_hd__nor2_2
XFILLER_0_39_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_1522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_84_2900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_1582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout276_X net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1397_A net1404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09646_ net1196 control.body\[745\] vssd1 vssd1 vccd1 vccd1 _04619_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_65_2310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_638 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09577_ net899 net902 net906 vssd1 vssd1 vccd1 vccd1 _04550_ sky130_fd_sc_hd__and3_4
XANTENNA_fanout822_A net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout443_X net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1185_X net1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1046 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10059__B1 net1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09464__A2 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17600__B net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16195__C1 net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout610_X net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_14_Right_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout708_X net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_2704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_968 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_2715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11470_ ag2.body\[488\] net1233 vssd1 vssd1 vccd1 vccd1 _06443_ sky130_fd_sc_hd__xor2_1
XANTENNA_clkbuf_4_6__f_clk_A clknet_3_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_2114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12744__B _07575_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_2125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20635__1552 vssd1 vssd1 vccd1 vccd1 _20635__1552/HI net1552 sky130_fd_sc_hd__conb_1
XFILLER_0_107_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_2136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10421_ net1135 control.body\[1068\] vssd1 vssd1 vccd1 vccd1 _05394_ sky130_fd_sc_hd__nand2_1
XFILLER_0_61_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20599_ net1531 vssd1 vssd1 vccd1 vccd1 gpio_oeb[11] sky130_fd_sc_hd__buf_2
XFILLER_0_21_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13140_ _07592_ _07639_ vssd1 vssd1 vccd1 vccd1 _07762_ sky130_fd_sc_hd__nor2_1
XFILLER_0_46_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10352_ ag2.body\[292\] net764 net757 ag2.body\[293\] _05324_ vssd1 vssd1 vccd1 vccd1
+ _05325_ sky130_fd_sc_hd__a221o_1
XFILLER_0_123_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13071_ _07558_ _07639_ vssd1 vssd1 vccd1 vccd1 _07729_ sky130_fd_sc_hd__nor2_1
X_10283_ ag2.body\[329\] net1212 vssd1 vssd1 vccd1 vccd1 _05256_ sky130_fd_sc_hd__or2_1
XFILLER_0_103_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16232__A net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout91_X net91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12022_ img_gen.tracker.frame\[195\] net612 net595 img_gen.tracker.frame\[201\] vssd1
+ vssd1 vccd1 vccd1 _06994_ sky130_fd_sc_hd__a22o_1
Xfanout1502 net1504 vssd1 vssd1 vccd1 vccd1 net1502 sky130_fd_sc_hd__buf_2
Xfanout1513 net1514 vssd1 vssd1 vccd1 vccd1 net1513 sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_23_Right_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16830_ ag2.body\[226\] net726 net711 ag2.body\[228\] _02503_ vssd1 vssd1 vccd1 vccd1
+ _02509_ sky130_fd_sc_hd__o221a_1
XANTENNA__19195__CLK clknet_leaf_53_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout570 net573 vssd1 vssd1 vccd1 vccd1 net570 sky130_fd_sc_hd__clkbuf_2
Xfanout581 net582 vssd1 vssd1 vccd1 vccd1 net581 sky130_fd_sc_hd__clkbuf_2
XANTENNA__11095__B net1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout592 _06524_ vssd1 vssd1 vccd1 vccd1 net592 sky130_fd_sc_hd__clkbuf_4
X_16761_ obsg2.obstacleArray\[20\] net494 net485 obsg2.obstacleArray\[21\] _02439_
+ vssd1 vssd1 vccd1 vccd1 _02440_ sky130_fd_sc_hd__a221o_1
X_13973_ _05162_ net60 vssd1 vssd1 vccd1 vccd1 _08158_ sky130_fd_sc_hd__nor2_2
XANTENNA__12287__A1 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10298__B1 _05255_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18500_ net1514 net1508 vssd1 vssd1 vccd1 vccd1 _00031_ sky130_fd_sc_hd__or2_1
X_15712_ _06041_ net67 vssd1 vssd1 vccd1 vccd1 _01630_ sky130_fd_sc_hd__and2_2
XANTENNA__20172__CLK clknet_leaf_83_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17214__A2 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12924_ net673 _07659_ vssd1 vssd1 vccd1 vccd1 _07660_ sky130_fd_sc_hd__nor2_1
X_16692_ _02262_ _02370_ _02362_ _02209_ vssd1 vssd1 vccd1 vccd1 _02371_ sky130_fd_sc_hd__a211oi_1
X_19480_ clknet_leaf_110_clk _00424_ net1418 vssd1 vssd1 vccd1 vccd1 control.body\[918\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18431_ _03914_ _03916_ _03919_ vssd1 vssd1 vccd1 vccd1 _03920_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_69_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15643_ ag2.body\[425\] net138 _01623_ ag2.body\[417\] vssd1 vssd1 vccd1 vccd1 _00907_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__17998__A net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12855_ net239 _07628_ _07629_ net1730 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[183\]
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_17_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11806_ img_gen.tracker.frame\[449\] net597 vssd1 vssd1 vccd1 vccd1 _06778_ sky130_fd_sc_hd__or2_1
XFILLER_0_69_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_96_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15574_ ag2.body\[492\] net135 _01615_ ag2.body\[484\] vssd1 vssd1 vccd1 vccd1 _00846_
+ sky130_fd_sc_hd__a22o_1
X_18362_ _07181_ _03819_ vssd1 vssd1 vccd1 vccd1 _03857_ sky130_fd_sc_hd__nor2_1
XFILLER_0_29_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12786_ net669 _07596_ vssd1 vssd1 vccd1 vccd1 _07597_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_32_Right_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18175__B1 net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17313_ _02986_ _02987_ _02990_ _02991_ vssd1 vssd1 vccd1 vccd1 _02992_ sky130_fd_sc_hd__a211o_1
X_14525_ net992 ag2.body\[249\] vssd1 vssd1 vccd1 vccd1 _08686_ sky130_fd_sc_hd__nand2_1
XFILLER_0_84_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17510__B net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11737_ img_gen.tracker.frame\[47\] net590 net553 img_gen.tracker.frame\[44\] _06708_
+ vssd1 vssd1 vccd1 vccd1 _06709_ sky130_fd_sc_hd__o221a_1
XFILLER_0_84_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19588__RESET_B net1386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18293_ _08052_ _03783_ _03788_ _08053_ vssd1 vssd1 vccd1 vccd1 _03789_ sky130_fd_sc_hd__a31o_1
XANTENNA__11893__S0 net1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12935__A _07476_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18190__A3 _03705_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14456_ net827 ag2.body\[434\] _04155_ net1008 _08616_ vssd1 vssd1 vccd1 vccd1 _08617_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_126_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17244_ ag2.body\[619\] net715 net698 ag2.body\[622\] vssd1 vssd1 vccd1 vccd1 _02923_
+ sky130_fd_sc_hd__o2bb2a_1
X_11668_ net1169 net1122 vssd1 vssd1 vccd1 vccd1 _06640_ sky130_fd_sc_hd__nand2_4
XFILLER_0_98_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13407_ net234 _07874_ _07875_ net1690 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[489\]
+ sky130_fd_sc_hd__a22o_1
X_17175_ ag2.body\[463\] net930 vssd1 vssd1 vccd1 vccd1 _02854_ sky130_fd_sc_hd__nand2_1
X_10619_ ag2.body\[55\] net1055 vssd1 vssd1 vccd1 vccd1 _05592_ sky130_fd_sc_hd__xor2_1
XANTENNA__15030__B net66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14387_ net975 _04098_ _04100_ net1022 vssd1 vssd1 vccd1 vccd1 _08548_ sky130_fd_sc_hd__a22o_1
X_11599_ obsg2.obstacleArray\[16\] obsg2.obstacleArray\[20\] net514 vssd1 vssd1 vccd1
+ vccd1 _06572_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16126_ obsg2.obstacleArray\[90\] obsg2.obstacleArray\[91\] net428 vssd1 vssd1 vccd1
+ vccd1 _01805_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13338_ net664 _07848_ vssd1 vssd1 vccd1 vccd1 _07849_ sky130_fd_sc_hd__nor2_1
XFILLER_0_45_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10174__B net1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16057_ net956 net538 vssd1 vssd1 vccd1 vccd1 _01736_ sky130_fd_sc_hd__nor2_2
XFILLER_0_122_684 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13269_ net670 _07821_ vssd1 vssd1 vccd1 vccd1 _07822_ sky130_fd_sc_hd__nor2_1
XANTENNA__12670__A net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_41_Right_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_1350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19538__CLK clknet_leaf_115_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15008_ control.body\[997\] net166 _01552_ control.body\[989\] vssd1 vssd1 vccd1
+ vccd1 _00343_ sky130_fd_sc_hd__a22o_1
XANTENNA__11317__A3 _05074_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_88_3000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_88_3011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13485__B net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_88_3022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11286__A net1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19816_ clknet_leaf_125_clk _00760_ net1410 vssd1 vssd1 vccd1 vccd1 ag2.body\[582\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__16110__C1 net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20515__CLK clknet_leaf_113_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19747_ clknet_leaf_129_clk net2417 net1325 vssd1 vssd1 vccd1 vccd1 control.body\[641\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__16288__S net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16959_ ag2.body\[288\] net885 vssd1 vssd1 vccd1 vccd1 _02638_ sky130_fd_sc_hd__xor2_1
XFILLER_0_75_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18562__CLK clknet_leaf_15_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18069__A net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09500_ ag2.body\[402\] net1185 vssd1 vssd1 vccd1 vccd1 _04473_ sky130_fd_sc_hd__nand2_1
XANTENNA__17205__A2 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19678_ clknet_leaf_135_clk _00622_ net1386 vssd1 vssd1 vccd1 vccd1 control.body\[716\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__16413__B1 net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09431_ net927 net1127 vssd1 vssd1 vccd1 vccd1 _04404_ sky130_fd_sc_hd__or2_1
XFILLER_0_2_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18629_ clknet_leaf_0_clk img_gen.tracker.next_frame\[67\] net1242 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[67\] sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_50_Right_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_1490 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09362_ sound_gen.osc1.stayCount\[11\] sound_gen.osc1.stayCount\[10\] _04363_ vssd1
+ vssd1 vccd1 vccd1 _04364_ sky130_fd_sc_hd__and3_1
XFILLER_0_136_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_250 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09293_ sound_gen.osc1.count\[2\] _04308_ _04309_ _04312_ vssd1 vssd1 vccd1 vccd1
+ _04313_ sky130_fd_sc_hd__a211o_1
XANTENNA__12450__A1 net1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10917__X _05890_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_11 _03446_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout236_A net247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_22 _08699_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_33 _03442_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20522_ clknet_leaf_93_clk track.nextCurrScore\[4\] net1413 vssd1 vssd1 vccd1 vccd1
+ control.body_update.curr_length\[4\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_62_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_676 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16036__B net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18469__A1 net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12202__A1 _07147_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20453_ clknet_leaf_38_clk _01340_ net1354 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[89\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_16_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10365__A net1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1145_A net1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20384_ clknet_leaf_41_clk _01271_ net1372 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[20\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_101_802 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17692__A2 net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12580__A _06671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11908__B net1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout772_A _04230_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout393_X net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11713__B1 net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18905__CLK clknet_leaf_144_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20195__CLK clknet_leaf_88_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1100_X net1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout560_X net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16198__S net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10970_ net1230 control.body\[1000\] vssd1 vssd1 vccd1 vccd1 _05943_ sky130_fd_sc_hd__xnor2_1
XANTENNA__14300__A net1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09629_ net910 net905 net918 net914 vssd1 vssd1 vccd1 vccd1 _04602_ sky130_fd_sc_hd__and4_2
XANTENNA_fanout825_X net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17170__X _02849_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12640_ _06671_ _07522_ vssd1 vssd1 vccd1 vccd1 _07523_ sky130_fd_sc_hd__or2_2
XANTENNA__09888__X _04861_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14966__B1 net51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12441__A1 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12571_ net267 _07484_ _07485_ net1769 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[43\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_13_1547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16227__A net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_50_clk clknet_4_6__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_50_clk
+ sky130_fd_sc_hd__clkbuf_8
X_14310_ net1034 ag2.body\[52\] vssd1 vssd1 vccd1 vccd1 _08471_ sky130_fd_sc_hd__nand2_1
XFILLER_0_13_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11522_ _06479_ _06482_ _06494_ vssd1 vssd1 vccd1 vccd1 _06495_ sky130_fd_sc_hd__a21o_1
XFILLER_0_87_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15290_ control.body\[751\] net87 _01584_ control.body\[743\] vssd1 vssd1 vccd1 vccd1
+ _00593_ sky130_fd_sc_hd__a22o_1
XFILLER_0_92_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14194__A1 net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14241_ _08399_ _08400_ _08401_ vssd1 vssd1 vccd1 vccd1 _08402_ sky130_fd_sc_hd__nor3b_1
XANTENNA__14194__B2 net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11453_ _06420_ _06421_ _06422_ _06425_ vssd1 vssd1 vccd1 vccd1 _06426_ sky130_fd_sc_hd__or4_4
XANTENNA__16661__S net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_12_Left_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18442__A net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10204__B1 _05160_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20515__RESET_B net1403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10404_ net1183 control.body\[1074\] vssd1 vssd1 vccd1 vccd1 _05377_ sky130_fd_sc_hd__xor2_1
X_14172_ _08328_ _08330_ _08332_ vssd1 vssd1 vccd1 vccd1 _08333_ sky130_fd_sc_hd__or3_1
XANTENNA__15785__B net60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11384_ net1146 control.body\[643\] vssd1 vssd1 vccd1 vccd1 _06357_ sky130_fd_sc_hd__nand2_1
XANTENNA__12761__Y _07584_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16233__Y _01912_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11952__B1 net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13123_ net243 _07752_ _07753_ net1686 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[327\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_104_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10335_ ag2.body\[524\] net1136 vssd1 vssd1 vccd1 vccd1 _05308_ sky130_fd_sc_hd__nand2_1
XFILLER_0_127_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17683__A2 net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18980_ clknet_leaf_8_clk img_gen.tracker.next_frame\[418\] net1270 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[418\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_131_492 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17931_ net298 _03562_ vssd1 vssd1 vccd1 vccd1 _03563_ sky130_fd_sc_hd__and2_1
X_13054_ net680 _07720_ vssd1 vssd1 vccd1 vccd1 _07721_ sky130_fd_sc_hd__nor2_1
X_10266_ _05237_ _05238_ vssd1 vssd1 vccd1 vccd1 _05239_ sky130_fd_sc_hd__and2_1
XFILLER_0_24_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18585__CLK clknet_leaf_15_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1310 net1311 vssd1 vssd1 vccd1 vccd1 net1310 sky130_fd_sc_hd__clkbuf_2
X_12005_ img_gen.tracker.frame\[478\] net578 net568 vssd1 vssd1 vccd1 vccd1 _06977_
+ sky130_fd_sc_hd__o21a_1
Xfanout1321 net1323 vssd1 vssd1 vccd1 vccd1 net1321 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_84_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17862_ _03500_ _03512_ vssd1 vssd1 vccd1 vccd1 _01236_ sky130_fd_sc_hd__and2_1
Xfanout1332 net1333 vssd1 vssd1 vccd1 vccd1 net1332 sky130_fd_sc_hd__clkbuf_2
X_10197_ _05164_ _05165_ _05166_ _05167_ vssd1 vssd1 vccd1 vccd1 _05170_ sky130_fd_sc_hd__a22o_1
Xfanout1343 net1344 vssd1 vssd1 vccd1 vccd1 net1343 sky130_fd_sc_hd__clkbuf_4
Xfanout1354 net1355 vssd1 vssd1 vccd1 vccd1 net1354 sky130_fd_sc_hd__clkbuf_4
X_19601_ clknet_leaf_118_clk _00545_ net1393 vssd1 vssd1 vccd1 vccd1 control.body\[799\]
+ sky130_fd_sc_hd__dfrtp_1
X_16813_ ag2.body\[82\] net865 vssd1 vssd1 vccd1 vccd1 _02492_ sky130_fd_sc_hd__xnor2_1
Xfanout1365 net1366 vssd1 vssd1 vccd1 vccd1 net1365 sky130_fd_sc_hd__clkbuf_4
Xfanout1376 net1377 vssd1 vssd1 vccd1 vccd1 net1376 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_75_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17793_ net1009 _03466_ _03464_ vssd1 vssd1 vccd1 vccd1 _01213_ sky130_fd_sc_hd__o21a_1
Xfanout1387 net1389 vssd1 vssd1 vccd1 vccd1 net1387 sky130_fd_sc_hd__clkbuf_4
Xfanout1398 net1400 vssd1 vssd1 vccd1 vccd1 net1398 sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_21_Left_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19532_ clknet_leaf_118_clk _00476_ net1388 vssd1 vssd1 vccd1 vccd1 control.body\[858\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_117_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16744_ obsg2.obstacleArray\[39\] net500 net486 obsg2.obstacleArray\[38\] _02420_
+ vssd1 vssd1 vccd1 vccd1 _02423_ sky130_fd_sc_hd__a221o_1
XANTENNA__14210__A net1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13956_ ag2.body\[96\] net189 _08156_ ag2.body\[88\] vssd1 vssd1 vccd1 vccd1 _00177_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12649__B _07528_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17738__A3 _02642_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19463_ clknet_leaf_110_clk net2282 net1418 vssd1 vssd1 vccd1 vccd1 control.body\[933\]
+ sky130_fd_sc_hd__dfrtp_1
X_12907_ net293 _07650_ _07651_ net1977 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[212\]
+ sky130_fd_sc_hd__a22o_1
X_16675_ obsg2.obstacleArray\[26\] net447 vssd1 vssd1 vccd1 vccd1 _02354_ sky130_fd_sc_hd__or2_1
X_13887_ ag2.body\[35\] net119 _08148_ ag2.body\[27\] vssd1 vssd1 vccd1 vccd1 _00116_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_53_1327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18414_ _03841_ _03890_ _03903_ _08144_ vssd1 vssd1 vccd1 vccd1 _03904_ sky130_fd_sc_hd__a211o_1
XFILLER_0_69_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15626_ ag2.body\[442\] net125 _01621_ ag2.body\[434\] vssd1 vssd1 vccd1 vccd1 _00892_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_97_991 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12838_ net261 _07619_ _07620_ net1679 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[175\]
+ sky130_fd_sc_hd__a22o_1
X_19394_ clknet_leaf_103_clk _00338_ net1427 vssd1 vssd1 vccd1 vccd1 control.body\[992\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18345_ net906 _04644_ _08030_ _08036_ _03820_ vssd1 vssd1 vccd1 vccd1 _03841_ sky130_fd_sc_hd__a311o_2
X_15557_ ag2.body\[510\] net187 _01612_ ag2.body\[502\] vssd1 vssd1 vccd1 vccd1 _00832_
+ sky130_fd_sc_hd__a22o_1
X_12769_ net672 _07588_ vssd1 vssd1 vccd1 vccd1 _07589_ sky130_fd_sc_hd__nor2_1
XFILLER_0_33_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_41_clk clknet_4_7__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_41_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_127_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14508_ net1037 ag2.body\[180\] vssd1 vssd1 vccd1 vccd1 _08669_ sky130_fd_sc_hd__xor2_1
X_18276_ net319 _03575_ obsg2.obstacleArray\[135\] vssd1 vssd1 vccd1 vccd1 _03777_
+ sky130_fd_sc_hd__a21oi_1
X_15488_ _05192_ net54 vssd1 vssd1 vccd1 vccd1 _01606_ sky130_fd_sc_hd__nor2_2
XFILLER_0_115_916 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__20068__CLK clknet_leaf_73_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17227_ ag2.body\[313\] net736 net713 ag2.body\[316\] _02905_ vssd1 vssd1 vccd1 vccd1
+ _02906_ sky130_fd_sc_hd__o221a_1
XANTENNA_clkbuf_leaf_20_clk_X clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14439_ net840 ag2.body\[16\] _03983_ net1035 _08599_ vssd1 vssd1 vccd1 vccd1 _08600_
+ sky130_fd_sc_hd__a221o_1
XANTENNA__16424__X _02103_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18352__A _04646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13932__B2 ag2.body\[67\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold804 sound_gen.osc1.stayCount\[3\] vssd1 vssd1 vccd1 vccd1 net2366 sky130_fd_sc_hd__dlygate4sd3_1
X_17158_ _02831_ _02832_ _02835_ _02836_ vssd1 vssd1 vccd1 vccd1 _02837_ sky130_fd_sc_hd__or4b_2
Xhold815 control.body\[676\] vssd1 vssd1 vccd1 vccd1 net2377 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold826 control.body\[916\] vssd1 vssd1 vccd1 vccd1 net2388 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold837 sound_gen.osc1.stayCount\[1\] vssd1 vssd1 vccd1 vccd1 net2399 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16109_ obsg2.obstacleArray\[87\] net431 net378 _01787_ vssd1 vssd1 vccd1 vccd1 _01788_
+ sky130_fd_sc_hd__o211a_1
XANTENNA__13496__A net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold848 _00400_ vssd1 vssd1 vccd1 vccd1 net2410 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__17674__A2 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09693__B net1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17089_ _02757_ _02762_ _02767_ vssd1 vssd1 vccd1 vccd1 _02768_ sky130_fd_sc_hd__or3_2
X_09980_ _04951_ _04952_ vssd1 vssd1 vccd1 vccd1 _04953_ sky130_fd_sc_hd__nand2_1
Xhold859 control.body\[717\] vssd1 vssd1 vccd1 vccd1 net2421 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12335__A_N _07301_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11728__B net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17831__C1 net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout186_A net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20634__1551 vssd1 vssd1 vccd1 vccd1 _20634__1551/HI net1551 sky130_fd_sc_hd__conb_1
XFILLER_0_100_1398 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14120__A net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12120__B1 net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12671__A1 net242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout353_A net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16746__S net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09414_ img_gen.control.current\[1\] img_gen.control.current\[0\] vssd1 vssd1 vccd1
+ vccd1 _04393_ sky130_fd_sc_hd__and2_4
XANTENNA_fanout1095_A net1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12846__Y _07624_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18246__B net35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09345_ sound_gen.osc1.stayCount\[19\] sound_gen.osc1.stayCount\[18\] sound_gen.osc1.stayCount\[17\]
+ _04348_ vssd1 vssd1 vccd1 vccd1 _04349_ sky130_fd_sc_hd__and4_1
XANTENNA__09868__B net1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout520_A net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17150__B net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12575__A net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14119__X _08280_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16047__A net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_32_clk clknet_4_5__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_32_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout239_X net239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1262_A net1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout618_A net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__20565__Q obsg2.randCord\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_1472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09276_ sound_gen.osc1.stayCount\[18\] _04288_ _04297_ _04298_ vssd1 vssd1 vccd1
+ vccd1 _04299_ sky130_fd_sc_hd__o211a_1
XANTENNA__17901__A3 net48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20505_ clknet_leaf_132_clk coll.nextBadColl net1304 vssd1 vssd1 vccd1 vccd1 coll.badColl
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__15373__B1 _01594_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16481__S net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10095__A net1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14790__A net1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout406_X net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1148_X net1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13923__A1 ag2.body\[67\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13923__B2 ag2.body\[59\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20436_ clknet_leaf_26_clk _01323_ net1343 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[72\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__16053__Y _01732_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout987_A net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11934__B1 net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11919__A net1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20367_ clknet_leaf_21_clk _01254_ net1362 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[3\]
+ sky130_fd_sc_hd__dfrtp_2
X_10120_ _05089_ _05090_ _05091_ _05092_ vssd1 vssd1 vccd1 vccd1 _05093_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout99_A net100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20298_ clknet_leaf_36_clk control.divider.next_count\[19\] net1347 vssd1 vssd1 vccd1
+ vccd1 control.divider.count\[19\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_100_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10542__B net1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout775_X net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_99_clk clknet_4_11__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_99_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_105_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17165__X _02844_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10051_ ag2.body\[486\] net1080 vssd1 vssd1 vccd1 vccd1 _05024_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09890__Y _04863_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout942_X net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11654__A net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13810_ control.divider.fsm.current_mode\[2\] control.divider.fsm.current_mode\[0\]
+ _08109_ vssd1 vssd1 vccd1 vccd1 _00078_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_19_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14790_ net1039 ag2.body\[548\] vssd1 vssd1 vccd1 vccd1 _01461_ sky130_fd_sc_hd__xor2_1
XFILLER_0_97_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout54_X net54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12111__B1 net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11373__B net1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1051 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13741_ _07209_ _07214_ vssd1 vssd1 vccd1 vccd1 _08062_ sky130_fd_sc_hd__or2_1
XFILLER_0_35_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10953_ ag2.body\[171\] net1154 vssd1 vssd1 vccd1 vccd1 _05926_ sky130_fd_sc_hd__xor2_1
XANTENNA__17979__C net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17050__B1 net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16460_ _02086_ _02135_ _02138_ _02104_ _02107_ vssd1 vssd1 vccd1 vccd1 _02139_ sky130_fd_sc_hd__o311a_1
X_13672_ net465 _08019_ _08020_ vssd1 vssd1 vccd1 vccd1 track.nextCurrScore\[0\] sky130_fd_sc_hd__and3_1
X_10884_ _04556_ _04601_ _05856_ vssd1 vssd1 vccd1 vccd1 _05857_ sky130_fd_sc_hd__o21ai_2
X_12623_ net231 _07513_ _07514_ net1837 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[66\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_6_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15411_ net2309 net83 _01597_ control.body\[627\] vssd1 vssd1 vccd1 vccd1 _00701_
+ sky130_fd_sc_hd__a22o_1
X_16391_ net398 _02069_ vssd1 vssd1 vccd1 vccd1 _02070_ sky130_fd_sc_hd__or2_1
XFILLER_0_52_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12485__A net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_23_clk clknet_4_6__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_23_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_38_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18130_ obsg2.obstacleArray\[64\] _03701_ net530 vssd1 vssd1 vccd1 vccd1 _01315_
+ sky130_fd_sc_hd__o21a_1
X_15342_ control.body\[701\] net72 _01590_ net2225 vssd1 vssd1 vccd1 vccd1 _00639_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__19383__CLK clknet_leaf_93_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12554_ net329 _07475_ vssd1 vssd1 vccd1 vccd1 _07476_ sky130_fd_sc_hd__or2_2
XFILLER_0_87_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_253 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11505_ net1197 net1174 vssd1 vssd1 vccd1 vccd1 _06478_ sky130_fd_sc_hd__xor2_2
XANTENNA__14167__A1 net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18061_ net42 _03656_ vssd1 vssd1 vccd1 vccd1 _03657_ sky130_fd_sc_hd__nor2_1
XANTENNA__14167__B2 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15364__B1 _01593_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15273_ _04605_ net54 vssd1 vssd1 vccd1 vccd1 _01583_ sky130_fd_sc_hd__nor2_2
XANTENNA__16561__C1 net357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12485_ net678 _07436_ vssd1 vssd1 vccd1 vccd1 _07437_ sky130_fd_sc_hd__nor2_1
XFILLER_0_48_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14224_ net843 ag2.body\[392\] ag2.body\[399\] net793 _08384_ vssd1 vssd1 vccd1 vccd1
+ _08385_ sky130_fd_sc_hd__a221o_1
X_17012_ ag2.body\[497\] net735 net932 _04183_ _02690_ vssd1 vssd1 vccd1 vccd1 _02691_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_80_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13914__A1 ag2.body\[59\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20360__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09794__A net1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11436_ ag2.body\[395\] net1162 vssd1 vssd1 vccd1 vccd1 _06409_ sky130_fd_sc_hd__xor2_1
XANTENNA__11925__B1 net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12932__B net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15116__B1 _01554_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11829__A net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14155_ net1034 ag2.body\[620\] vssd1 vssd1 vccd1 vccd1 _08316_ sky130_fd_sc_hd__xor2_1
X_11367_ _06329_ _06330_ _06338_ _06339_ vssd1 vssd1 vccd1 vccd1 _06340_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13106_ net673 _07745_ vssd1 vssd1 vccd1 vccd1 _07746_ sky130_fd_sc_hd__nor2_1
XFILLER_0_123_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16864__B1 net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10318_ ag2.body\[612\] net1120 vssd1 vssd1 vccd1 vccd1 _05291_ sky130_fd_sc_hd__nand2_1
XFILLER_0_123_1354 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14086_ net983 ag2.body\[282\] vssd1 vssd1 vccd1 vccd1 _08247_ sky130_fd_sc_hd__or2_1
X_18963_ clknet_leaf_7_clk img_gen.tracker.next_frame\[401\] net1266 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[401\] sky130_fd_sc_hd__dfrtp_1
X_11298_ net1118 control.body\[684\] vssd1 vssd1 vccd1 vccd1 _06271_ sky130_fd_sc_hd__xor2_1
XANTENNA__13678__B1 net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10452__B net1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17914_ _01691_ _03535_ _03548_ vssd1 vssd1 vccd1 vccd1 _03549_ sky130_fd_sc_hd__a21o_2
X_13037_ net342 _07542_ vssd1 vssd1 vccd1 vccd1 _07713_ sky130_fd_sc_hd__nor2_1
XANTENNA__17408__A2 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10249_ _05210_ _05212_ _05217_ _05221_ vssd1 vssd1 vccd1 vccd1 _05222_ sky130_fd_sc_hd__or4_4
XFILLER_0_119_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18894_ clknet_leaf_26_clk img_gen.tracker.next_frame\[332\] net1339 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[332\] sky130_fd_sc_hd__dfrtp_1
Xfanout1140 net1142 vssd1 vssd1 vccd1 vccd1 net1140 sky130_fd_sc_hd__buf_4
Xfanout1151 net1156 vssd1 vssd1 vccd1 vccd1 net1151 sky130_fd_sc_hd__buf_2
X_17845_ _04277_ _03500_ vssd1 vssd1 vccd1 vccd1 _03501_ sky130_fd_sc_hd__nor2_1
Xfanout1162 net1166 vssd1 vssd1 vccd1 vccd1 net1162 sky130_fd_sc_hd__buf_4
XANTENNA__16711__S0 net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1173 net1189 vssd1 vssd1 vccd1 vccd1 net1173 sky130_fd_sc_hd__clkbuf_4
XANTENNA__16092__A1 net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1184 net1188 vssd1 vssd1 vccd1 vccd1 net1184 sky130_fd_sc_hd__buf_4
Xfanout1195 net1200 vssd1 vssd1 vccd1 vccd1 net1195 sky130_fd_sc_hd__buf_4
XFILLER_0_59_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17776_ _03410_ _03437_ _03454_ _03385_ _02468_ vssd1 vssd1 vccd1 vccd1 _03455_ sky130_fd_sc_hd__a2111o_1
XANTENNA__18369__B1 net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14988_ control.body\[1011\] net151 _01549_ net2539 vssd1 vssd1 vccd1 vccd1 _00325_
+ sky130_fd_sc_hd__a22o_1
X_19515_ clknet_leaf_121_clk _00459_ net1401 vssd1 vssd1 vccd1 vccd1 control.body\[873\]
+ sky130_fd_sc_hd__dfrtp_1
X_16727_ obsg2.obstacleArray\[115\] net957 net537 vssd1 vssd1 vccd1 vccd1 _02406_
+ sky130_fd_sc_hd__and3_1
X_13939_ ag2.body\[81\] net197 _08154_ ag2.body\[73\] vssd1 vssd1 vccd1 vccd1 _00162_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_89_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10113__C1 _04551_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12653__A1 net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_62_clk_A clknet_4_13__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17041__B1 net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19446_ clknet_leaf_110_clk _00390_ net1422 vssd1 vssd1 vccd1 vccd1 control.body\[948\]
+ sky130_fd_sc_hd__dfrtp_1
X_16658_ net390 _02334_ net362 vssd1 vssd1 vccd1 vccd1 _02337_ sky130_fd_sc_hd__a21o_1
XANTENNA__17592__A1 ag2.body\[57\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_3361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17592__B2 ag2.body\[63\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18066__B _03582_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15609_ ag2.body\[458\] net123 _01620_ ag2.body\[450\] vssd1 vssd1 vccd1 vccd1 _00876_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_100_3372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_100_3383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19377_ clknet_leaf_93_clk _00321_ net1436 vssd1 vssd1 vccd1 vccd1 control.body\[1023\]
+ sky130_fd_sc_hd__dfrtp_1
X_16589_ obsg2.obstacleArray\[70\] net446 net392 _02267_ vssd1 vssd1 vccd1 vccd1 _02268_
+ sky130_fd_sc_hd__o211a_1
XANTENNA__10908__A net1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_14_clk clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_14_clk
+ sky130_fd_sc_hd__clkbuf_8
X_09130_ ag2.body\[439\] vssd1 vssd1 vccd1 vccd1 _04155_ sky130_fd_sc_hd__inv_2
XANTENNA__18136__A3 net37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13133__A_N _07486_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18328_ net902 _04519_ _04638_ _08140_ vssd1 vssd1 vccd1 vccd1 _03824_ sky130_fd_sc_hd__a31oi_2
XFILLER_0_60_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_77_clk_A clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14158__A1 net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09061_ ag2.body\[257\] vssd1 vssd1 vccd1 vccd1 _04086_ sky130_fd_sc_hd__inv_2
XANTENNA__13003__B _07639_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14158__B2 net1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18259_ net526 _03768_ vssd1 vssd1 vccd1 vccd1 _01377_ sky130_fd_sc_hd__and2_1
XANTENNA__15355__B1 _01592_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17895__A2 _03531_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_117_3880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18082__A net39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_117_3891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_120_clk_A clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_113_3755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_407 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold601 img_gen.tracker.frame\[90\] vssd1 vssd1 vccd1 vccd1 net2163 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkload40_A clknet_leaf_127_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_113_3766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14323__A1_N net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold612 obsg2.obstacleCount\[3\] vssd1 vssd1 vccd1 vccd1 net2174 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_113_3777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20221_ clknet_leaf_60_clk _01165_ net1466 vssd1 vssd1 vccd1 vccd1 ag2.body\[171\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_4_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold623 _00272_ vssd1 vssd1 vccd1 vccd1 net2185 sky130_fd_sc_hd__dlygate4sd3_1
Xhold634 control.body\[917\] vssd1 vssd1 vccd1 vccd1 net2196 sky130_fd_sc_hd__dlygate4sd3_1
Xhold645 control.body\[832\] vssd1 vssd1 vccd1 vccd1 net2207 sky130_fd_sc_hd__dlygate4sd3_1
Xhold656 control.body\[962\] vssd1 vssd1 vccd1 vccd1 net2218 sky130_fd_sc_hd__dlygate4sd3_1
Xhold667 control.body\[651\] vssd1 vssd1 vccd1 vccd1 net2229 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__17250__A1_N net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09963_ _04013_ net1163 net747 ag2.body\[87\] vssd1 vssd1 vccd1 vccd1 _04936_ sky130_fd_sc_hd__a22o_1
XANTENNA__11458__B net1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_4_Right_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold678 control.body\[729\] vssd1 vssd1 vccd1 vccd1 net2240 sky130_fd_sc_hd__dlygate4sd3_1
X_20152_ clknet_leaf_101_clk _01096_ net1452 vssd1 vssd1 vccd1 vccd1 ag2.body\[246\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__09209__A net1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_135_clk_A clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold689 control.body\[830\] vssd1 vssd1 vccd1 vccd1 net2251 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14330__A1 net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14330__B2 net1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09894_ ag2.body\[72\] net1234 vssd1 vssd1 vccd1 vccd1 _04867_ sky130_fd_sc_hd__xor2_1
X_20083_ clknet_leaf_77_clk _01027_ net1491 vssd1 vssd1 vccd1 vccd1 ag2.body\[305\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA_fanout1010_A net1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_15_clk_A clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1108_A net1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19256__CLK clknet_leaf_75_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout470_A _06648_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout568_A net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17280__B1 net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13392__C _07306_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20233__CLK clknet_leaf_66_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12644__A1 net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16476__S net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout735_A _04263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17032__B1 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1477_A net1478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1098_X net1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09879__A ag2.body\[166\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11852__C1 _06724_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_1523 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14397__B2 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_2788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout523_X net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_2799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_1642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout902_A control.body_update.curr_length\[5\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_14_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_685 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__20178__RESET_B net1461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09328_ _04337_ _04338_ vssd1 vssd1 vccd1 vccd1 _01433_ sky130_fd_sc_hd__and2b_1
XANTENNA__11604__C1 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_430 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10537__B net1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_713 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14149__A1 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09259_ sound_gen.osc1.keepCounting sound_gen.posDetector1.N\[0\] vssd1 vssd1 vccd1
+ vccd1 _04284_ sky130_fd_sc_hd__and2b_2
XANTENNA__14149__B2 net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17886__A2 _04445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12270_ _07190_ _07233_ _07239_ _07238_ vssd1 vssd1 vccd1 vccd1 _07240_ sky130_fd_sc_hd__o31a_1
XFILLER_0_121_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_1316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17099__B1 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11221_ net1099 control.body\[861\] vssd1 vssd1 vccd1 vccd1 _06194_ sky130_fd_sc_hd__xor2_1
X_20419_ clknet_leaf_33_clk _01306_ net1346 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[55\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__11649__A _06511_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14025__A net996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16846__B1 net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11152_ ag2.body\[603\] net1146 vssd1 vssd1 vccd1 vccd1 _06125_ sky130_fd_sc_hd__or2_1
XANTENNA__10272__B net1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14857__C1 _08499_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10103_ net638 _05073_ net892 vssd1 vssd1 vccd1 vccd1 _05076_ sky130_fd_sc_hd__a21o_1
X_15960_ ag2.body\[148\] net198 _01657_ ag2.body\[140\] vssd1 vssd1 vccd1 vccd1 _01190_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__14321__B2 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11083_ ag2.body\[541\] net1108 vssd1 vssd1 vccd1 vccd1 _06056_ sky130_fd_sc_hd__nand2_1
XANTENNA__16240__A _01918_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11135__A1 _04421_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14911_ control.body\[1087\] net178 _01541_ control.body\[1079\] vssd1 vssd1 vccd1
+ vccd1 _00257_ sky130_fd_sc_hd__a22o_1
X_10034_ ag2.body\[510\] net751 net1064 _04187_ vssd1 vssd1 vccd1 vccd1 _05007_ sky130_fd_sc_hd__a22o_1
X_15891_ ag2.body\[215\] net184 _01649_ ag2.body\[207\] vssd1 vssd1 vccd1 vccd1 _01129_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_21_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12883__A1 net245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_4062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17630_ _03306_ _03307_ _03308_ vssd1 vssd1 vccd1 vccd1 _03309_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_51_1880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_123_4073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14842_ _08363_ _08368_ _01509_ _01510_ _01512_ vssd1 vssd1 vccd1 vccd1 _01513_ sky130_fd_sc_hd__o2111a_1
XTAP_TAPCELL_ROW_51_1891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_32_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12199__B _07169_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16894__B net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_1460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12096__C1 net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17561_ ag2.body\[580\] net959 vssd1 vssd1 vccd1 vccd1 _03240_ sky130_fd_sc_hd__nand2_1
X_14773_ _08930_ _08931_ _08925_ vssd1 vssd1 vccd1 vccd1 _01444_ sky130_fd_sc_hd__a21o_1
X_11985_ _06952_ _06954_ _06956_ net558 vssd1 vssd1 vccd1 vccd1 _06957_ sky130_fd_sc_hd__a22o_1
XANTENNA__12767__X _07587_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16239__X _01918_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19300_ clknet_leaf_99_clk net2486 net1445 vssd1 vssd1 vccd1 vccd1 control.body\[1090\]
+ sky130_fd_sc_hd__dfrtp_1
X_16512_ obsg2.obstacleArray\[5\] _02059_ net402 _02190_ vssd1 vssd1 vccd1 vccd1 _02191_
+ sky130_fd_sc_hd__o211a_1
X_10936_ net907 _04982_ _05074_ _05798_ vssd1 vssd1 vccd1 vccd1 _05909_ sky130_fd_sc_hd__o31a_2
XANTENNA__09789__A net1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13724_ toggle1.bcd_ones\[0\] toggle1.nextBlinkToggle\[0\] toggle1.nextBlinkToggle\[1\]
+ net2233 _08054_ vssd1 vssd1 vccd1 vccd1 toggle1.nextDisplayOut\[0\] sky130_fd_sc_hd__a221o_1
X_17492_ ag2.body\[362\] net725 net718 ag2.body\[363\] vssd1 vssd1 vccd1 vccd1 _03171_
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_131_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19231_ clknet_leaf_75_clk _00175_ net1483 vssd1 vssd1 vccd1 vccd1 ag2.body\[94\]
+ sky130_fd_sc_hd__dfrtp_4
X_16443_ obsg2.obstacleArray\[64\] obsg2.obstacleArray\[65\] net456 vssd1 vssd1 vccd1
+ vccd1 _02122_ sky130_fd_sc_hd__mux2_1
X_13655_ control.divider.count\[19\] _08009_ vssd1 vssd1 vccd1 vccd1 _08011_ sky130_fd_sc_hd__and2_1
XFILLER_0_39_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10867_ ag2.body\[532\] net1132 vssd1 vssd1 vccd1 vccd1 _05840_ sky130_fd_sc_hd__or2_1
XANTENNA__18773__CLK clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_136_4456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16782__C1 net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_1529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_4467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12646__C net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_4478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19162_ clknet_leaf_52_clk _00106_ net1368 vssd1 vssd1 vccd1 vccd1 ag2.body\[25\]
+ sky130_fd_sc_hd__dfrtp_4
X_12606_ net277 _07503_ _07504_ net1735 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[59\]
+ sky130_fd_sc_hd__a22o_1
X_13586_ _03960_ control.divider.count\[4\] _07958_ vssd1 vssd1 vccd1 vccd1 _07961_
+ sky130_fd_sc_hd__or3_1
X_16374_ _01888_ _02052_ vssd1 vssd1 vccd1 vccd1 _02053_ sky130_fd_sc_hd__nor2_1
XANTENNA__16129__A2 net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10798_ ag2.body\[34\] net1175 vssd1 vssd1 vccd1 vccd1 _05771_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_45_1695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10447__B net1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11611__C_N _06497_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18113_ net300 _03627_ vssd1 vssd1 vccd1 vccd1 _03691_ sky130_fd_sc_hd__nand2_1
XFILLER_0_42_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15325_ net2568 net74 _01589_ net2222 vssd1 vssd1 vccd1 vccd1 _00623_ sky130_fd_sc_hd__a22o_1
XANTENNA__15337__B1 _01590_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_1559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12537_ net225 _07465_ vssd1 vssd1 vccd1 vccd1 _07466_ sky130_fd_sc_hd__nor2_1
X_19093_ clknet_leaf_146_clk img_gen.tracker.next_frame\[531\] net1239 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[531\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_121_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19129__CLK clknet_leaf_132_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18044_ net42 _03645_ vssd1 vssd1 vccd1 vccd1 _03646_ sky130_fd_sc_hd__nor2_1
X_12468_ _07307_ _07422_ vssd1 vssd1 vccd1 vccd1 _07423_ sky130_fd_sc_hd__nor2_2
X_15256_ net2599 net108 net50 control.body\[762\] vssd1 vssd1 vccd1 vccd1 _00564_
+ sky130_fd_sc_hd__a22o_1
X_20633__1550 vssd1 vssd1 vccd1 vccd1 _20633__1550/HI net1550 sky130_fd_sc_hd__conb_1
XFILLER_0_124_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12662__B _07444_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14207_ _08364_ _08365_ _08366_ _08367_ vssd1 vssd1 vccd1 vccd1 _08368_ sky130_fd_sc_hd__or4b_1
XANTENNA__14560__A1 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11419_ net1130 control.body\[852\] vssd1 vssd1 vccd1 vccd1 _06392_ sky130_fd_sc_hd__xor2_1
XANTENNA__14560__B2 net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17629__A2 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15187_ control.body\[836\] net102 _01572_ net2391 vssd1 vssd1 vccd1 vccd1 _00502_
+ sky130_fd_sc_hd__a22o_1
X_12399_ net1194 _07354_ _07361_ _07362_ _07298_ vssd1 vssd1 vccd1 vccd1 _07363_ sky130_fd_sc_hd__a2111o_1
XANTENNA__10463__A net1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_3084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_91_3095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16837__B1 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11374__B2 ag2.body\[478\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14138_ net989 ag2.body\[169\] vssd1 vssd1 vccd1 vccd1 _08299_ sky130_fd_sc_hd__nand2_1
XFILLER_0_26_1568 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10182__B net1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19995_ clknet_leaf_58_clk _00939_ net1472 vssd1 vssd1 vccd1 vccd1 ag2.body\[393\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_61_1459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14848__C1 _01515_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_39_1499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13115__A2 net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14069_ net1021 ag2.body\[214\] vssd1 vssd1 vccd1 vccd1 _08230_ sky130_fd_sc_hd__xor2_1
X_18946_ clknet_leaf_5_clk img_gen.tracker.next_frame\[384\] net1269 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[384\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__09971__B _04427_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_3_clk clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_3_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_94_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12874__A1 net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18877_ clknet_leaf_12_clk img_gen.tracker.next_frame\[315\] net1281 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[315\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__15057__A_N _04759_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17828_ net987 ag2.apple_cord\[1\] net224 vssd1 vssd1 vccd1 vccd1 _03491_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_106_3570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_3423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17759_ net354 _03409_ vssd1 vssd1 vccd1 vccd1 _03438_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_102_3434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11581__X _06554_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_3445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09699__A ag2.body\[67\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_1566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1122 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19429_ clknet_leaf_108_clk net2460 net1434 vssd1 vssd1 vccd1 vccd1 control.body\[963\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_110_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10197__X _05170_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout39 _03592_ vssd1 vssd1 vccd1 vccd1 net39 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10638__A net1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_119_3942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout149_A net154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13014__A net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_994 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_3953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13051__A1 net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_3964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10357__B net1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09113_ ag2.body\[383\] vssd1 vssd1 vccd1 vccd1 _04138_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_115_3817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_3828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_115_3839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12853__A _07431_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1058_A net1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09044_ ag2.body\[218\] vssd1 vssd1 vccd1 vccd1 _04069_ sky130_fd_sc_hd__inv_2
XFILLER_0_66_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_226 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold420 img_gen.tracker.frame\[533\] vssd1 vssd1 vccd1 vccd1 net1982 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold431 img_gen.tracker.frame\[361\] vssd1 vssd1 vccd1 vccd1 net1993 sky130_fd_sc_hd__dlygate4sd3_1
Xhold442 img_gen.tracker.frame\[207\] vssd1 vssd1 vccd1 vccd1 net2004 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1225_A ag2.y\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16979__B net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20204_ clknet_leaf_56_clk _01148_ net1457 vssd1 vssd1 vccd1 vccd1 ag2.body\[186\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_74_2570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold453 img_gen.tracker.frame\[480\] vssd1 vssd1 vccd1 vccd1 net2015 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__16828__B1 net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_2581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold464 img_gen.tracker.frame\[46\] vssd1 vssd1 vccd1 vccd1 net2026 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold475 img_gen.tracker.frame\[152\] vssd1 vssd1 vccd1 vccd1 net2037 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__15883__B net67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold486 img_gen.tracker.frame\[215\] vssd1 vssd1 vccd1 vccd1 net2048 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout685_A net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout900 net901 vssd1 vssd1 vccd1 vccd1 net900 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_70_2445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14303__A1 net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold497 img_gen.tracker.frame\[15\] vssd1 vssd1 vccd1 vccd1 net2059 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout911 net912 vssd1 vssd1 vccd1 vccd1 net911 sky130_fd_sc_hd__clkbuf_2
XANTENNA__13684__A _04944_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09881__B net1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14303__B2 net1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout922 net923 vssd1 vssd1 vccd1 vccd1 net922 sky130_fd_sc_hd__clkbuf_8
XANTENNA__10523__D _05495_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_2456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20135_ clknet_leaf_80_clk _01079_ net1485 vssd1 vssd1 vccd1 vccd1 ag2.body\[261\]
+ sky130_fd_sc_hd__dfrtp_4
X_09946_ net1146 control.body\[739\] vssd1 vssd1 vccd1 vccd1 _04919_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_70_2467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1013_X net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout933 net936 vssd1 vssd1 vccd1 vccd1 net933 sky130_fd_sc_hd__buf_4
XFILLER_0_42_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11117__A1 net1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout944 net945 vssd1 vssd1 vccd1 vccd1 net944 sky130_fd_sc_hd__buf_4
Xfanout955 obsg2.randCord\[5\] vssd1 vssd1 vccd1 vccd1 net955 sky130_fd_sc_hd__buf_4
Xfanout966 net967 vssd1 vssd1 vccd1 vccd1 net966 sky130_fd_sc_hd__buf_4
Xfanout977 ag2.randCord\[3\] vssd1 vssd1 vccd1 vccd1 net977 sky130_fd_sc_hd__buf_4
X_20066_ clknet_leaf_73_clk _01010_ net1501 vssd1 vssd1 vccd1 vccd1 ag2.body\[320\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA_fanout852_A net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09877_ ag2.body\[165\] net1105 vssd1 vssd1 vccd1 vccd1 _04850_ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout473_X net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout988 net995 vssd1 vssd1 vccd1 vccd1 net988 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_5_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout999 net1000 vssd1 vssd1 vccd1 vccd1 net999 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_5_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_2964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1466 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_87_2975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_79_Right_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_87_2986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17603__B net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12617__A1 net250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout640_X net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_68_2385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout738_X net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_2396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_1644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11770_ img_gen.tracker.frame\[86\] net624 net608 img_gen.tracker.frame\[89\] vssd1
+ vssd1 vccd1 vccd1 _06742_ sky130_fd_sc_hd__o22a_1
XANTENNA__13290__A1 net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10721_ _04223_ net1169 net743 ag2.body\[623\] _05688_ vssd1 vssd1 vccd1 vccd1 _05694_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_36_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11840__A2 net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15031__A2 _04607_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13440_ _07575_ net302 vssd1 vssd1 vccd1 vccd1 _07888_ sky130_fd_sc_hd__nor2_1
XANTENNA__12466__C net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10652_ ag2.body\[285\] net1115 vssd1 vssd1 vccd1 vccd1 _05625_ sky130_fd_sc_hd__xor2_1
XFILLER_0_113_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13042__A1 net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10267__B net1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_4320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13371_ net274 _07860_ _07861_ net1868 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[467\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_49_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_131_4331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10583_ _05552_ _05553_ _05554_ _05555_ vssd1 vssd1 vccd1 vccd1 _05556_ sky130_fd_sc_hd__or4_1
XFILLER_0_35_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12763__A net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_88_Right_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12322_ _07251_ _07254_ _07285_ _07287_ vssd1 vssd1 vccd1 vccd1 _07289_ sky130_fd_sc_hd__a22o_1
X_15110_ net2110 net145 _01564_ control.body\[903\] vssd1 vssd1 vccd1 vccd1 _00433_
+ sky130_fd_sc_hd__a22o_1
X_16090_ obsg2.obstacleArray\[102\] net421 vssd1 vssd1 vccd1 vccd1 _01769_ sky130_fd_sc_hd__or2_1
X_15041_ control.body\[961\] net163 _01556_ net2475 vssd1 vssd1 vccd1 vccd1 _00371_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__09549__A1 _04445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12253_ _07210_ _07222_ vssd1 vssd1 vccd1 vccd1 _07223_ sky130_fd_sc_hd__or2_1
XANTENNA__16819__B1 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11204_ _05051_ _06173_ _06174_ _06175_ _06176_ vssd1 vssd1 vccd1 vccd1 _06177_ sky130_fd_sc_hd__o2111a_1
XANTENNA__11098__B net1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12184_ net1078 ag2.apple_cord\[6\] vssd1 vssd1 vccd1 vccd1 _07156_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_129_4260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_4271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18800_ clknet_leaf_17_clk img_gen.tracker.next_frame\[238\] net1319 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[238\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__17492__B1 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11135_ _04421_ _05051_ _06106_ _06107_ vssd1 vssd1 vccd1 vccd1 _06108_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_53_1931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19780_ clknet_leaf_127_clk _00724_ net1326 vssd1 vssd1 vccd1 vccd1 ag2.body\[610\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_125_4124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16992_ _02663_ _02664_ _02665_ _02668_ vssd1 vssd1 vccd1 vccd1 _02671_ sky130_fd_sc_hd__or4b_1
XTAP_TAPCELL_ROW_53_1942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18731_ clknet_leaf_142_clk img_gen.tracker.next_frame\[169\] net1261 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[169\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_34_1352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11066_ _06028_ _06033_ _06038_ vssd1 vssd1 vccd1 vccd1 _06039_ sky130_fd_sc_hd__and3_1
X_15943_ ag2.body\[165\] net195 _01653_ ag2.body\[157\] vssd1 vssd1 vccd1 vccd1 _01175_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_34_1363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12856__A1 net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_97_Right_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_1544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10017_ ag2.body\[267\] net1164 vssd1 vssd1 vccd1 vccd1 _04990_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_30_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17244__B1 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18662_ clknet_leaf_11_clk img_gen.tracker.next_frame\[100\] net1282 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[100\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__19195__RESET_B net1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15874_ _05740_ net65 vssd1 vssd1 vccd1 vccd1 _01648_ sky130_fd_sc_hd__and2_2
X_17613_ ag2.body\[600\] net879 vssd1 vssd1 vccd1 vccd1 _03292_ sky130_fd_sc_hd__xor2_1
X_14825_ net986 _04045_ ag2.body\[158\] net802 _01490_ vssd1 vssd1 vccd1 vccd1 _01496_
+ sky130_fd_sc_hd__o221a_1
XANTENNA__12497__X _07443_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18593_ clknet_leaf_13_clk img_gen.tracker.next_frame\[31\] net1284 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[31\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_138_4518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_138_4529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17544_ _03219_ _03221_ _03222_ _03220_ vssd1 vssd1 vccd1 vccd1 _03223_ sky130_fd_sc_hd__or4b_1
XFILLER_0_118_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13281__A1 net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14756_ net1034 ag2.body\[44\] vssd1 vssd1 vccd1 vccd1 _08917_ sky130_fd_sc_hd__xor2_1
XANTENNA__12084__A2 net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11968_ img_gen.tracker.frame\[505\] net620 net599 img_gen.tracker.frame\[508\] _06939_
+ vssd1 vssd1 vccd1 vccd1 _06940_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_47_1746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13707_ track.highScore\[7\] _08035_ vssd1 vssd1 vccd1 vccd1 _08048_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_47_1768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_1442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17475_ ag2.body\[132\] net966 vssd1 vssd1 vccd1 vccd1 _03154_ sky130_fd_sc_hd__xor2_1
X_10919_ ag2.body\[460\] net1127 vssd1 vssd1 vccd1 vccd1 _05892_ sky130_fd_sc_hd__or2_1
XFILLER_0_58_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14687_ net986 _04018_ _04019_ net977 vssd1 vssd1 vccd1 vccd1 _08848_ sky130_fd_sc_hd__o22a_1
XANTENNA__11831__A2 net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11899_ net1215 net1190 img_gen.tracker.frame\[49\] vssd1 vssd1 vccd1 vccd1 _06871_
+ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_28_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19214_ clknet_leaf_58_clk _00158_ net1473 vssd1 vssd1 vccd1 vccd1 ag2.body\[77\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_89_1326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_28_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16426_ net355 _02084_ vssd1 vssd1 vccd1 vccd1 _02105_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_28_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13638_ net2043 _07997_ _07999_ vssd1 vssd1 vccd1 vccd1 control.divider.next_count\[13\]
+ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_15_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13033__A1 net238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_4_Left_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10177__B net1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16770__A2 net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19145_ clknet_leaf_47_clk _00089_ net1377 vssd1 vssd1 vccd1 vccd1 ag2.body\[9\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_97_3271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09966__B net1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_97_3282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16357_ obsg2.obstacleArray\[2\] obsg2.obstacleArray\[3\] net409 vssd1 vssd1 vccd1
+ vccd1 _02036_ sky130_fd_sc_hd__mux2_1
XANTENNA__14217__X _08378_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13569_ ssdec1.in\[1\] _07941_ _07945_ _04281_ ssdec1.in\[3\] vssd1 vssd1 vccd1 vccd1
+ net22 sky130_fd_sc_hd__o32a_1
XTAP_TAPCELL_ROW_97_3293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_3146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15308_ control.body\[735\] net77 _01586_ control.body\[727\] vssd1 vssd1 vccd1 vccd1
+ _00609_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_93_3157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19076_ clknet_leaf_29_clk img_gen.tracker.next_frame\[514\] net1334 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[514\] sky130_fd_sc_hd__dfrtp_1
X_16288_ obsg2.obstacleArray\[120\] obsg2.obstacleArray\[121\] net407 vssd1 vssd1
+ vccd1 vccd1 _01967_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_93_3168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16522__A2 _02199_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18027_ obsg2.obstacleArray\[28\] _03634_ net527 vssd1 vssd1 vccd1 vccd1 _01279_
+ sky130_fd_sc_hd__o21a_1
XANTENNA__15984__A ag2.body\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11289__A net1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14533__A1 net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_395 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15239_ net2587 net96 _01578_ control.body\[778\] vssd1 vssd1 vccd1 vccd1 _00548_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_26_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14533__B2 net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_1392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11898__A2 net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17483__B1 net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout207 net210 vssd1 vssd1 vccd1 vccd1 net207 sky130_fd_sc_hd__clkbuf_2
X_09800_ net1134 control.body\[964\] vssd1 vssd1 vccd1 vccd1 _04773_ sky130_fd_sc_hd__xor2_1
Xfanout218 net219 vssd1 vssd1 vccd1 vccd1 net218 sky130_fd_sc_hd__buf_4
X_19978_ clknet_leaf_64_clk _00922_ net1474 vssd1 vssd1 vccd1 vccd1 ag2.body\[408\]
+ sky130_fd_sc_hd__dfrtp_4
Xfanout229 net233 vssd1 vssd1 vccd1 vccd1 net229 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_61_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_108_3610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_3621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_3632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09731_ _04701_ _04702_ _04703_ _04700_ vssd1 vssd1 vccd1 vccd1 _04704_ sky130_fd_sc_hd__a211o_1
X_18929_ clknet_leaf_140_clk img_gen.tracker.next_frame\[367\] net1290 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[367\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__11736__B net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17235__B1 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_3507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09662_ net919 net922 vssd1 vssd1 vccd1 vccd1 _04635_ sky130_fd_sc_hd__xnor2_2
XANTENNA__13009__A net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1028 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16589__A2 net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17423__B net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09593_ net1179 control.body\[906\] vssd1 vssd1 vccd1 vccd1 _04566_ sky130_fd_sc_hd__xor2_1
XANTENNA__14644__A2_N net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12848__A net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout266_A net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12075__A2 net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13272__A1 net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11471__B net1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10368__A net1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16210__A1 net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1175_A net1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_59_Left_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13024__A1 net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16761__A2 net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14772__A1 net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09876__B net1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14772__B2 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout600_A net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout319_X net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_76_2632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17710__A1 net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_2643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_2654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20421__CLK clknet_leaf_37_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09027_ ag2.body\[168\] vssd1 vssd1 vccd1 vccd1 _04052_ sky130_fd_sc_hd__inv_2
XFILLER_0_108_1433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_2507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1130_X net1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_2053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_2064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_72_2529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1228_X net1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_2075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19594__CLK clknet_leaf_118_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold250 img_gen.tracker.frame\[509\] vssd1 vssd1 vccd1 vccd1 net1812 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold261 img_gen.tracker.frame\[146\] vssd1 vssd1 vccd1 vccd1 net1823 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11889__A2 net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout590_X net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16502__B _02057_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout688_X net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold272 img_gen.tracker.frame\[399\] vssd1 vssd1 vccd1 vccd1 net1834 sky130_fd_sc_hd__dlygate4sd3_1
Xhold283 img_gen.tracker.frame\[201\] vssd1 vssd1 vccd1 vccd1 net1845 sky130_fd_sc_hd__dlygate4sd3_1
Xhold294 img_gen.tracker.frame\[401\] vssd1 vssd1 vccd1 vccd1 net1856 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11927__A net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout730 net731 vssd1 vssd1 vccd1 vccd1 net730 sky130_fd_sc_hd__buf_4
Xfanout741 _04262_ vssd1 vssd1 vccd1 vccd1 net741 sky130_fd_sc_hd__clkbuf_4
X_20118_ clknet_leaf_80_clk _01062_ net1488 vssd1 vssd1 vccd1 vccd1 ag2.body\[276\]
+ sky130_fd_sc_hd__dfrtp_4
XPHY_EDGE_ROW_130_Right_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12838__A1 net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout752 _04233_ vssd1 vssd1 vccd1 vccd1 net752 sky130_fd_sc_hd__buf_4
X_09929_ _04598_ _04661_ _04783_ _04901_ vssd1 vssd1 vccd1 vccd1 _04902_ sky130_fd_sc_hd__nand4_1
XFILLER_0_102_1076 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout763 net765 vssd1 vssd1 vccd1 vccd1 net763 sky130_fd_sc_hd__buf_4
XANTENNA__10550__B net1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout855_X net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout774 _04229_ vssd1 vssd1 vccd1 vccd1 net774 sky130_fd_sc_hd__clkbuf_8
XANTENNA__17226__B1 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout785 net789 vssd1 vssd1 vccd1 vccd1 net785 sky130_fd_sc_hd__buf_4
Xfanout796 net797 vssd1 vssd1 vccd1 vccd1 net796 sky130_fd_sc_hd__buf_4
XFILLER_0_99_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20049_ clknet_leaf_74_clk _00993_ net1495 vssd1 vssd1 vccd1 vccd1 ag2.body\[351\]
+ sky130_fd_sc_hd__dfrtp_4
X_12940_ net343 _07480_ vssd1 vssd1 vccd1 vccd1 _07667_ sky130_fd_sc_hd__nor2_1
XANTENNA__11227__A1_N net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14957__B _04646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17333__B net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12871_ net678 _07636_ vssd1 vssd1 vccd1 vccd1 _07637_ sky130_fd_sc_hd__nor2_1
X_14610_ net810 ag2.body\[133\] ag2.body\[132\] net815 vssd1 vssd1 vccd1 vccd1 _08771_
+ sky130_fd_sc_hd__o2bb2a_1
X_11822_ img_gen.tracker.frame\[413\] net600 vssd1 vssd1 vccd1 vccd1 _06794_ sky130_fd_sc_hd__or2_1
XANTENNA__09467__B1 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15590_ ag2.body\[473\] net122 _01618_ ag2.body\[465\] vssd1 vssd1 vccd1 vccd1 _00859_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12066__A2 _07036_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11753_ img_gen.tracker.frame\[245\] net598 net559 vssd1 vssd1 vccd1 vccd1 _06725_
+ sky130_fd_sc_hd__o21a_1
XANTENNA__10077__B2 _05035_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14541_ net1038 ag2.body\[244\] vssd1 vssd1 vccd1 vccd1 _08702_ sky130_fd_sc_hd__nand2_1
XFILLER_0_138_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10704_ ag2.body\[21\] net1102 vssd1 vssd1 vccd1 vccd1 _05677_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_42_1610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17260_ ag2.body\[252\] net964 vssd1 vssd1 vccd1 vccd1 _02939_ sky130_fd_sc_hd__nand2_1
X_11684_ img_gen.tracker.frame\[131\] net585 net546 img_gen.tracker.frame\[128\] _06655_
+ vssd1 vssd1 vccd1 vccd1 _06656_ sky130_fd_sc_hd__o221a_1
X_14472_ net983 _04090_ ag2.body\[271\] net795 _08628_ vssd1 vssd1 vccd1 vccd1 _08633_
+ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_12_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08971__A ag2.body\[60\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16752__A2 net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16211_ net461 net496 vssd1 vssd1 vccd1 vccd1 _01890_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_23_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10635_ net1095 control.body\[669\] vssd1 vssd1 vccd1 vccd1 _05608_ sky130_fd_sc_hd__or2_1
X_13423_ net256 _07880_ _07881_ net1612 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[499\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__09786__B _04758_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_912 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17191_ ag2.body\[575\] net929 vssd1 vssd1 vccd1 vccd1 _02870_ sky130_fd_sc_hd__or2_1
XANTENNA__11601__S net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkload109 clknet_leaf_87_clk vssd1 vssd1 vccd1 vccd1 clkload109/Y sky130_fd_sc_hd__clkinv_4
X_16142_ obsg2.obstacleArray\[2\] net426 vssd1 vssd1 vccd1 vccd1 _01821_ sky130_fd_sc_hd__or2_1
X_13354_ net228 _07854_ _07855_ net1806 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[456\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_49_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10566_ _04189_ net1180 _05536_ _05537_ _05538_ vssd1 vssd1 vccd1 vccd1 _05539_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_63_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17701__A1 net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12305_ _07202_ _07228_ vssd1 vssd1 vccd1 vccd1 _07272_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_126_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13318__A2 _07807_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16073_ obsg2.obstacleArray\[124\] obsg2.obstacleArray\[125\] net424 vssd1 vssd1
+ vccd1 vccd1 _01752_ sky130_fd_sc_hd__mux2_1
X_13285_ net234 _07827_ _07828_ net1893 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[414\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_49_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10497_ _04200_ net1203 net762 ag2.body\[548\] _05465_ vssd1 vssd1 vccd1 vccd1 _05470_
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_122_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19901_ clknet_leaf_57_clk _00845_ net1464 vssd1 vssd1 vccd1 vccd1 ag2.body\[491\]
+ sky130_fd_sc_hd__dfrtp_4
X_12236_ _07197_ _07205_ vssd1 vssd1 vccd1 vccd1 _07206_ sky130_fd_sc_hd__or2_1
X_15024_ control.body\[978\] net167 _01555_ net2209 vssd1 vssd1 vccd1 vccd1 _00356_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_127_4208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09915__D_N net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12940__B _07480_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16268__A1 _01918_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16412__B net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11396__X _06369_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19832_ clknet_leaf_122_clk _00776_ net1408 vssd1 vssd1 vccd1 vccd1 ag2.body\[566\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__15309__A _04520_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12167_ img_gen.tracker.frame\[408\] net616 net545 img_gen.tracker.frame\[414\] _07138_
+ vssd1 vssd1 vccd1 vccd1 _07139_ sky130_fd_sc_hd__o221a_1
XANTENNA__14213__A net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11118_ _06066_ _06075_ _06077_ _06087_ _06090_ vssd1 vssd1 vccd1 vccd1 _06091_ sky130_fd_sc_hd__a32o_1
X_19763_ clknet_leaf_16_clk _00707_ net1322 vssd1 vssd1 vccd1 vccd1 control.body\[625\]
+ sky130_fd_sc_hd__dfrtp_1
X_16975_ ag2.body\[426\] net861 vssd1 vssd1 vccd1 vccd1 _02654_ sky130_fd_sc_hd__xnor2_1
X_12098_ img_gen.tracker.frame\[339\] net609 net554 img_gen.tracker.frame\[342\] _07069_
+ vssd1 vssd1 vccd1 vccd1 _07070_ sky130_fd_sc_hd__a221o_1
XANTENNA__10460__B net1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18714_ clknet_leaf_144_clk img_gen.tracker.next_frame\[152\] net1252 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[152\] sky130_fd_sc_hd__dfrtp_1
X_11049_ ag2.body\[386\] net1176 vssd1 vssd1 vccd1 vccd1 _06022_ sky130_fd_sc_hd__xnor2_1
X_15926_ ag2.body\[181\] net124 _01654_ ag2.body\[173\] vssd1 vssd1 vccd1 vccd1 _01159_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_127_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19694_ clknet_leaf_135_clk _00638_ net1301 vssd1 vssd1 vccd1 vccd1 control.body\[700\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput7 gpio_in[30] vssd1 vssd1 vccd1 vccd1 net7 sky130_fd_sc_hd__clkbuf_1
XANTENNA__14867__B net51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18645_ clknet_leaf_141_clk img_gen.tracker.next_frame\[83\] net1295 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[83\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_49_1808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11073__A2_N net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15857_ ag2.body\[232\] net172 _01646_ ag2.body\[224\] vssd1 vssd1 vccd1 vccd1 _01098_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12668__A _06671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1347 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14808_ net1028 ag2.body\[381\] vssd1 vssd1 vccd1 vccd1 _01479_ sky130_fd_sc_hd__xor2_1
XFILLER_0_73_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13490__C _07813_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12057__A2 net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18576_ clknet_leaf_14_clk img_gen.tracker.next_frame\[14\] net1279 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[14\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_133_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15788_ ag2.body\[298\] net208 _01639_ ag2.body\[290\] vssd1 vssd1 vccd1 vccd1 _01036_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_15_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16991__A2 net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17527_ _03201_ _03203_ _03205_ vssd1 vssd1 vccd1 vccd1 _03206_ sky130_fd_sc_hd__or3_2
XFILLER_0_34_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14739_ net1023 ag2.body\[334\] vssd1 vssd1 vccd1 vccd1 _08900_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_99_3333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11804__A2 net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_3344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_99_3355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17458_ ag2.body\[433\] net732 net703 ag2.body\[437\] vssd1 vssd1 vccd1 vccd1 _03137_
+ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__13006__A1 net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_95_3208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_3219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16743__A2 net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16409_ obsg2.obstacleArray\[99\] _02059_ net397 _02087_ vssd1 vssd1 vccd1 vccd1
+ _02088_ sky130_fd_sc_hd__o211a_1
XANTENNA__09696__B _04493_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17389_ ag2.body\[489\] net734 net728 ag2.body\[490\] vssd1 vssd1 vccd1 vccd1 _03068_
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_15_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11568__A1 _06485_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19128_ clknet_leaf_140_clk img_gen.tracker.next_frame\[566\] net1294 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[566\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13011__B net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12553__D net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19059_ clknet_leaf_9_clk img_gen.tracker.next_frame\[497\] net1274 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[497\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__18090__A net44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13946__B net67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16259__A1 net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17456__B1 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17766__A_N _02662_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14123__A net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09714_ net903 _04602_ net642 vssd1 vssd1 vccd1 vccd1 _04687_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_138_1437 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13493__A1 net250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_65_2300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09645_ _04613_ _04614_ _04615_ _04617_ vssd1 vssd1 vccd1 vccd1 _04618_ sky130_fd_sc_hd__or4_4
XANTENNA_fanout171_X net171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout550_A net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_2311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1292_A net1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout648_A net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout269_X net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12048__A2 net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09576_ _04541_ _04545_ _04547_ _04548_ vssd1 vssd1 vccd1 vccd1 _04549_ sky130_fd_sc_hd__or4_1
XANTENNA__13245__A1 net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_67_Left_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_1058 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10098__A net1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1080_X net1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout815_A net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout436_X net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1178_X net1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18834__CLK clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16734__A2 net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16056__Y _01735_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_2705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_78_2716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10385__X _05358_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout603_X net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11559__A1 net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1345_X net1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1464 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_2115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13202__A net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10420_ net1135 control.body\[1068\] vssd1 vssd1 vccd1 vccd1 _05393_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_59_2126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_2137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20598_ net1530 vssd1 vssd1 vccd1 vccd1 gpio_oeb[10] sky130_fd_sc_hd__buf_2
XFILLER_0_61_753 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10545__B net1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17695__B1 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10351_ ag2.body\[295\] net1066 vssd1 vssd1 vccd1 vccd1 _05324_ sky130_fd_sc_hd__xor2_1
XANTENNA__18984__CLK clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17609__A net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_76_Left_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13070_ net293 _07726_ _07727_ net2008 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[299\]
+ sky130_fd_sc_hd__a22o_1
X_10282_ _04982_ _05254_ _05253_ vssd1 vssd1 vccd1 vccd1 _05255_ sky130_fd_sc_hd__o21a_2
XANTENNA_fanout972_X net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17328__B net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12021_ net566 _06989_ _06992_ vssd1 vssd1 vccd1 vccd1 _06993_ sky130_fd_sc_hd__o21a_1
XFILLER_0_104_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11657__A net1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14033__A net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1503 net1504 vssd1 vssd1 vccd1 vccd1 net1503 sky130_fd_sc_hd__clkbuf_4
Xfanout1514 net1 vssd1 vssd1 vccd1 vccd1 net1514 sky130_fd_sc_hd__buf_2
XANTENNA__16659__S net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout560 net562 vssd1 vssd1 vccd1 vccd1 net560 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_1571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout571 net573 vssd1 vssd1 vccd1 vccd1 net571 sky130_fd_sc_hd__clkbuf_4
X_16760_ obsg2.obstacleArray\[23\] net503 net489 obsg2.obstacleArray\[22\] vssd1 vssd1
+ vccd1 vccd1 _02439_ sky130_fd_sc_hd__a22o_1
XFILLER_0_22_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout582 net592 vssd1 vssd1 vccd1 vccd1 net582 sky130_fd_sc_hd__buf_2
X_13972_ ag2.body\[111\] net202 _08157_ ag2.body\[103\] vssd1 vssd1 vccd1 vccd1 _00192_
+ sky130_fd_sc_hd__a22o_1
Xfanout593 net595 vssd1 vssd1 vccd1 vccd1 net593 sky130_fd_sc_hd__clkbuf_4
X_15711_ ag2.body\[375\] net141 _01629_ ag2.body\[367\] vssd1 vssd1 vccd1 vccd1 _00969_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__09414__X _04393_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10298__B2 _05270_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12923_ _07467_ net340 net335 vssd1 vssd1 vccd1 vccd1 _07659_ sky130_fd_sc_hd__and3b_1
X_16691_ _02364_ _02369_ vssd1 vssd1 vccd1 vccd1 _02370_ sky130_fd_sc_hd__nor2_1
XFILLER_0_87_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_1547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16422__A1 _02075_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_85_Left_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11392__A net1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18430_ net321 _03798_ _03797_ vssd1 vssd1 vccd1 vccd1 _03919_ sky130_fd_sc_hd__a21o_1
X_15642_ ag2.body\[424\] net126 _01623_ ag2.body\[416\] vssd1 vssd1 vccd1 vccd1 _00906_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_115_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12854_ net675 _07628_ vssd1 vssd1 vccd1 vccd1 _07629_ sky130_fd_sc_hd__nor2_1
XANTENNA__12039__A2 net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_1318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11805_ img_gen.tracker.frame\[437\] net597 net540 img_gen.tracker.frame\[440\] _06776_
+ vssd1 vssd1 vccd1 vccd1 _06777_ sky130_fd_sc_hd__o221a_1
X_18361_ _03823_ _03855_ _03821_ vssd1 vssd1 vccd1 vccd1 _03856_ sky130_fd_sc_hd__o21bai_1
X_15573_ ag2.body\[491\] net135 _01615_ ag2.body\[483\] vssd1 vssd1 vccd1 vccd1 _00845_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_68_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12785_ net316 _07595_ vssd1 vssd1 vccd1 vccd1 _07596_ sky130_fd_sc_hd__nor2_1
XFILLER_0_51_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11798__A1 net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17312_ ag2.body\[396\] net963 vssd1 vssd1 vccd1 vccd1 _02991_ sky130_fd_sc_hd__xor2_1
XANTENNA__09797__A net1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14524_ net1038 ag2.body\[252\] vssd1 vssd1 vccd1 vccd1 _08685_ sky130_fd_sc_hd__nand2_1
X_18292_ track.nextHighScore\[1\] _03787_ vssd1 vssd1 vccd1 vccd1 _03788_ sky130_fd_sc_hd__nor2_1
X_11736_ img_gen.tracker.frame\[38\] net623 vssd1 vssd1 vccd1 vccd1 _06708_ sky130_fd_sc_hd__or2_1
XANTENNA__16725__A2 net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17922__A1 net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11893__S1 net1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12935__B _07639_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14736__A1 net1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17243_ _02918_ _02919_ _02921_ vssd1 vssd1 vccd1 vccd1 _02922_ sky130_fd_sc_hd__or3b_1
X_14455_ net1027 ag2.body\[437\] vssd1 vssd1 vccd1 vccd1 _08616_ sky130_fd_sc_hd__xor2_1
XANTENNA__14736__B2 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11667_ net1144 _06636_ vssd1 vssd1 vccd1 vccd1 _06639_ sky130_fd_sc_hd__xnor2_4
XANTENNA__14208__A net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12654__C net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13406_ net672 _07874_ vssd1 vssd1 vccd1 vccd1 _07875_ sky130_fd_sc_hd__nor2_1
X_17174_ ag2.body\[457\] net870 vssd1 vssd1 vccd1 vccd1 _02853_ sky130_fd_sc_hd__nand2_1
X_10618_ ag2.body\[54\] net1074 vssd1 vssd1 vccd1 vccd1 _05591_ sky130_fd_sc_hd__xor2_1
X_14386_ net823 ag2.body\[299\] ag2.body\[303\] net795 vssd1 vssd1 vccd1 vccd1 _08547_
+ sky130_fd_sc_hd__a22o_1
X_11598_ _06485_ _06565_ _06570_ _06497_ vssd1 vssd1 vccd1 vccd1 _06571_ sky130_fd_sc_hd__a211o_1
XANTENNA__10455__B net1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16489__A1 net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_94_Left_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16125_ obsg2.obstacleArray\[88\] net428 net375 _01803_ vssd1 vssd1 vccd1 vccd1 _01804_
+ sky130_fd_sc_hd__o211a_1
X_13337_ net332 _07508_ _07813_ vssd1 vssd1 vccd1 vccd1 _07848_ sky130_fd_sc_hd__and3_1
XFILLER_0_24_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10549_ ag2.body\[227\] net1159 vssd1 vssd1 vccd1 vccd1 _05522_ sky130_fd_sc_hd__or2_1
XFILLER_0_11_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16056_ net536 _01725_ _01733_ vssd1 vssd1 vccd1 vccd1 _01735_ sky130_fd_sc_hd__o21ai_2
X_13268_ net310 _07457_ vssd1 vssd1 vccd1 vccd1 _07821_ sky130_fd_sc_hd__nor2_1
XFILLER_0_62_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16142__B net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17438__B1 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15007_ control.body\[996\] net152 _01552_ net2344 vssd1 vssd1 vccd1 vccd1 _00342_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_122_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12219_ img_gen.updater.commands.count\[1\] img_gen.updater.commands.count\[0\] vssd1
+ vssd1 vccd1 vccd1 _07189_ sky130_fd_sc_hd__or2_1
XFILLER_0_62_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_88_3001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13199_ img_gen.tracker.frame\[367\] net658 vssd1 vssd1 vccd1 vccd1 _07790_ sky130_fd_sc_hd__and2_1
XANTENNA__13485__C net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10471__A net1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_3012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19815_ clknet_leaf_89_clk _00759_ net1410 vssd1 vssd1 vccd1 vccd1 ag2.body\[581\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__10190__B net1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_1447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16958_ ag2.body\[291\] net854 vssd1 vssd1 vccd1 vccd1 _02637_ sky130_fd_sc_hd__xor2_1
X_19746_ clknet_leaf_129_clk _00690_ net1327 vssd1 vssd1 vccd1 vccd1 control.body\[640\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__18069__B _03586_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15909_ ag2.body\[199\] net129 _01651_ ag2.body\[191\] vssd1 vssd1 vccd1 vccd1 _01145_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_79_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19677_ clknet_leaf_136_clk _00621_ net1384 vssd1 vssd1 vccd1 vccd1 control.body\[715\]
+ sky130_fd_sc_hd__dfrtp_1
X_16889_ _04068_ net863 net706 ag2.body\[213\] _02567_ vssd1 vssd1 vccd1 vccd1 _02568_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_36_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09430_ net927 net1127 vssd1 vssd1 vccd1 vccd1 _04403_ sky130_fd_sc_hd__nand2_1
XFILLER_0_56_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18628_ clknet_leaf_0_clk img_gen.tracker.next_frame\[66\] net1242 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[66\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_1481 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13227__A1 net239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10189__Y _05162_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09361_ sound_gen.osc1.stayCount\[9\] _04354_ vssd1 vssd1 vccd1 vccd1 _04363_ sky130_fd_sc_hd__and2_1
XFILLER_0_133_1356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18559_ clknet_leaf_132_clk _00085_ net1303 vssd1 vssd1 vccd1 vccd1 ag2.x\[1\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__18166__A1 net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18085__A net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16177__B1 net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09292_ sound_gen.osc1.count\[1\] sound_gen.osc1.count\[0\] vssd1 vssd1 vccd1 vccd1
+ _04312_ sky130_fd_sc_hd__or2_1
XFILLER_0_30_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12450__A2 net1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16716__A2 net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_12 _03446_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_23 control.button3.Q\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20521_ clknet_leaf_93_clk track.nextCurrScore\[3\] net1413 vssd1 vssd1 vccd1 vccd1
+ control.body_update.curr_length\[3\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_34 _06676_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout131_A net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14118__A net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout229_A net233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16036__C net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09994__X _04967_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20452_ clknet_leaf_38_clk _01339_ net1354 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[88\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_103_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18469__A2 net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_455 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17677__B1 net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20383_ clknet_leaf_40_clk _01270_ net1374 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[19\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__13950__A2 net191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1040_A net1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_1572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1138_A net1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13676__B _07181_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17148__B net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19227__RESET_B net1482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17429__B1 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout598_A _06476_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10516__A2 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16987__B net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout386_X net386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout765_A net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15236__X _01578_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout932_A net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout553_X net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17601__B1 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09628_ _04236_ net901 _04239_ vssd1 vssd1 vccd1 vccd1 _04601_ sky130_fd_sc_hd__or3_2
XANTENNA_fanout44_A net46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19782__CLK clknet_leaf_127_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout720_X net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_7_0_clk_X clknet_3_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09559_ net1096 control.body\[725\] vssd1 vssd1 vccd1 vccd1 _04532_ sky130_fd_sc_hd__xor2_1
XANTENNA__17611__B net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout818_X net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12570_ net245 _07484_ _07485_ net1908 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[42\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__16168__B1 net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16707__A2 net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12441__A2 net1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11521_ _06490_ _06493_ vssd1 vssd1 vccd1 vccd1 _06494_ sky130_fd_sc_hd__xnor2_1
XANTENNA__15915__B1 _01652_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14240_ net836 ag2.body\[481\] ag2.body\[486\] net799 vssd1 vssd1 vccd1 vccd1 _08401_
+ sky130_fd_sc_hd__o22a_1
X_11452_ _06414_ _06415_ _06423_ _06424_ vssd1 vssd1 vccd1 vccd1 _06425_ sky130_fd_sc_hd__or4_1
XFILLER_0_123_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14194__A2 ag2.body\[161\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10275__B net1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10204__A1 _05162_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10403_ net1160 control.body\[1075\] vssd1 vssd1 vccd1 vccd1 _05376_ sky130_fd_sc_hd__xor2_1
XANTENNA__10204__B2 _05151_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14171_ net988 _04063_ _04065_ net1029 _08331_ vssd1 vssd1 vccd1 vccd1 _08332_ sky130_fd_sc_hd__a221o_1
XFILLER_0_81_1204 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11383_ net1146 control.body\[643\] vssd1 vssd1 vccd1 vccd1 _06356_ sky130_fd_sc_hd__or2_1
XFILLER_0_127_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19162__CLK clknet_leaf_52_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13122_ net683 _07752_ vssd1 vssd1 vccd1 vccd1 _07753_ sky130_fd_sc_hd__nor2_1
X_10334_ ag2.body\[523\] net1159 vssd1 vssd1 vccd1 vccd1 _05307_ sky130_fd_sc_hd__or2_1
X_17930_ net380 net493 _03561_ vssd1 vssd1 vccd1 vccd1 _03562_ sky130_fd_sc_hd__and3_1
XFILLER_0_24_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11387__A net1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13053_ net338 _07421_ net329 vssd1 vssd1 vccd1 vccd1 _07720_ sky130_fd_sc_hd__and3_2
X_10265_ net907 net923 vssd1 vssd1 vccd1 vccd1 _05238_ sky130_fd_sc_hd__nand2_4
XFILLER_0_123_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12052__S1 net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1300 net1302 vssd1 vssd1 vccd1 vccd1 net1300 sky130_fd_sc_hd__clkbuf_4
X_12004_ net558 _06975_ _06973_ vssd1 vssd1 vccd1 vccd1 _06976_ sky130_fd_sc_hd__a21o_1
Xfanout1311 net1333 vssd1 vssd1 vccd1 vccd1 net1311 sky130_fd_sc_hd__buf_2
XFILLER_0_24_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17861_ _04279_ _03499_ _04278_ vssd1 vssd1 vccd1 vccd1 _03512_ sky130_fd_sc_hd__o21ai_1
X_10196_ ag2.body\[118\] net1090 vssd1 vssd1 vccd1 vccd1 _05169_ sky130_fd_sc_hd__xor2_1
Xfanout1322 net1323 vssd1 vssd1 vccd1 vccd1 net1322 sky130_fd_sc_hd__clkbuf_2
XANTENNA__14698__A net1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1333 net1505 vssd1 vssd1 vccd1 vccd1 net1333 sky130_fd_sc_hd__clkbuf_8
Xfanout1344 net1345 vssd1 vssd1 vccd1 vccd1 net1344 sky130_fd_sc_hd__clkbuf_2
Xfanout1355 net1356 vssd1 vssd1 vccd1 vccd1 net1355 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_108_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16812_ _02484_ _02486_ _02489_ _02490_ vssd1 vssd1 vccd1 vccd1 _02491_ sky130_fd_sc_hd__or4_2
X_19600_ clknet_leaf_119_clk _00544_ net1390 vssd1 vssd1 vccd1 vccd1 control.body\[798\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1366 net1370 vssd1 vssd1 vccd1 vccd1 net1366 sky130_fd_sc_hd__buf_2
X_17792_ _03466_ _03467_ vssd1 vssd1 vccd1 vccd1 _01212_ sky130_fd_sc_hd__nor2_1
XANTENNA__13457__A1 net235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1377 net1383 vssd1 vssd1 vccd1 vccd1 net1377 sky130_fd_sc_hd__clkbuf_4
Xfanout390 net393 vssd1 vssd1 vccd1 vccd1 net390 sky130_fd_sc_hd__clkbuf_4
Xfanout1388 net1389 vssd1 vssd1 vccd1 vccd1 net1388 sky130_fd_sc_hd__clkbuf_4
Xfanout1399 net1400 vssd1 vssd1 vccd1 vccd1 net1399 sky130_fd_sc_hd__clkbuf_4
X_19531_ clknet_leaf_118_clk _00475_ net1394 vssd1 vssd1 vccd1 vccd1 control.body\[857\]
+ sky130_fd_sc_hd__dfrtp_1
X_16743_ obsg2.obstacleArray\[32\] net490 net481 obsg2.obstacleArray\[33\] _02421_
+ vssd1 vssd1 vccd1 vccd1 _02422_ sky130_fd_sc_hd__a221o_1
XFILLER_0_17_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13955_ _04421_ net634 net67 vssd1 vssd1 vccd1 vccd1 _08156_ sky130_fd_sc_hd__o21a_2
XANTENNA__17199__A2 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11563__S0 net1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkload7_A clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19462_ clknet_leaf_110_clk _00406_ net1418 vssd1 vssd1 vccd1 vccd1 control.body\[932\]
+ sky130_fd_sc_hd__dfrtp_1
X_12906_ _07652_ net268 _07650_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[211\]
+ sky130_fd_sc_hd__mux2_1
X_16674_ obsg2.obstacleArray\[24\] obsg2.obstacleArray\[25\] net447 vssd1 vssd1 vccd1
+ vccd1 _02353_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14406__B1 net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13886_ ag2.body\[34\] net119 _08148_ ag2.body\[26\] vssd1 vssd1 vccd1 vccd1 _00115_
+ sky130_fd_sc_hd__a22o_1
XANTENNA_output25_A net25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18413_ _03823_ _03901_ _03902_ vssd1 vssd1 vccd1 vccd1 _03903_ sky130_fd_sc_hd__o21a_1
XFILLER_0_134_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15625_ ag2.body\[441\] net125 _01621_ ag2.body\[433\] vssd1 vssd1 vccd1 vccd1 _00891_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_75_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_1104 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1620 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17521__B net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12837_ net239 _07619_ _07620_ net1835 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[174\]
+ sky130_fd_sc_hd__a22o_1
X_19393_ clknet_leaf_102_clk _00337_ net1428 vssd1 vssd1 vccd1 vccd1 control.body\[1007\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_68_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11850__A net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18344_ _03837_ _03839_ _03823_ vssd1 vssd1 vccd1 vccd1 _03840_ sky130_fd_sc_hd__a21oi_1
X_15556_ ag2.body\[509\] net187 _01612_ ag2.body\[501\] vssd1 vssd1 vccd1 vccd1 _00831_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_31_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12768_ net305 _07587_ vssd1 vssd1 vccd1 vccd1 _07588_ sky130_fd_sc_hd__nor2_1
XANTENNA__10737__Y _05710_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14507_ net1016 ag2.body\[182\] vssd1 vssd1 vccd1 vccd1 _08668_ sky130_fd_sc_hd__xor2_1
XANTENNA__14709__A1 net1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18275_ net517 _03776_ vssd1 vssd1 vccd1 vccd1 _01385_ sky130_fd_sc_hd__nor2_1
X_11719_ _06641_ _06644_ _06671_ net466 vssd1 vssd1 vccd1 vccd1 _06691_ sky130_fd_sc_hd__a31o_1
XANTENNA__14709__B2 net1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10466__A net1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15487_ ag2.body\[575\] net109 _01605_ ag2.body\[567\] vssd1 vssd1 vccd1 vccd1 _00769_
+ sky130_fd_sc_hd__a22o_1
X_12699_ net237 net311 _07553_ _07554_ net1634 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[102\]
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_25_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_928 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17226_ _04103_ net887 net720 ag2.body\[315\] vssd1 vssd1 vccd1 vccd1 _02905_ sky130_fd_sc_hd__o22a_1
X_14438_ net1026 ag2.body\[21\] vssd1 vssd1 vccd1 vccd1 _08599_ sky130_fd_sc_hd__xor2_1
XANTENNA__19505__CLK clknet_leaf_113_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_614 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15976__B net56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10185__B net1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09974__B _04695_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17157_ ag2.body\[610\] net722 net928 _04221_ vssd1 vssd1 vccd1 vccd1 _02836_ sky130_fd_sc_hd__o22a_1
XANTENNA__12681__A _06671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold805 control.body\[867\] vssd1 vssd1 vccd1 vccd1 net2367 sky130_fd_sc_hd__dlygate4sd3_1
X_14369_ _08523_ _08524_ _08525_ _08527_ vssd1 vssd1 vccd1 vccd1 _08530_ sky130_fd_sc_hd__and4_1
XFILLER_0_106_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold816 control.body\[638\] vssd1 vssd1 vccd1 vccd1 net2378 sky130_fd_sc_hd__dlygate4sd3_1
X_16108_ obsg2.obstacleArray\[86\] net428 vssd1 vssd1 vccd1 vccd1 _01787_ sky130_fd_sc_hd__or2_1
Xhold827 _00414_ vssd1 vssd1 vccd1 vccd1 net2389 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold838 control.body\[699\] vssd1 vssd1 vccd1 vccd1 net2400 sky130_fd_sc_hd__dlygate4sd3_1
X_17088_ _02763_ _02764_ _02766_ vssd1 vssd1 vccd1 vccd1 _02767_ sky130_fd_sc_hd__nand3b_1
Xhold849 control.body\[864\] vssd1 vssd1 vccd1 vccd1 net2411 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10913__B net1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11297__A net1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20296__RESET_B net1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16039_ _01716_ _01717_ vssd1 vssd1 vccd1 vccd1 _01718_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_111_3694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09990__A net1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_1480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16600__B net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13448__A1 net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19729_ clknet_leaf_132_clk _00673_ net1304 vssd1 vssd1 vccd1 vccd1 control.body\[671\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_74_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09989__X _04962_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09413_ _04392_ vssd1 vssd1 vccd1 vccd1 img_gen.updater.update.wr sky130_fd_sc_hd__inv_2
XFILLER_0_88_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout346_A _01732_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1088_A net1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09344_ sound_gen.osc1.stayCount\[12\] sound_gen.osc1.stayCount\[11\] sound_gen.osc1.stayCount\[8\]
+ vssd1 vssd1 vccd1 vccd1 _04348_ sky130_fd_sc_hd__and3_1
XFILLER_0_47_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12575__B net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11631__B1 net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09275_ sound_gen.osc1.stayCount\[20\] _04287_ net535 sound_gen.osc1.stayCount\[19\]
+ vssd1 vssd1 vccd1 vccd1 _04298_ sky130_fd_sc_hd__o22a_1
XANTENNA__16762__S net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout513_A net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19185__CLK clknet_leaf_53_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_986 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20504_ clknet_leaf_130_clk coll.nextGoodColl net1317 vssd1 vssd1 vccd1 vccd1 ag2.goodColl
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_133_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20435_ clknet_leaf_23_clk _01322_ net1359 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[71\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_71_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout301_X net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10737__A2 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20366_ clknet_leaf_21_clk _01253_ net1360 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[2\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__11919__B net1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10820__A1_N net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout882_A net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1210_X net1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20297_ clknet_leaf_36_clk control.divider.next_count\[18\] net1347 vssd1 vssd1 vccd1
+ vccd1 control.divider.count\[18\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_41_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11000__A _05253_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10050_ _04931_ _04962_ _04997_ _05022_ vssd1 vssd1 vccd1 vccd1 _05023_ sky130_fd_sc_hd__and4_1
XANTENNA_fanout670_X net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout768_X net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15407__A _04574_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13439__A1 net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14311__A net1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11654__B net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout935_X net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18378__B2 net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13740_ net320 vssd1 vssd1 vccd1 vccd1 _08061_ sky130_fd_sc_hd__inv_2
X_10952_ ag2.body\[170\] net1176 vssd1 vssd1 vccd1 vccd1 _05925_ sky130_fd_sc_hd__xor2_1
XANTENNA__16928__A2 net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17341__B net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13671_ net922 track.current_collision vssd1 vssd1 vccd1 vccd1 _08020_ sky130_fd_sc_hd__nand2_1
XANTENNA__10838__X _05811_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10883_ net896 net905 _04471_ net636 vssd1 vssd1 vccd1 vccd1 _05856_ sky130_fd_sc_hd__a31oi_4
XANTENNA__16238__A net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15410_ net2289 net81 _01597_ control.body\[626\] vssd1 vssd1 vccd1 vccd1 _00700_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_109_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12622_ net666 _07513_ vssd1 vssd1 vccd1 vccd1 _07514_ sky130_fd_sc_hd__nor2_1
X_16390_ obsg2.obstacleArray\[120\] obsg2.obstacleArray\[121\] net455 vssd1 vssd1
+ vccd1 vccd1 _02069_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15341_ net2307 net71 _01590_ net2546 vssd1 vssd1 vccd1 vccd1 _00638_ sky130_fd_sc_hd__a22o_1
XANTENNA__11622__B1 _06485_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12553_ net618 net439 net469 net561 vssd1 vssd1 vccd1 vccd1 _07475_ sky130_fd_sc_hd__or4_1
XANTENNA__16672__S net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18060_ net352 _03577_ vssd1 vssd1 vccd1 vccd1 _03656_ sky130_fd_sc_hd__nand2_1
XFILLER_0_80_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11504_ net773 net605 vssd1 vssd1 vccd1 vccd1 _06477_ sky130_fd_sc_hd__nand2_1
XANTENNA__20505__CLK clknet_leaf_132_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15272_ net2162 net108 _01582_ net2238 vssd1 vssd1 vccd1 vccd1 _00577_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_134_4395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12484_ net311 _07435_ vssd1 vssd1 vccd1 vccd1 _07436_ sky130_fd_sc_hd__and2_1
XANTENNA__18552__CLK clknet_leaf_37_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17011_ ag2.body\[496\] net886 vssd1 vssd1 vccd1 vccd1 _02690_ sky130_fd_sc_hd__xor2_1
XFILLER_0_22_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14223_ net793 ag2.body\[399\] ag2.body\[393\] net833 vssd1 vssd1 vccd1 vccd1 _08384_
+ sky130_fd_sc_hd__a2bb2o_1
X_11435_ ag2.body\[396\] net1139 vssd1 vssd1 vccd1 vccd1 _06408_ sky130_fd_sc_hd__xor2_1
XFILLER_0_110_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17105__A2 net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11366_ net1099 control.body\[813\] vssd1 vssd1 vccd1 vccd1 _06339_ sky130_fd_sc_hd__nand2_1
X_14154_ _08309_ _08311_ _08313_ _08314_ vssd1 vssd1 vccd1 vccd1 _08315_ sky130_fd_sc_hd__or4b_4
XFILLER_0_123_1311 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10733__B net1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1491 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10317_ ag2.body\[612\] net1120 vssd1 vssd1 vccd1 vccd1 _05290_ sky130_fd_sc_hd__or2_1
X_13105_ net344 _07575_ vssd1 vssd1 vccd1 vccd1 _07745_ sky130_fd_sc_hd__nor2_1
XFILLER_0_131_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11548__C _06503_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11297_ net1072 control.body\[686\] vssd1 vssd1 vccd1 vccd1 _06270_ sky130_fd_sc_hd__xor2_1
X_18962_ clknet_leaf_7_clk img_gen.tracker.next_frame\[400\] net1266 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[400\] sky130_fd_sc_hd__dfrtp_1
X_14085_ _08238_ _08239_ _08242_ _08245_ vssd1 vssd1 vccd1 vccd1 _08246_ sky130_fd_sc_hd__or4_1
XFILLER_0_123_1366 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13678__B2 net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10248_ _05208_ _05209_ _05218_ _05219_ _05220_ vssd1 vssd1 vccd1 vccd1 _05221_ sky130_fd_sc_hd__a221o_1
X_17913_ _01818_ _03536_ vssd1 vssd1 vccd1 vccd1 _03548_ sky130_fd_sc_hd__nor2_1
X_13036_ net283 _07710_ _07711_ net1677 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[281\]
+ sky130_fd_sc_hd__a22o_1
X_18893_ clknet_leaf_26_clk img_gen.tracker.next_frame\[331\] net1342 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[331\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1130 net1131 vssd1 vssd1 vccd1 vccd1 net1130 sky130_fd_sc_hd__clkbuf_4
Xfanout1141 net1142 vssd1 vssd1 vccd1 vccd1 net1141 sky130_fd_sc_hd__buf_4
XFILLER_0_119_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17844_ _04278_ _04279_ _03499_ vssd1 vssd1 vccd1 vccd1 _03500_ sky130_fd_sc_hd__or3_1
XFILLER_0_121_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10179_ _04427_ net638 net642 vssd1 vssd1 vccd1 vccd1 _05152_ sky130_fd_sc_hd__a21oi_2
Xfanout1152 net1153 vssd1 vssd1 vccd1 vccd1 net1152 sky130_fd_sc_hd__buf_4
XANTENNA__14221__A net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1163 net1166 vssd1 vssd1 vccd1 vccd1 net1163 sky130_fd_sc_hd__clkbuf_4
Xfanout1174 net1178 vssd1 vssd1 vccd1 vccd1 net1174 sky130_fd_sc_hd__clkbuf_8
Xfanout1185 net1188 vssd1 vssd1 vccd1 vccd1 net1185 sky130_fd_sc_hd__buf_4
XFILLER_0_94_1439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17775_ _03029_ _03057_ _03439_ _03453_ vssd1 vssd1 vccd1 vccd1 _03454_ sky130_fd_sc_hd__or4b_1
Xfanout1196 net1200 vssd1 vssd1 vccd1 vccd1 net1196 sky130_fd_sc_hd__clkbuf_4
X_14987_ control.body\[1010\] net154 _01549_ net2516 vssd1 vssd1 vccd1 vccd1 _00324_
+ sky130_fd_sc_hd__a22o_1
X_16726_ obsg2.obstacleArray\[118\] net487 net483 obsg2.obstacleArray\[117\] net495
+ vssd1 vssd1 vccd1 vccd1 _02405_ sky130_fd_sc_hd__a221o_1
X_19514_ clknet_leaf_121_clk _00458_ net1401 vssd1 vssd1 vccd1 vccd1 control.body\[872\]
+ sky130_fd_sc_hd__dfrtp_1
X_13938_ ag2.body\[80\] net197 _08154_ ag2.body\[72\] vssd1 vssd1 vccd1 vccd1 _00161_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__16919__A2 net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_4_8__f_clk_X clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19445_ clknet_leaf_110_clk _00389_ net1422 vssd1 vssd1 vccd1 vccd1 control.body\[947\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_134_1451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16657_ obsg2.obstacleArray\[8\] net443 net394 _02335_ vssd1 vssd1 vccd1 vccd1 _02336_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_48_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11861__B1 net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17251__B net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13869_ net742 _08030_ _08142_ vssd1 vssd1 vccd1 vccd1 _08143_ sky130_fd_sc_hd__and3_1
XANTENNA__12676__A net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17592__A2 net731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15608_ ag2.body\[457\] net124 _01620_ ag2.body\[449\] vssd1 vssd1 vccd1 vccd1 _00875_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_100_3362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_3373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19376_ clknet_leaf_93_clk _00320_ net1437 vssd1 vssd1 vccd1 vccd1 control.body\[1022\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_100_3384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16588_ obsg2.obstacleArray\[71\] net451 vssd1 vssd1 vccd1 vccd1 _02267_ sky130_fd_sc_hd__or2_1
XFILLER_0_57_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18327_ net893 _08031_ _03822_ _08140_ vssd1 vssd1 vccd1 vccd1 _03823_ sky130_fd_sc_hd__o31a_2
XFILLER_0_45_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15539_ ag2.body\[525\] net161 _01611_ ag2.body\[517\] vssd1 vssd1 vccd1 vccd1 _00815_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_71_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09060_ ag2.body\[256\] vssd1 vssd1 vccd1 vccd1 _04085_ sky130_fd_sc_hd__inv_2
X_18258_ net353 _03638_ net37 obsg2.obstacleArray\[126\] vssd1 vssd1 vccd1 vccd1 _03768_
+ sky130_fd_sc_hd__a31o_1
XANTENNA__09985__A net1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_117_3881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_117_3892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17209_ ag2.body\[52\] net959 vssd1 vssd1 vccd1 vccd1 _02888_ sky130_fd_sc_hd__or2_1
XANTENNA__13905__A2 net90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18189_ obsg2.obstacleArray\[91\] _03733_ net531 vssd1 vssd1 vccd1 vccd1 _01342_
+ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_113_3756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold602 control.body\[906\] vssd1 vssd1 vccd1 vccd1 net2164 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10719__A2 net1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20220_ clknet_leaf_61_clk _01164_ net1382 vssd1 vssd1 vccd1 vccd1 ag2.body\[170\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_113_3767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold613 obsg2.obstacleCount\[2\] vssd1 vssd1 vccd1 vccd1 net2175 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_113_3778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold624 control.body\[1091\] vssd1 vssd1 vccd1 vccd1 net2186 sky130_fd_sc_hd__dlygate4sd3_1
Xhold635 _00415_ vssd1 vssd1 vccd1 vccd1 net2197 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11739__B net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold646 control.body\[807\] vssd1 vssd1 vccd1 vccd1 net2208 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10643__B _04791_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15658__A2 net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold657 _00364_ vssd1 vssd1 vccd1 vccd1 net2219 sky130_fd_sc_hd__dlygate4sd3_1
Xhold668 control.body\[694\] vssd1 vssd1 vccd1 vccd1 net2230 sky130_fd_sc_hd__dlygate4sd3_1
X_20151_ clknet_leaf_98_clk _01095_ net1452 vssd1 vssd1 vccd1 vccd1 ag2.body\[245\]
+ sky130_fd_sc_hd__dfrtp_4
X_09962_ ag2.body\[86\] net1088 vssd1 vssd1 vccd1 vccd1 _04935_ sky130_fd_sc_hd__or2_1
Xhold679 control.body\[670\] vssd1 vssd1 vccd1 vccd1 net2241 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17232__A2_N net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20082_ clknet_leaf_77_clk _01026_ net1490 vssd1 vssd1 vccd1 vccd1 ag2.body\[304\]
+ sky130_fd_sc_hd__dfrtp_4
X_09893_ ag2.body\[76\] net1139 vssd1 vssd1 vccd1 vccd1 _04866_ sky130_fd_sc_hd__or2_1
XANTENNA__16068__C1 net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16607__A1 net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10352__B1 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1003_A net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14618__B1 ag2.body\[62\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16083__A2 net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11474__B net1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17161__B net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09879__B net1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout630_A _06473_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16058__A net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12586__A net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout349_X net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout728_A net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_40_Left_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_1535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_1670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_81_2789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_826 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09327_ sound_gen.dac1.dacCount\[5\] _04336_ sound_gen.dac1.dacCount\[6\] vssd1 vssd1
+ vccd1 vccd1 _04338_ sky130_fd_sc_hd__a21o_1
XFILLER_0_34_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_62_2199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16492__S net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_1529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09258_ track.highScore\[5\] vssd1 vssd1 vccd1 vccd1 _04283_ sky130_fd_sc_hd__inv_2
XFILLER_0_133_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17886__A3 _03523_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16064__Y _01743_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15897__A2 net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09189_ ag2.body\[586\] vssd1 vssd1 vccd1 vccd1 _04214_ sky130_fd_sc_hd__inv_2
XFILLER_0_62_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11220_ _06180_ _06182_ _06187_ _06192_ vssd1 vssd1 vccd1 vccd1 _06193_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_43_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20418_ clknet_leaf_34_clk _01305_ net1346 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[54\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_102_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout885_X net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15649__A2 net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11151_ ag2.body\[603\] net1146 vssd1 vssd1 vccd1 vccd1 _06124_ sky130_fd_sc_hd__nand2_1
XFILLER_0_124_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20349_ clknet_leaf_139_clk _01240_ net1292 vssd1 vssd1 vccd1 vccd1 img_gen.updater.commands.rR1.rainbowRNG\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_31_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14857__B1 _08437_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_997 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10102_ net638 _05073_ vssd1 vssd1 vccd1 vccd1 _05075_ sky130_fd_sc_hd__nand2_2
XANTENNA__18048__B1 net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11082_ ag2.body\[541\] net1108 vssd1 vssd1 vccd1 vccd1 _06055_ sky130_fd_sc_hd__or2_1
XANTENNA__17336__B net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10840__Y _05813_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19200__CLK clknet_leaf_53_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10033_ ag2.body\[505\] net1210 vssd1 vssd1 vccd1 vccd1 _05006_ sky130_fd_sc_hd__or2_1
XANTENNA__11665__A net1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14910_ net2573 net177 _01541_ control.body\[1078\] vssd1 vssd1 vccd1 vccd1 _00256_
+ sky130_fd_sc_hd__a22o_1
X_15890_ ag2.body\[214\] net184 _01649_ ag2.body\[206\] vssd1 vssd1 vccd1 vccd1 _01128_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__10343__B1 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14841_ _08932_ _01445_ _01511_ _08830_ vssd1 vssd1 vccd1 vccd1 _01512_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_51_1881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_51_1892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_32_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17560_ _03231_ _03232_ _03234_ _03238_ vssd1 vssd1 vccd1 vccd1 _03239_ sky130_fd_sc_hd__or4_1
X_14772_ net823 ag2.body\[99\] ag2.body\[101\] net808 _08929_ vssd1 vssd1 vccd1 vccd1
+ _01443_ sky130_fd_sc_hd__a221o_1
XANTENNA__08974__A ag2.body\[65\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11984_ img_gen.tracker.frame\[529\] net613 net579 img_gen.tracker.frame\[538\] _06955_
+ vssd1 vssd1 vccd1 vccd1 _06956_ sky130_fd_sc_hd__o221a_1
XANTENNA__19350__CLK clknet_leaf_102_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16511_ obsg2.obstacleArray\[4\] net457 vssd1 vssd1 vccd1 vccd1 _02190_ sky130_fd_sc_hd__or2_1
X_13723_ net26 toggle1.bcd_hundreds\[0\] vssd1 vssd1 vccd1 vccd1 _08054_ sky130_fd_sc_hd__and2_1
XFILLER_0_58_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17491_ ag2.body\[363\] net718 net706 ag2.body\[365\] vssd1 vssd1 vccd1 vccd1 _03170_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_105_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10935_ _05885_ _05890_ _05897_ _05907_ _04646_ vssd1 vssd1 vccd1 vccd1 _05908_ sky130_fd_sc_hd__a32o_1
XANTENNA__11843__B1 net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18918__CLK clknet_leaf_142_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12496__A net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17574__A2 net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19230_ clknet_leaf_75_clk _00174_ net1482 vssd1 vssd1 vccd1 vccd1 ag2.body\[93\]
+ sky130_fd_sc_hd__dfrtp_4
X_16442_ obsg2.obstacleArray\[66\] obsg2.obstacleArray\[67\] net456 vssd1 vssd1 vccd1
+ vccd1 _02121_ sky130_fd_sc_hd__mux2_1
X_13654_ control.divider.count\[18\] _08008_ _08010_ net221 vssd1 vssd1 vccd1 vccd1
+ control.divider.next_count\[18\] sky130_fd_sc_hd__o211a_1
X_10866_ _05496_ _05619_ _05725_ _05838_ vssd1 vssd1 vccd1 vccd1 _05839_ sky130_fd_sc_hd__or4b_1
XTAP_TAPCELL_ROW_136_4457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12399__A1 net1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_136_4468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19161_ clknet_leaf_52_clk _00105_ net1363 vssd1 vssd1 vccd1 vccd1 ag2.body\[24\]
+ sky130_fd_sc_hd__dfrtp_4
X_12605_ net252 _07503_ _07504_ net1764 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[58\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_27_826 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_136_4479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16373_ net956 net948 net939 net930 vssd1 vssd1 vccd1 vccd1 _02052_ sky130_fd_sc_hd__and4b_1
XANTENNA__12646__D net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13585_ control.divider.count\[7\] _07959_ vssd1 vssd1 vccd1 vccd1 _07960_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_45_1685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_563 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10797_ _05766_ _05767_ _05768_ _05769_ vssd1 vssd1 vccd1 vccd1 _05770_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_45_1696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18112_ obsg2.obstacleArray\[57\] _03690_ net525 vssd1 vssd1 vccd1 vccd1 _01308_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_121_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15324_ net2576 net74 _01589_ net2247 vssd1 vssd1 vccd1 vccd1 _00622_ sky130_fd_sc_hd__a22o_1
XFILLER_0_26_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19092_ clknet_leaf_146_clk img_gen.tracker.next_frame\[530\] net1239 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[530\] sky130_fd_sc_hd__dfrtp_1
X_12536_ net2081 net649 _07465_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[28\]
+ sky130_fd_sc_hd__and3_1
XFILLER_0_13_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12943__B net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18043_ net301 _03554_ vssd1 vssd1 vccd1 vccd1 _03645_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_10_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15255_ net2243 net97 net50 net2443 vssd1 vssd1 vccd1 vccd1 _00563_ sky130_fd_sc_hd__a22o_1
X_12467_ net385 _07306_ vssd1 vssd1 vccd1 vccd1 _07422_ sky130_fd_sc_hd__nor2_1
XANTENNA__12662__C _07535_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14206_ net843 ag2.body\[360\] ag2.body\[366\] net801 _08359_ vssd1 vssd1 vccd1 vccd1
+ _08367_ sky130_fd_sc_hd__o221a_1
XFILLER_0_112_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11418_ net1201 control.body\[849\] vssd1 vssd1 vccd1 vccd1 _06391_ sky130_fd_sc_hd__xor2_1
XANTENNA__12020__B1 net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15186_ net2262 net101 _01572_ net2477 vssd1 vssd1 vccd1 vccd1 _00501_ sky130_fd_sc_hd__a22o_1
X_12398_ _06636_ _07299_ _07351_ net1095 vssd1 vssd1 vccd1 vccd1 _07362_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_91_3085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11374__A2 net1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16298__C1 net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14137_ net989 ag2.body\[169\] vssd1 vssd1 vccd1 vccd1 _08298_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_91_3096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11349_ ag2.body\[441\] net1198 vssd1 vssd1 vccd1 vccd1 _06322_ sky130_fd_sc_hd__nand2_1
X_19994_ clknet_leaf_58_clk _00938_ net1471 vssd1 vssd1 vccd1 vccd1 ag2.body\[392\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_39_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18039__B1 net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14068_ net1002 ag2.body\[208\] vssd1 vssd1 vccd1 vccd1 _08229_ sky130_fd_sc_hd__xor2_1
X_18945_ clknet_leaf_139_clk img_gen.tracker.next_frame\[383\] net1290 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[383\] sky130_fd_sc_hd__dfrtp_1
X_13019_ net288 _07702_ _07703_ net1851 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[272\]
+ sky130_fd_sc_hd__a22o_1
X_18876_ clknet_leaf_12_clk img_gen.tracker.next_frame\[314\] net1282 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[314\] sky130_fd_sc_hd__dfrtp_1
X_17827_ ag2.apple_cord\[0\] net224 _03490_ net686 vssd1 vssd1 vccd1 vccd1 _01223_
+ sky130_fd_sc_hd__a211o_1
XANTENNA__14076__A1 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14076__B2 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_3560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_3571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12087__B1 net557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17758_ net350 _02211_ _03393_ _03436_ vssd1 vssd1 vccd1 vccd1 _03437_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_102_3424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_3435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_102_3446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18211__B1 net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire317_X net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16709_ obsg2.obstacleArray\[76\] net492 net483 obsg2.obstacleArray\[77\] _02387_
+ vssd1 vssd1 vccd1 vccd1 _02388_ sky130_fd_sc_hd__a221o_1
XANTENNA__11834__B1 net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18598__CLK clknet_leaf_13_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17689_ ag2.body\[152\] net888 vssd1 vssd1 vccd1 vccd1 _03368_ sky130_fd_sc_hd__xor2_1
XANTENNA__09699__B net1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15025__B1 _01555_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17565__A2 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19428_ clknet_leaf_108_clk _00372_ net1423 vssd1 vssd1 vccd1 vccd1 control.body\[962\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_3943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_3954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19359_ clknet_leaf_101_clk net2541 net1439 vssd1 vssd1 vccd1 vccd1 control.body\[1037\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_119_3965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13051__A2 _07718_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11598__C1 _06497_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_115_3818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09112_ ag2.body\[381\] vssd1 vssd1 vccd1 vccd1 _04137_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_21_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_115_3829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19993__CLK clknet_leaf_66_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09043_ ag2.body\[210\] vssd1 vssd1 vccd1 vccd1 _04068_ sky130_fd_sc_hd__inv_2
XFILLER_0_88_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15879__A2 net192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14000__A1 net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout211_A net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14000__B2 net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11102__X _06075_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_111_Right_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold410 img_gen.tracker.frame\[320\] vssd1 vssd1 vccd1 vccd1 net1972 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11469__B net1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold421 img_gen.tracker.frame\[40\] vssd1 vssd1 vccd1 vccd1 net1983 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold432 img_gen.tracker.frame\[350\] vssd1 vssd1 vccd1 vccd1 net1994 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20203_ clknet_leaf_55_clk _01147_ net1458 vssd1 vssd1 vccd1 vccd1 ag2.body\[185\]
+ sky130_fd_sc_hd__dfrtp_4
Xhold443 img_gen.tracker.frame\[154\] vssd1 vssd1 vccd1 vccd1 net2005 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_74_2571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold454 img_gen.tracker.frame\[13\] vssd1 vssd1 vccd1 vccd1 net2016 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14413__X _08574_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_2582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1120_A net1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold465 img_gen.tracker.frame\[30\] vssd1 vssd1 vccd1 vccd1 net2027 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_74_2593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold476 img_gen.tracker.frame\[498\] vssd1 vssd1 vccd1 vccd1 net2038 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1218_A net1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold487 img_gen.tracker.frame\[107\] vssd1 vssd1 vccd1 vccd1 net2049 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout901 control.body_update.curr_length\[5\] vssd1 vssd1 vccd1 vccd1 net901 sky130_fd_sc_hd__buf_2
Xhold498 img_gen.tracker.frame\[501\] vssd1 vssd1 vccd1 vccd1 net2060 sky130_fd_sc_hd__dlygate4sd3_1
X_20134_ clknet_leaf_96_clk _01078_ net1485 vssd1 vssd1 vccd1 vccd1 ag2.body\[260\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_70_2446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09945_ net758 control.body\[740\] control.body\[742\] net748 _04917_ vssd1 vssd1
+ vccd1 vccd1 _04918_ sky130_fd_sc_hd__a221o_1
Xfanout912 control.body_update.curr_length\[3\] vssd1 vssd1 vccd1 vccd1 net912 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_70_2457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout580_A net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout923 control.body_update.curr_length\[0\] vssd1 vssd1 vccd1 vccd1 net923 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_70_2468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout934 net935 vssd1 vssd1 vccd1 vccd1 net934 sky130_fd_sc_hd__buf_4
XANTENNA__20200__CLK clknet_leaf_88_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout945 obsg2.randCord\[6\] vssd1 vssd1 vccd1 vccd1 net945 sky130_fd_sc_hd__buf_4
XANTENNA_fanout678_A net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout956 net957 vssd1 vssd1 vccd1 vccd1 net956 sky130_fd_sc_hd__buf_2
X_20065_ clknet_leaf_72_clk _01009_ net1501 vssd1 vssd1 vccd1 vccd1 ag2.body\[335\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_77_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout967 net968 vssd1 vssd1 vccd1 vccd1 net967 sky130_fd_sc_hd__clkbuf_4
X_09876_ ag2.body\[163\] net1154 vssd1 vssd1 vccd1 vccd1 _04849_ sky130_fd_sc_hd__nand2_1
Xfanout978 ag2.randCord\[3\] vssd1 vssd1 vccd1 vccd1 net978 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout1006_X net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19373__CLK clknet_leaf_102_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout989 net990 vssd1 vssd1 vccd1 vccd1 net989 sky130_fd_sc_hd__buf_4
XANTENNA__16995__B net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_5_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout845_A net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout466_X net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_2965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_87_2976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_2987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_2386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_2397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11932__B net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11825__B1 net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15016__B1 _01553_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10720_ ag2.body\[618\] net774 net1047 _04226_ _05689_ vssd1 vssd1 vccd1 vccd1 _05693_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_95_578 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16764__B1 net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10548__B net1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12466__D _07312_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout800_X net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10651_ _05620_ _05621_ _05622_ _05623_ vssd1 vssd1 vccd1 vccd1 _05624_ sky130_fd_sc_hd__a22o_1
XFILLER_0_14_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_131_4310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_131_4321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10582_ ag2.body\[184\] net1233 vssd1 vssd1 vccd1 vccd1 _05555_ sky130_fd_sc_hd__xor2_1
X_13370_ net1648 _07861_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[466\]
+ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_131_4332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12321_ _07287_ vssd1 vssd1 vccd1 vccd1 _07288_ sky130_fd_sc_hd__inv_2
XFILLER_0_133_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14036__A net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11012__X _05985_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15040_ net2312 net164 _01556_ net2506 vssd1 vssd1 vccd1 vccd1 _00370_ sky130_fd_sc_hd__a22o_1
XANTENNA__09549__A2 net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12002__B1 net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12252_ _07218_ _07221_ vssd1 vssd1 vccd1 vccd1 _07222_ sky130_fd_sc_hd__or2_1
XANTENNA__10283__B net1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11203_ net1202 control.body\[873\] vssd1 vssd1 vccd1 vccd1 _06176_ sky130_fd_sc_hd__xnor2_1
XANTENNA__17347__A net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12183_ net1078 ag2.apple_cord\[6\] vssd1 vssd1 vccd1 vccd1 _07155_ sky130_fd_sc_hd__nand2_1
XANTENNA_clkbuf_leaf_61_clk_A clknet_4_13__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_4250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_4261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_1472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_129_4272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11134_ net1076 control.body\[870\] vssd1 vssd1 vccd1 vccd1 _06107_ sky130_fd_sc_hd__xnor2_1
XANTENNA__11666__Y _06638_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16991_ _04018_ net863 net711 ag2.body\[92\] vssd1 vssd1 vccd1 vccd1 _02670_ sky130_fd_sc_hd__a22o_1
XANTENNA__17066__B net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10570__Y _05543_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11065_ _06034_ _06035_ _06036_ _06037_ vssd1 vssd1 vccd1 vccd1 _06038_ sky130_fd_sc_hd__and4_1
X_15942_ ag2.body\[164\] net195 _01653_ ag2.body\[156\] vssd1 vssd1 vccd1 vccd1 _01174_
+ sky130_fd_sc_hd__a22o_1
X_18730_ clknet_leaf_141_clk img_gen.tracker.next_frame\[168\] net1261 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[168\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_34_1353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_1364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10016_ ag2.body\[268\] net1140 vssd1 vssd1 vccd1 vccd1 _04989_ sky130_fd_sc_hd__xor2_1
XANTENNA_clkbuf_leaf_76_clk_A clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18661_ clknet_leaf_13_clk img_gen.tracker.next_frame\[99\] net1282 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[99\] sky130_fd_sc_hd__dfrtp_1
X_15873_ ag2.body\[231\] net161 _01647_ ag2.body\[223\] vssd1 vssd1 vccd1 vccd1 _01113_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12778__X _07592_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18740__CLK clknet_leaf_142_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15255__B1 net50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14824_ net1040 _04047_ ag2.body\[157\] net809 _01491_ vssd1 vssd1 vccd1 vccd1 _01495_
+ sky130_fd_sc_hd__a221o_1
X_17612_ ag2.body\[604\] net959 vssd1 vssd1 vccd1 vccd1 _03291_ sky130_fd_sc_hd__xor2_1
XANTENNA__12069__B1 net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18592_ clknet_leaf_13_clk img_gen.tracker.next_frame\[30\] net1284 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[30\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_99_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13805__A1 net1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17543_ ag2.body\[325\] net954 vssd1 vssd1 vccd1 vccd1 _03222_ sky130_fd_sc_hd__xor2_1
XFILLER_0_25_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_138_4519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14322__A1_N net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14755_ net987 ag2.body\[41\] vssd1 vssd1 vccd1 vccd1 _08916_ sky130_fd_sc_hd__xor2_1
XANTENNA__10298__X _05271_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09485__A1 _04447_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11967_ img_gen.tracker.frame\[514\] net583 vssd1 vssd1 vccd1 vccd1 _06939_ sky130_fd_sc_hd__or2_1
XANTENNA__15007__B1 _01552_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13281__A2 _07825_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13706_ track.highScore\[5\] _08028_ _08031_ track.highScore\[6\] vssd1 vssd1 vccd1
+ vccd1 _08047_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_47_1758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17474_ ag2.body\[133\] net953 vssd1 vssd1 vccd1 vccd1 _03153_ sky130_fd_sc_hd__or2_1
X_10918_ ag2.body\[460\] net1127 vssd1 vssd1 vccd1 vccd1 _05891_ sky130_fd_sc_hd__nand2_1
XANTENNA__16755__B1 net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14686_ net837 ag2.body\[89\] _04022_ net1011 _08846_ vssd1 vssd1 vccd1 vccd1 _08847_
+ sky130_fd_sc_hd__o221a_1
XANTENNA__19164__RESET_B net1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_1769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10458__B net1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11898_ img_gen.tracker.frame\[70\] net579 net568 _06869_ vssd1 vssd1 vccd1 vccd1
+ _06870_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_131_1454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_28_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16425_ _02057_ _02103_ _02102_ _02086_ vssd1 vssd1 vccd1 vccd1 _02104_ sky130_fd_sc_hd__o211ai_1
X_19213_ clknet_leaf_85_clk _00157_ net1463 vssd1 vssd1 vccd1 vccd1 ag2.body\[76\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA_clkbuf_leaf_134_clk_A clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13637_ control.divider.count\[13\] _07997_ net222 vssd1 vssd1 vccd1 vccd1 _07999_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_131_1487 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10849_ ag2.body\[45\] net1097 vssd1 vssd1 vccd1 vccd1 _05822_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_15_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19144_ clknet_leaf_51_clk _00088_ net1377 vssd1 vssd1 vccd1 vccd1 ag2.body\[8\]
+ sky130_fd_sc_hd__dfrtp_4
X_16356_ obsg2.obstacleArray\[0\] obsg2.obstacleArray\[1\] net409 vssd1 vssd1 vccd1
+ vccd1 _02035_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_14_clk_A clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_97_3272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13568_ ssdec1.in\[3\] _07943_ _07946_ vssd1 vssd1 vccd1 vccd1 net20 sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_97_3283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16145__B net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_97_3294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15794__A_N _04983_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11595__A2 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15307_ net2570 net75 _01586_ net2308 vssd1 vssd1 vccd1 vccd1 _00608_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_93_3147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19075_ clknet_leaf_29_clk img_gen.tracker.next_frame\[513\] net1334 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[513\] sky130_fd_sc_hd__dfrtp_1
X_12519_ net226 _07455_ _07456_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[20\]
+ sky130_fd_sc_hd__o21bai_1
X_16287_ _01964_ _01965_ net419 vssd1 vssd1 vccd1 vccd1 _01966_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_3158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13499_ net276 _07910_ _07911_ net2012 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[545\]
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_93_3169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18026_ net351 net38 _03633_ vssd1 vssd1 vccd1 vccd1 _03634_ sky130_fd_sc_hd__and3_1
X_15238_ control.body\[785\] net96 _01578_ net2439 vssd1 vssd1 vccd1 vccd1 _00547_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__10193__B net1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_29_clk_A clknet_4_4__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15169_ control.body\[852\] net102 _01570_ net2449 vssd1 vssd1 vccd1 vccd1 _00486_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_103_1501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19396__CLK clknet_leaf_103_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout208 net209 vssd1 vssd1 vccd1 vccd1 net208 sky130_fd_sc_hd__buf_2
Xfanout219 _08130_ vssd1 vssd1 vccd1 vccd1 net219 sky130_fd_sc_hd__buf_4
XANTENNA__09960__A2 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16901__A2_N net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19977_ clknet_leaf_62_clk _00921_ net1470 vssd1 vssd1 vccd1 vccd1 ag2.body\[423\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_10_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_108_3611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09730_ ag2.body\[94\] net1089 vssd1 vssd1 vccd1 vccd1 _04703_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_108_3622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18928_ clknet_leaf_140_clk img_gen.tracker.next_frame\[366\] net1290 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[366\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_66_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_105_Left_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_104_3508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09661_ net919 net638 _04632_ vssd1 vssd1 vccd1 vccd1 _04634_ sky130_fd_sc_hd__or3_1
XANTENNA__14049__A1 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18859_ clknet_leaf_18_clk img_gen.tracker.next_frame\[297\] net1323 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[297\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__14049__B2 net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16100__S net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15797__A1 ag2.body\[290\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09592_ net1084 control.body\[910\] vssd1 vssd1 vccd1 vccd1 _04565_ sky130_fd_sc_hd__xor2_1
XFILLER_0_82_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout161_A net162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17538__A2 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout259_A net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_2250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16210__A2 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__20492__RESET_B net1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_114_Left_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10936__X _05909_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_1549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout426_A net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1168_A net1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12783__A1 net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout214_X net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_76_2633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_76_2644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09026_ ag2.body\[166\] vssd1 vssd1 vccd1 vccd1 _04051_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_76_2655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_1445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_72_2508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_57_2054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_2065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout795_A net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_1433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_57_2076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09892__B net1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold240 img_gen.tracker.frame\[444\] vssd1 vssd1 vccd1 vccd1 net1802 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1502_A net1504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold251 img_gen.tracker.frame\[227\] vssd1 vssd1 vccd1 vccd1 net1813 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1123_X net1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold262 img_gen.tracker.frame\[93\] vssd1 vssd1 vccd1 vccd1 net1824 sky130_fd_sc_hd__dlygate4sd3_1
Xhold273 img_gen.tracker.frame\[174\] vssd1 vssd1 vccd1 vccd1 net1835 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11486__Y _06459_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold284 img_gen.tracker.frame\[439\] vssd1 vssd1 vccd1 vccd1 net1846 sky130_fd_sc_hd__dlygate4sd3_1
Xhold295 img_gen.tracker.frame\[389\] vssd1 vssd1 vccd1 vccd1 net1857 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_123_Left_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10831__B net1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout962_A net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout583_X net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout720 net721 vssd1 vssd1 vccd1 vccd1 net720 sky130_fd_sc_hd__buf_4
XANTENNA__18763__CLK clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15485__B1 _01605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19889__CLK clknet_leaf_83_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout731 _04263_ vssd1 vssd1 vccd1 vccd1 net731 sky130_fd_sc_hd__clkbuf_4
X_20117_ clknet_leaf_80_clk _01061_ net1488 vssd1 vssd1 vccd1 vccd1 ag2.body\[275\]
+ sky130_fd_sc_hd__dfrtp_4
Xfanout742 _04235_ vssd1 vssd1 vccd1 vccd1 net742 sky130_fd_sc_hd__buf_4
X_09928_ _04818_ _04846_ _04876_ _04900_ vssd1 vssd1 vccd1 vccd1 _04901_ sky130_fd_sc_hd__and4_1
Xfanout753 net754 vssd1 vssd1 vccd1 vccd1 net753 sky130_fd_sc_hd__buf_4
Xfanout764 net765 vssd1 vssd1 vccd1 vccd1 net764 sky130_fd_sc_hd__buf_2
XFILLER_0_102_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout775 _04229_ vssd1 vssd1 vccd1 vccd1 net775 sky130_fd_sc_hd__buf_4
X_20048_ clknet_leaf_68_clk _00992_ net1498 vssd1 vssd1 vccd1 vccd1 ag2.body\[350\]
+ sky130_fd_sc_hd__dfrtp_4
Xfanout786 net787 vssd1 vssd1 vccd1 vccd1 net786 sky130_fd_sc_hd__clkbuf_4
Xfanout797 _03973_ vssd1 vssd1 vccd1 vccd1 net797 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout750_X net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09859_ net903 _04238_ _04420_ _04470_ _04831_ vssd1 vssd1 vccd1 vccd1 _04832_ sky130_fd_sc_hd__o41a_2
XFILLER_0_99_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1492_X net1492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15237__B1 _01578_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout848_X net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19119__CLK clknet_leaf_141_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14957__C net65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12870_ _06673_ _07305_ _07444_ vssd1 vssd1 vccd1 vccd1 _07636_ sky130_fd_sc_hd__and3_1
XFILLER_0_99_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15788__B2 ag2.body\[290\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16985__B1 net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11821_ net560 _06792_ _06790_ vssd1 vssd1 vccd1 vccd1 _06793_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_115_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_1464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14540_ net1001 ag2.body\[240\] vssd1 vssd1 vccd1 vccd1 _08701_ sky130_fd_sc_hd__or2_1
XFILLER_0_96_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_1546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11752_ net466 _06673_ _06722_ vssd1 vssd1 vccd1 vccd1 _06724_ sky130_fd_sc_hd__a21o_2
XANTENNA__16737__B1 net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_132_Left_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10703_ _05672_ _05673_ _05674_ _05675_ vssd1 vssd1 vccd1 vccd1 _05676_ sky130_fd_sc_hd__a22o_1
X_14471_ net975 _04091_ _04092_ net1010 _08627_ vssd1 vssd1 vccd1 vccd1 _08632_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_42_1600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14318__X _08479_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11683_ img_gen.tracker.frame\[122\] net619 net601 img_gen.tracker.frame\[125\] vssd1
+ vssd1 vccd1 vccd1 _06655_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_12_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16210_ net956 net703 net696 net690 _01888_ vssd1 vssd1 vccd1 vccd1 _01889_ sky130_fd_sc_hd__a41o_1
XTAP_TAPCELL_ROW_23_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_740 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13422_ net236 _07880_ _07881_ net2038 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[498\]
+ sky130_fd_sc_hd__a22o_1
X_10634_ net1070 control.body\[670\] vssd1 vssd1 vccd1 vccd1 _05607_ sky130_fd_sc_hd__or2_1
XFILLER_0_52_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17190_ ag2.body\[572\] net710 net705 ag2.body\[573\] _02865_ vssd1 vssd1 vccd1 vccd1
+ _02869_ sky130_fd_sc_hd__a221o_1
XFILLER_0_11_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_1322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16141_ obsg2.obstacleArray\[0\] obsg2.obstacleArray\[1\] net427 vssd1 vssd1 vccd1
+ vccd1 _01820_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13353_ net670 _07854_ vssd1 vssd1 vccd1 vccd1 _07855_ sky130_fd_sc_hd__nor2_1
X_10565_ net1132 ag2.body\[516\] vssd1 vssd1 vccd1 vccd1 _05538_ sky130_fd_sc_hd__and2b_1
XFILLER_0_107_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12304_ _07228_ _07267_ _07269_ _07265_ _07266_ vssd1 vssd1 vccd1 vccd1 _07271_ sky130_fd_sc_hd__a311o_1
X_16072_ net348 _01750_ _01747_ _01743_ vssd1 vssd1 vccd1 vccd1 _01751_ sky130_fd_sc_hd__o211a_1
XFILLER_0_106_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13284_ net670 _07827_ vssd1 vssd1 vccd1 vccd1 _07828_ sky130_fd_sc_hd__nor2_1
X_10496_ ag2.body\[544\] net1228 vssd1 vssd1 vccd1 vccd1 _05469_ sky130_fd_sc_hd__xnor2_1
X_19900_ clknet_leaf_57_clk _00844_ net1464 vssd1 vssd1 vccd1 vccd1 ag2.body\[490\]
+ sky130_fd_sc_hd__dfrtp_4
X_15023_ control.body\[977\] net167 _01555_ control.body\[969\] vssd1 vssd1 vccd1
+ vccd1 _00355_ sky130_fd_sc_hd__a22o_1
XFILLER_0_60_990 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11677__X _06649_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12235_ _04274_ _07196_ vssd1 vssd1 vccd1 vccd1 _07205_ sky130_fd_sc_hd__and2_1
XFILLER_0_47_1090 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_127_4209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_36_1415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_1566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19831_ clknet_leaf_124_clk _00775_ net1408 vssd1 vssd1 vccd1 vccd1 ag2.body\[565\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_102_591 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09942__A2 net1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15309__B net53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12166_ img_gen.tracker.frame\[411\] net600 net584 img_gen.tracker.frame\[417\] vssd1
+ vssd1 vccd1 vccd1 _07138_ sky130_fd_sc_hd__o22a_1
XANTENNA__10741__B net1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11117_ net1232 _04256_ _04861_ _06089_ control.body_update.curr_length\[7\] vssd1
+ vssd1 vccd1 vccd1 _06090_ sky130_fd_sc_hd__o2111a_4
X_19762_ clknet_leaf_127_clk _00706_ net1326 vssd1 vssd1 vccd1 vccd1 control.body\[624\]
+ sky130_fd_sc_hd__dfrtp_1
X_16974_ ag2.body\[427\] net851 vssd1 vssd1 vccd1 vccd1 _02653_ sky130_fd_sc_hd__xnor2_1
X_12097_ img_gen.tracker.frame\[336\] net627 net593 img_gen.tracker.frame\[345\] vssd1
+ vssd1 vccd1 vccd1 _07069_ sky130_fd_sc_hd__a22o_1
XFILLER_0_120_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18713_ clknet_leaf_144_clk img_gen.tracker.next_frame\[151\] net1252 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[151\] sky130_fd_sc_hd__dfrtp_1
X_11048_ ag2.body\[391\] net1056 vssd1 vssd1 vccd1 vccd1 _06021_ sky130_fd_sc_hd__xor2_1
X_15925_ ag2.body\[180\] net124 _01654_ ag2.body\[172\] vssd1 vssd1 vccd1 vccd1 _01158_
+ sky130_fd_sc_hd__a22o_1
X_19693_ clknet_leaf_136_clk _00637_ net1300 vssd1 vssd1 vccd1 vccd1 control.body\[699\]
+ sky130_fd_sc_hd__dfrtp_1
Xinput8 gpio_in[31] vssd1 vssd1 vccd1 vccd1 net8 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_56_1304 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18644_ clknet_leaf_15_clk img_gen.tracker.next_frame\[82\] net1312 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[82\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_49_1809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15856_ _04740_ net59 vssd1 vssd1 vccd1 vccd1 _01646_ sky130_fd_sc_hd__nor2_2
XFILLER_0_56_1359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14807_ _01472_ _01477_ vssd1 vssd1 vccd1 vccd1 _01478_ sky130_fd_sc_hd__nand2b_1
X_15787_ ag2.body\[297\] net209 _01639_ ag2.body\[289\] vssd1 vssd1 vccd1 vccd1 _01035_
+ sky130_fd_sc_hd__a22o_1
X_18575_ clknet_leaf_14_clk img_gen.tracker.next_frame\[13\] net1279 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[13\] sky130_fd_sc_hd__dfrtp_1
X_12999_ net229 _07694_ _07695_ net2039 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[261\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_98_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11265__A1 _05543_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14738_ net839 ag2.body\[329\] ag2.body\[330\] net830 _08898_ vssd1 vssd1 vccd1 vccd1
+ _08899_ sky130_fd_sc_hd__a221o_1
X_17526_ _04175_ net852 net710 ag2.body\[484\] _03204_ vssd1 vssd1 vccd1 vccd1 _03205_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_15_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16728__B1 net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_3334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_99_3345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17457_ ag2.body\[432\] net737 net930 _04155_ vssd1 vssd1 vccd1 vccd1 _03136_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_99_3356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14669_ _08823_ _08824_ _08828_ _08829_ vssd1 vssd1 vccd1 vccd1 _08830_ sky130_fd_sc_hd__or4b_1
XTAP_TAPCELL_ROW_95_3209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15400__B1 _01581_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16408_ obsg2.obstacleArray\[98\] net452 vssd1 vssd1 vccd1 vccd1 _02087_ sky130_fd_sc_hd__or2_1
XFILLER_0_129_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18636__CLK clknet_leaf_131_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17388_ ag2.body\[489\] net734 net693 ag2.body\[495\] vssd1 vssd1 vccd1 vccd1 _03067_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__10916__B net1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12765__A1 net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16339_ obsg2.obstacleArray\[82\] obsg2.obstacleArray\[83\] net411 vssd1 vssd1 vccd1
+ vccd1 _02018_ sky130_fd_sc_hd__mux2_1
X_19127_ clknet_leaf_140_clk img_gen.tracker.next_frame\[565\] net1296 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[565\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__17539__X _03218_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16590__S net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17153__B1 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19058_ clknet_leaf_9_clk img_gen.tracker.next_frame\[496\] net1271 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[496\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__16900__B1 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18786__CLK clknet_leaf_13_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18009_ net432 net463 net495 net491 vssd1 vssd1 vccd1 vccd1 _03621_ sky130_fd_sc_hd__and4_1
XANTENNA__14404__A net1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_1099 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15467__B1 _01603_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09713_ net912 _04427_ net642 vssd1 vssd1 vccd1 vccd1 _04686_ sky130_fd_sc_hd__a21oi_4
XANTENNA__17434__B net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12859__A _07431_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout376_A net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09644_ net775 control.body\[1018\] control.body\[1023\] net746 _04616_ vssd1 vssd1
+ vccd1 vccd1 _04617_ sky130_fd_sc_hd__a221o_1
XFILLER_0_74_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_65_2301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_2312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09575_ ag2.body\[203\] net1162 vssd1 vssd1 vccd1 vccd1 _04548_ sky130_fd_sc_hd__xor2_1
XANTENNA__19411__CLK clknet_leaf_105_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout543_A net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10059__A2 net1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16719__B1 net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09520__X _04493_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16195__A1 net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout331_X net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout710_A net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout429_X net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout808_A net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1073_X net1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1452_A net1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15942__A1 ag2.body\[164\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_367 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_2706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19561__CLK clknet_leaf_115_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_2717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10826__B net1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_2116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_2127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_592 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20597_ net1529 vssd1 vssd1 vccd1 vccd1 gpio_oeb[9] sky130_fd_sc_hd__buf_2
XANTENNA__17144__B1 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1338_X net1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_765 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10350_ _05320_ _05321_ _05322_ _04418_ vssd1 vssd1 vccd1 vccd1 _05323_ sky130_fd_sc_hd__a211o_1
XANTENNA__17609__B net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_798 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout798_X net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09009_ ag2.body\[130\] vssd1 vssd1 vccd1 vccd1 _04034_ sky130_fd_sc_hd__inv_2
XFILLER_0_130_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10281_ net905 net918 net914 net910 vssd1 vssd1 vccd1 vccd1 _05254_ sky130_fd_sc_hd__or4b_4
XANTENNA__10519__B1 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1505_X net1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_3_0_clk_X clknet_3_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11716__C1 _06660_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12020_ img_gen.tracker.frame\[216\] net630 net577 _06991_ vssd1 vssd1 vccd1 vccd1
+ _06992_ sky130_fd_sc_hd__a211o_1
XANTENNA__11657__B net1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout965_X net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10561__B net1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1504 net1505 vssd1 vssd1 vccd1 vccd1 net1504 sky130_fd_sc_hd__buf_2
XANTENNA__15458__B1 _01602_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1515 net1517 vssd1 vssd1 vccd1 vccd1 net1515 sky130_fd_sc_hd__clkbuf_2
Xfanout550 net553 vssd1 vssd1 vccd1 vccd1 net550 sky130_fd_sc_hd__buf_2
Xfanout561 net562 vssd1 vssd1 vccd1 vccd1 net561 sky130_fd_sc_hd__buf_2
Xfanout572 net573 vssd1 vssd1 vccd1 vccd1 net572 sky130_fd_sc_hd__clkbuf_2
X_13971_ ag2.body\[110\] net202 _08157_ ag2.body\[102\] vssd1 vssd1 vccd1 vccd1 _00191_
+ sky130_fd_sc_hd__a22o_1
Xfanout583 net586 vssd1 vssd1 vccd1 vccd1 net583 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09688__A1 _04647_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12769__A net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout594 net595 vssd1 vssd1 vccd1 vccd1 net594 sky130_fd_sc_hd__buf_4
XANTENNA__09688__B2 _04606_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15710_ ag2.body\[374\] net140 _01629_ ag2.body\[366\] vssd1 vssd1 vccd1 vccd1 _00968_
+ sky130_fd_sc_hd__a22o_1
X_12922_ net290 _07656_ _07657_ net1792 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[221\]
+ sky130_fd_sc_hd__a22o_1
X_16690_ _02278_ _02365_ _02367_ _02368_ _02243_ vssd1 vssd1 vccd1 vccd1 _02369_ sky130_fd_sc_hd__o221a_1
X_15641_ _06066_ net64 vssd1 vssd1 vccd1 vccd1 _01623_ sky130_fd_sc_hd__and2_2
XFILLER_0_57_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19091__CLK clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12853_ _07431_ _07627_ vssd1 vssd1 vccd1 vccd1 _07628_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_17_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15630__B1 _01621_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11804_ img_gen.tracker.frame\[434\] net613 net582 img_gen.tracker.frame\[443\] vssd1
+ vssd1 vccd1 vccd1 _06776_ sky130_fd_sc_hd__o22a_1
X_18360_ _03830_ _03834_ _03824_ vssd1 vssd1 vccd1 vccd1 _03855_ sky130_fd_sc_hd__o21a_1
X_15572_ ag2.body\[490\] net135 _01615_ ag2.body\[482\] vssd1 vssd1 vccd1 vccd1 _00844_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_90_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__20343__RESET_B net1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1488 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18659__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12784_ net336 net332 _07493_ vssd1 vssd1 vccd1 vccd1 _07595_ sky130_fd_sc_hd__or3_1
XFILLER_0_29_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17311_ ag2.body\[392\] net738 net733 ag2.body\[393\] _02989_ vssd1 vssd1 vccd1 vccd1
+ _02990_ sky130_fd_sc_hd__a221o_1
XFILLER_0_95_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12995__A1 net254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14523_ net1038 ag2.body\[252\] vssd1 vssd1 vccd1 vccd1 _08684_ sky130_fd_sc_hd__or2_1
XFILLER_0_113_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18291_ net326 net325 vssd1 vssd1 vccd1 vccd1 _03787_ sky130_fd_sc_hd__or2_2
X_11735_ img_gen.tracker.frame\[35\] net585 net546 img_gen.tracker.frame\[32\] _06706_
+ vssd1 vssd1 vccd1 vccd1 _06707_ sky130_fd_sc_hd__o221a_1
XFILLER_0_138_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17242_ _04222_ net879 net710 ag2.body\[620\] _02920_ vssd1 vssd1 vccd1 vccd1 _02921_
+ sky130_fd_sc_hd__o221a_1
X_14454_ net812 ag2.body\[436\] ag2.body\[438\] net800 _08614_ vssd1 vssd1 vccd1 vccd1
+ _08615_ sky130_fd_sc_hd__a221o_1
X_11666_ net767 _06636_ vssd1 vssd1 vccd1 vccd1 _06638_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_37_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15933__B2 ag2.body\[163\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12747__A1 net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13405_ net313 _07555_ vssd1 vssd1 vccd1 vccd1 _07874_ sky130_fd_sc_hd__and2_1
X_17173_ ag2.body\[457\] net870 vssd1 vssd1 vccd1 vccd1 _02852_ sky130_fd_sc_hd__or2_1
X_10617_ ag2.body\[50\] net774 net753 ag2.body\[53\] _05589_ vssd1 vssd1 vccd1 vccd1
+ _05590_ sky130_fd_sc_hd__a221o_1
XANTENNA__12654__D net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14385_ net844 ag2.body\[296\] _04099_ net1039 _08545_ vssd1 vssd1 vccd1 vccd1 _08546_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_3_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11597_ net507 _06566_ _06569_ net475 vssd1 vssd1 vccd1 vccd1 _06570_ sky130_fd_sc_hd__o211a_1
X_16124_ obsg2.obstacleArray\[89\] net431 vssd1 vssd1 vccd1 vccd1 _01803_ sky130_fd_sc_hd__or2_1
X_13336_ net274 _07846_ _07847_ net1911 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[446\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_49_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10548_ ag2.body\[225\] net1206 vssd1 vssd1 vccd1 vccd1 _05521_ sky130_fd_sc_hd__or2_1
Xclkbuf_4_5__f_clk clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_5__leaf_clk sky130_fd_sc_hd__clkbuf_16
XANTENNA__17519__B net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16055_ _01715_ _01725_ _01733_ vssd1 vssd1 vccd1 vccd1 _01734_ sky130_fd_sc_hd__o21a_1
X_13267_ net280 _07819_ _07820_ net1788 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[404\]
+ sky130_fd_sc_hd__a22o_1
X_10479_ net637 _05450_ vssd1 vssd1 vccd1 vccd1 _05452_ sky130_fd_sc_hd__nand2_1
XFILLER_0_110_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13172__A1 net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15006_ net2584 net152 _01552_ control.body\[987\] vssd1 vssd1 vccd1 vccd1 _00341_
+ sky130_fd_sc_hd__a22o_1
X_12218_ img_gen.updater.commands.mode\[1\] _04391_ vssd1 vssd1 vccd1 vccd1 _07188_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_23_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_88_3002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13198_ net240 _07788_ _07789_ net1884 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[366\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_104_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15449__B1 _01601_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16646__C1 net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_3013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19814_ clknet_leaf_125_clk _00758_ net1410 vssd1 vssd1 vccd1 vccd1 ag2.body\[580\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__16110__A1 net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12149_ img_gen.tracker.frame\[447\] net597 net578 img_gen.tracker.frame\[453\] vssd1
+ vssd1 vccd1 vccd1 _07121_ sky130_fd_sc_hd__o22a_1
XFILLER_0_47_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19745_ clknet_leaf_131_clk _00689_ net1304 vssd1 vssd1 vccd1 vccd1 control.body\[655\]
+ sky130_fd_sc_hd__dfrtp_1
X_16957_ ag2.body\[294\] net700 net692 ag2.body\[295\] vssd1 vssd1 vccd1 vccd1 _02636_
+ sky130_fd_sc_hd__o22a_1
XANTENNA__18399__C1 net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14672__B2 net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11583__A net1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15908_ ag2.body\[198\] net129 _01651_ ag2.body\[190\] vssd1 vssd1 vccd1 vccd1 _01144_
+ sky130_fd_sc_hd__a22o_1
X_19676_ clknet_leaf_117_clk _00620_ net1384 vssd1 vssd1 vccd1 vccd1 control.body\[714\]
+ sky130_fd_sc_hd__dfrtp_1
X_16888_ ag2.body\[208\] net739 net727 ag2.body\[210\] vssd1 vssd1 vccd1 vccd1 _02567_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__17610__A1 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1025 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16413__A2 _02059_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18627_ clknet_leaf_0_clk img_gen.tracker.next_frame\[65\] net1243 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[65\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_133_1313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1167 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15839_ ag2.body\[248\] net181 _01644_ ag2.body\[240\] vssd1 vssd1 vccd1 vccd1 _01082_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_137_1493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09360_ _04361_ vssd1 vssd1 vccd1 vccd1 _04362_ sky130_fd_sc_hd__inv_2
X_18558_ clknet_leaf_132_clk _00084_ net1303 vssd1 vssd1 vccd1 vccd1 ag2.x\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_34_1432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18166__A2 _03539_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17509_ ag2.body\[588\] net961 vssd1 vssd1 vccd1 vccd1 _03188_ sky130_fd_sc_hd__xor2_1
X_09291_ sound_gen.osc1.count\[4\] sound_gen.osc1.count\[3\] _04310_ _04309_ sound_gen.osc1.count\[6\]
+ vssd1 vssd1 vccd1 vccd1 _04311_ sky130_fd_sc_hd__a32o_1
X_18489_ net1516 net1510 vssd1 vssd1 vccd1 vccd1 _00020_ sky130_fd_sc_hd__or2_1
XANTENNA__09851__A1 net1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10997__B1 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09851__B2 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12450__A3 net1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_13 _03446_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13303__A net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09500__B net1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20520_ clknet_leaf_93_clk track.nextCurrScore\[2\] net1413 vssd1 vssd1 vccd1 vccd1
+ control.body_update.curr_length\[2\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_24 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_35 _06837_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkload63_A clknet_leaf_52_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20451_ clknet_leaf_41_clk _01338_ net1371 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[87\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_133_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18469__A3 net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout124_A net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20382_ clknet_leaf_40_clk _01269_ net1374 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[18\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_70_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14134__A net1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10662__A net1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1033_A ag2.randCord\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11477__B net1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout493_A _01736_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10381__B net1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16637__C1 net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13973__A _05162_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11713__A2 net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1200_A ag2.y\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19267__RESET_B net1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13692__B _04427_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17164__B net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout281_X net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout758_A net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout379_X net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17732__X _03411_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19927__CLK clknet_leaf_51_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09627_ net897 _04237_ net921 vssd1 vssd1 vccd1 vccd1 _04600_ sky130_fd_sc_hd__and3_2
XANTENNA_fanout1190_X net1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout925_A net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15612__B1 _01620_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_459 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14415__B2 net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout546_X net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09558_ net1148 control.body\[723\] vssd1 vssd1 vccd1 vccd1 _04531_ sky130_fd_sc_hd__xor2_1
XFILLER_0_91_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout37_A _03705_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout713_X net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09489_ ag2.body\[371\] net1154 vssd1 vssd1 vccd1 vccd1 _04462_ sky130_fd_sc_hd__xor2_1
XANTENNA__18951__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_403 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14309__A net1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1455_X net1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13213__A net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11520_ _06491_ _06492_ vssd1 vssd1 vccd1 vccd1 _06493_ sky130_fd_sc_hd__or2_1
XFILLER_0_92_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_1216 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12729__A1 net237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11451_ net1110 control.body\[957\] vssd1 vssd1 vccd1 vccd1 _06424_ sky130_fd_sc_hd__xor2_1
XANTENNA__17117__B1 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11937__C1 net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10402_ _04632_ _04758_ vssd1 vssd1 vccd1 vccd1 _05375_ sky130_fd_sc_hd__nor2_1
XFILLER_0_61_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10204__A2 _05170_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14170_ net997 _04062_ ag2.body\[201\] net836 vssd1 vssd1 vccd1 vccd1 _08331_ sky130_fd_sc_hd__a22o_1
X_11382_ net1220 control.body\[640\] vssd1 vssd1 vccd1 vccd1 _06355_ sky130_fd_sc_hd__or2_1
X_20589__1521 vssd1 vssd1 vccd1 vccd1 _20589__1521/HI net1521 sky130_fd_sc_hd__conb_1
XANTENNA__15679__B1 _01627_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1216 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11072__A2_N net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11952__A2 net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11668__A net1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13121_ net343 _07584_ vssd1 vssd1 vccd1 vccd1 _07752_ sky130_fd_sc_hd__nor2_1
XANTENNA__17907__X _03542_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10333_ ag2.body\[523\] net1159 vssd1 vssd1 vccd1 vccd1 _05306_ sky130_fd_sc_hd__nand2_1
XFILLER_0_127_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14044__A net997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13052_ net293 _07718_ _07719_ net1870 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[290\]
+ sky130_fd_sc_hd__a22o_1
X_10264_ net908 _04471_ _04419_ vssd1 vssd1 vccd1 vccd1 _05237_ sky130_fd_sc_hd__a21oi_4
XANTENNA__10291__B net1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16628__C1 net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12003_ img_gen.tracker.frame\[442\] net578 net540 img_gen.tracker.frame\[439\] _06974_
+ vssd1 vssd1 vccd1 vccd1 _06975_ sky130_fd_sc_hd__o221a_1
XANTENNA__12901__A1 net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18093__A1 net38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13883__A _05670_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1301 net1302 vssd1 vssd1 vccd1 vccd1 net1301 sky130_fd_sc_hd__clkbuf_4
X_10195_ ag2.body\[116\] net1141 vssd1 vssd1 vccd1 vccd1 _05168_ sky130_fd_sc_hd__xor2_1
X_17860_ net2177 _03499_ vssd1 vssd1 vccd1 vccd1 _01235_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_20_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1312 net1314 vssd1 vssd1 vccd1 vccd1 net1312 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_24_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1323 net1324 vssd1 vssd1 vccd1 vccd1 net1323 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08977__A ag2.body\[71\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1334 net1338 vssd1 vssd1 vccd1 vccd1 net1334 sky130_fd_sc_hd__clkbuf_4
X_16811_ ag2.body\[66\] net728 net720 ag2.body\[67\] _02482_ vssd1 vssd1 vccd1 vccd1
+ _02490_ sky130_fd_sc_hd__a221o_1
Xfanout1345 net1357 vssd1 vssd1 vccd1 vccd1 net1345 sky130_fd_sc_hd__buf_2
Xfanout1356 net1357 vssd1 vssd1 vccd1 vccd1 net1356 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_108_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17074__B net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17791_ net1017 _03463_ _03464_ net1036 vssd1 vssd1 vccd1 vccd1 _03467_ sky130_fd_sc_hd__o22ai_1
Xfanout1367 net1369 vssd1 vssd1 vccd1 vccd1 net1367 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12499__A net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14654__A1 net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1378 net1380 vssd1 vssd1 vccd1 vccd1 net1378 sky130_fd_sc_hd__clkbuf_4
Xclkbuf_4_13__f_clk clknet_3_6_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_13__leaf_clk
+ sky130_fd_sc_hd__clkbuf_16
Xfanout380 net381 vssd1 vssd1 vccd1 vccd1 net380 sky130_fd_sc_hd__buf_2
XANTENNA__14654__B2 net1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout391 net393 vssd1 vssd1 vccd1 vccd1 net391 sky130_fd_sc_hd__buf_2
Xfanout1389 net1404 vssd1 vssd1 vccd1 vccd1 net1389 sky130_fd_sc_hd__clkbuf_4
X_19530_ clknet_leaf_120_clk _00474_ net1393 vssd1 vssd1 vccd1 vccd1 control.body\[856\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11468__A1 net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13954_ ag2.body\[95\] net190 _08155_ ag2.body\[87\] vssd1 vssd1 vccd1 vccd1 _00176_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_92_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16742_ obsg2.obstacleArray\[35\] net500 net486 obsg2.obstacleArray\[34\] vssd1 vssd1
+ vccd1 vccd1 _02421_ sky130_fd_sc_hd__a22o_1
XANTENNA__11563__S1 net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12905_ img_gen.tracker.frame\[211\] net661 vssd1 vssd1 vccd1 vccd1 _07652_ sky130_fd_sc_hd__and2_1
X_16673_ _02350_ _02351_ net392 vssd1 vssd1 vccd1 vccd1 _02352_ sky130_fd_sc_hd__mux2_1
X_19461_ clknet_leaf_112_clk _00405_ net1425 vssd1 vssd1 vccd1 vccd1 control.body\[931\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14406__A1 net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13885_ ag2.body\[33\] net118 _08148_ ag2.body\[25\] vssd1 vssd1 vccd1 vccd1 _00114_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_18_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14406__B2 net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15603__B1 _01619_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1190 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17090__A ag2.body\[303\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18412_ _04639_ _03823_ _03841_ vssd1 vssd1 vccd1 vccd1 _03902_ sky130_fd_sc_hd__a21oi_1
X_15624_ ag2.body\[440\] net125 _01621_ ag2.body\[432\] vssd1 vssd1 vccd1 vccd1 _00890_
+ sky130_fd_sc_hd__a22o_1
X_12836_ net676 _07619_ vssd1 vssd1 vccd1 vccd1 _07620_ sky130_fd_sc_hd__nor2_1
X_19392_ clknet_leaf_102_clk _00336_ net1428 vssd1 vssd1 vccd1 vccd1 control.body\[1006\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_1632 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18148__A2 _03574_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12946__B net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12968__A1 net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15555_ ag2.body\[508\] net186 _01612_ ag2.body\[500\] vssd1 vssd1 vccd1 vccd1 _00830_
+ sky130_fd_sc_hd__a22o_1
X_18343_ _04236_ _08028_ _08031_ _03838_ _08035_ vssd1 vssd1 vccd1 vccd1 _03839_ sky130_fd_sc_hd__o221a_1
XFILLER_0_70_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12767_ net333 _07483_ vssd1 vssd1 vccd1 vccd1 _07587_ sky130_fd_sc_hd__or2_2
XFILLER_0_29_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14506_ net973 ag2.body\[179\] vssd1 vssd1 vccd1 vccd1 _08667_ sky130_fd_sc_hd__xor2_1
XFILLER_0_31_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18274_ net319 _03571_ obsg2.obstacleArray\[134\] vssd1 vssd1 vccd1 vccd1 _03776_
+ sky130_fd_sc_hd__a21oi_1
X_11718_ net466 _06673_ vssd1 vssd1 vccd1 vccd1 _06690_ sky130_fd_sc_hd__nor2_1
XFILLER_0_86_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15486_ ag2.body\[574\] net112 _01605_ ag2.body\[566\] vssd1 vssd1 vccd1 vccd1 _00768_
+ sky130_fd_sc_hd__a22o_1
X_12698_ net310 _07553_ net673 vssd1 vssd1 vccd1 vccd1 _07554_ sky130_fd_sc_hd__a21oi_1
X_17225_ _04107_ net944 net694 ag2.body\[319\] _02903_ vssd1 vssd1 vccd1 vccd1 _02904_
+ sky130_fd_sc_hd__o221a_1
X_14437_ net1006 ag2.body\[23\] vssd1 vssd1 vccd1 vccd1 _08598_ sky130_fd_sc_hd__xor2_1
XANTENNA__17089__X _02768_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17108__B1 net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11649_ _06511_ _06528_ vssd1 vssd1 vccd1 vccd1 _06622_ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_626 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09597__B1 _04569_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17156_ _02828_ _02829_ _02834_ _02827_ vssd1 vssd1 vccd1 vccd1 _02835_ sky130_fd_sc_hd__a211o_1
XFILLER_0_64_1403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14368_ net817 ag2.body\[603\] ag2.body\[607\] net790 _08522_ vssd1 vssd1 vccd1 vccd1
+ _08529_ sky130_fd_sc_hd__o221a_1
XANTENNA__16153__B net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold806 control.body\[1009\] vssd1 vssd1 vccd1 vccd1 net2368 sky130_fd_sc_hd__dlygate4sd3_1
X_16107_ obsg2.obstacleArray\[84\] obsg2.obstacleArray\[85\] net428 vssd1 vssd1 vccd1
+ vccd1 _01786_ sky130_fd_sc_hd__mux2_1
Xhold817 control.body\[675\] vssd1 vssd1 vccd1 vccd1 net2379 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap536 _01715_ vssd1 vssd1 vccd1 vccd1 net536 sky130_fd_sc_hd__buf_1
XFILLER_0_3_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold828 control.body\[914\] vssd1 vssd1 vccd1 vccd1 net2390 sky130_fd_sc_hd__dlygate4sd3_1
X_13319_ net229 net316 _07495_ _07841_ net1733 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[435\]
+ sky130_fd_sc_hd__a32o_1
X_17087_ ag2.body\[193\] net731 net725 ag2.body\[194\] _02765_ vssd1 vssd1 vccd1 vccd1
+ _02766_ sky130_fd_sc_hd__o221a_1
Xhold839 control.body\[839\] vssd1 vssd1 vccd1 vccd1 net2401 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__15134__A2 net107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14299_ net808 ag2.body\[221\] ag2.body\[220\] net814 vssd1 vssd1 vccd1 vccd1 _08460_
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_42_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16038_ net709 net948 net939 net930 vssd1 vssd1 vccd1 vccd1 _01717_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_111_3695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_1047 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18084__A1 net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16095__B1 net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17989_ net45 _03606_ vssd1 vssd1 vccd1 vccd1 _03607_ sky130_fd_sc_hd__nor2_1
XANTENNA__14645__A1 net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15842__B1 _01644_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14645__B2 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19728_ clknet_leaf_133_clk _00672_ net1305 vssd1 vssd1 vccd1 vccd1 control.body\[670\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13017__B net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19659_ clknet_leaf_119_clk _00603_ net1391 vssd1 vssd1 vccd1 vccd1 control.body\[729\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__18096__A net44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18974__CLK clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09412_ img_gen.updater.commands.mode\[1\] net687 _04389_ vssd1 vssd1 vccd1 vccd1
+ _04392_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_71_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09343_ sound_gen.osc1.stayCount\[16\] sound_gen.osc1.stayCount\[14\] sound_gen.osc1.stayCount\[10\]
+ sound_gen.osc1.stayCount\[9\] vssd1 vssd1 vccd1 vccd1 _04347_ sky130_fd_sc_hd__and4_1
XFILLER_0_34_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout241_A net242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout339_A net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09274_ sound_gen.osc1.stayCount\[15\] net535 _04295_ _04296_ sound_gen.osc1.stayCount\[17\]
+ vssd1 vssd1 vccd1 vccd1 _04297_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_90_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10376__B net1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20503_ clknet_leaf_23_clk _01390_ net1359 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[139\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_74_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1150_A net1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1369 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout127_X net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout506_A net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1248_A net1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20434_ clknet_leaf_23_clk _01321_ net1358 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[70\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_47_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17159__B net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11488__A net1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11934__A2 net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20365_ clknet_leaf_21_clk _01252_ net1360 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__10392__A net1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1415_A net1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1036_X net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16998__B net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_1392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20296_ clknet_leaf_36_clk control.divider.next_count\[17\] net1351 vssd1 vssd1 vccd1
+ vccd1 control.divider.count\[17\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_100_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14799__A net1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout496_X net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout875_A net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1203_X net1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input1_X net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11935__B net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15407__B net52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08989_ ag2.body\[86\] vssd1 vssd1 vccd1 vccd1 _04014_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout663_X net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14636__A1 net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14636__B2 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17903__A net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13208__A _07624_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10353__A_N ag2.body\[288\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12111__A2 net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout830_X net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10951_ ag2.body\[175\] net1056 vssd1 vssd1 vccd1 vccd1 _05924_ sky130_fd_sc_hd__xor2_1
XFILLER_0_98_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout928_X net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17050__A2 net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1075 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13670_ _04239_ _04402_ vssd1 vssd1 vccd1 vccd1 _08019_ sky130_fd_sc_hd__nand2_1
X_10882_ _05844_ _05849_ _05854_ _05304_ vssd1 vssd1 vccd1 vccd1 _05855_ sky130_fd_sc_hd__or4b_2
XFILLER_0_112_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12621_ net307 _07512_ vssd1 vssd1 vccd1 vccd1 _07513_ sky130_fd_sc_hd__nor2_1
XFILLER_0_66_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09815__B2 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_125_Right_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15340_ net2612 net71 _01590_ net2283 vssd1 vssd1 vccd1 vccd1 _00637_ sky130_fd_sc_hd__a22o_1
XFILLER_0_66_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11622__A1 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12552_ net285 net334 _07444_ _07471_ _07474_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[35\]
+ sky130_fd_sc_hd__a41o_1
XANTENNA__17889__A1 _08141_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10286__B net1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1171 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11503_ net1199 net1225 vssd1 vssd1 vccd1 vccd1 _06476_ sky130_fd_sc_hd__nand2b_4
XFILLER_0_19_581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15271_ control.body\[766\] net108 _01582_ net2257 vssd1 vssd1 vccd1 vccd1 _00576_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__16561__A1 net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12483_ net338 _07434_ vssd1 vssd1 vccd1 vccd1 _07435_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_134_4396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17010_ ag2.body\[500\] net712 net706 ag2.body\[501\] _02688_ vssd1 vssd1 vccd1 vccd1
+ _02689_ sky130_fd_sc_hd__a221o_1
XFILLER_0_0_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14222_ _08379_ _08380_ _08381_ _08382_ vssd1 vssd1 vccd1 vccd1 _08383_ sky130_fd_sc_hd__nand4b_1
XFILLER_0_11_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13375__A1 net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11434_ ag2.body\[397\] net1113 vssd1 vssd1 vccd1 vccd1 _06407_ sky130_fd_sc_hd__xor2_1
XANTENNA__17069__B net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_893 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11925__A2 net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14153_ _08307_ _08308_ _08310_ vssd1 vssd1 vccd1 vccd1 _08314_ sky130_fd_sc_hd__and3_1
X_11365_ net1099 control.body\[813\] vssd1 vssd1 vccd1 vccd1 _06338_ sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_100_clk clknet_4_11__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_100_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_104_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_1323 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18847__CLK clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13104_ net291 _07742_ _07743_ net1946 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[317\]
+ sky130_fd_sc_hd__a22o_1
X_10316_ ag2.body\[611\] net1147 vssd1 vssd1 vccd1 vccd1 _05289_ sky130_fd_sc_hd__xor2_1
XANTENNA__16864__A2 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18961_ clknet_leaf_7_clk img_gen.tracker.next_frame\[399\] net1266 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[399\] sky130_fd_sc_hd__dfrtp_1
X_14084_ _08244_ _08240_ _08243_ vssd1 vssd1 vccd1 vccd1 _08245_ sky130_fd_sc_hd__or3b_1
XFILLER_0_123_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11296_ net1145 control.body\[683\] vssd1 vssd1 vccd1 vccd1 _06269_ sky130_fd_sc_hd__xor2_1
XANTENNA__12006__B net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1480 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1378 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17912_ net355 _03542_ net298 vssd1 vssd1 vccd1 vccd1 _03547_ sky130_fd_sc_hd__and3_1
X_13035_ _07712_ net262 _07710_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[280\]
+ sky130_fd_sc_hd__mux2_1
X_10247_ ag2.body\[322\] net1186 vssd1 vssd1 vccd1 vccd1 _05220_ sky130_fd_sc_hd__xor2_1
X_18892_ clknet_leaf_26_clk img_gen.tracker.next_frame\[330\] net1342 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[330\] sky130_fd_sc_hd__dfrtp_1
Xfanout1120 net1121 vssd1 vssd1 vccd1 vccd1 net1120 sky130_fd_sc_hd__buf_4
Xfanout1131 net1132 vssd1 vssd1 vccd1 vccd1 net1131 sky130_fd_sc_hd__clkbuf_4
Xfanout1142 net1143 vssd1 vssd1 vccd1 vccd1 net1142 sky130_fd_sc_hd__clkbuf_4
X_17843_ _07304_ _07316_ _03498_ vssd1 vssd1 vccd1 vccd1 _03499_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_20_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_8_clk_X clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10178_ _05147_ _05148_ _05149_ _05150_ vssd1 vssd1 vccd1 vccd1 _05151_ sky130_fd_sc_hd__or4_2
Xfanout1153 net1156 vssd1 vssd1 vccd1 vccd1 net1153 sky130_fd_sc_hd__clkbuf_4
XANTENNA__15824__B1 _01643_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1164 net1166 vssd1 vssd1 vccd1 vccd1 net1164 sky130_fd_sc_hd__clkbuf_8
Xfanout1175 net1178 vssd1 vssd1 vccd1 vccd1 net1175 sky130_fd_sc_hd__clkbuf_4
Xfanout1186 net1188 vssd1 vssd1 vccd1 vccd1 net1186 sky130_fd_sc_hd__buf_4
X_17774_ _03440_ _03442_ _03445_ _03452_ vssd1 vssd1 vccd1 vccd1 _03453_ sky130_fd_sc_hd__and4_1
Xfanout1197 net1198 vssd1 vssd1 vccd1 vccd1 net1197 sky130_fd_sc_hd__buf_4
X_14986_ net2643 net151 _01549_ control.body\[1001\] vssd1 vssd1 vccd1 vccd1 _00323_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__09503__B1 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19513_ clknet_leaf_121_clk _00457_ net1403 vssd1 vssd1 vccd1 vccd1 control.body\[887\]
+ sky130_fd_sc_hd__dfrtp_1
X_16725_ obsg2.obstacleArray\[119\] net501 net492 obsg2.obstacleArray\[116\] vssd1
+ vssd1 vccd1 vccd1 _02404_ sky130_fd_sc_hd__a22o_1
X_13937_ _04862_ net61 vssd1 vssd1 vccd1 vccd1 _08154_ sky130_fd_sc_hd__nor2_2
XFILLER_0_88_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17532__B net965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13850__A2 net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17041__A2 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19444_ clknet_leaf_109_clk _00388_ net1420 vssd1 vssd1 vccd1 vccd1 control.body\[946\]
+ sky130_fd_sc_hd__dfrtp_1
X_16656_ obsg2.obstacleArray\[9\] net449 vssd1 vssd1 vccd1 vccd1 _02335_ sky130_fd_sc_hd__or2_1
X_13868_ _04639_ _04642_ _08141_ _08028_ vssd1 vssd1 vccd1 vccd1 _08142_ sky130_fd_sc_hd__a31o_1
XFILLER_0_53_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_1463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15607_ ag2.body\[456\] net121 _01620_ ag2.body\[448\] vssd1 vssd1 vccd1 vccd1 _00874_
+ sky130_fd_sc_hd__a22o_1
X_12819_ net232 _07610_ _07611_ net1667 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[165\]
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_100_3363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19375_ clknet_leaf_93_clk _00319_ net1436 vssd1 vssd1 vccd1 vccd1 control.body\[1021\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_100_3374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16587_ net392 _02263_ _02265_ net362 vssd1 vssd1 vccd1 vccd1 _02266_ sky130_fd_sc_hd__a211o_1
X_13799_ _07178_ net465 vssd1 vssd1 vccd1 vccd1 _08103_ sky130_fd_sc_hd__and2_1
XFILLER_0_31_1413 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_3385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18326_ _04944_ _05697_ _08025_ vssd1 vssd1 vccd1 vccd1 _03822_ sky130_fd_sc_hd__a21o_1
XFILLER_0_84_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15538_ ag2.body\[524\] net160 _01611_ ag2.body\[516\] vssd1 vssd1 vccd1 vccd1 _00814_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__10196__B net1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18257_ obsg2.obstacleArray\[125\] _03767_ net526 vssd1 vssd1 vccd1 vccd1 _01376_
+ sky130_fd_sc_hd__o21a_1
X_15469_ ag2.body\[591\] net110 _01603_ ag2.body\[583\] vssd1 vssd1 vccd1 vccd1 _00753_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12692__A net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_117_3882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17208_ ag2.body\[52\] net959 vssd1 vssd1 vccd1 vccd1 _02887_ sky130_fd_sc_hd__nand2_1
XFILLER_0_71_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_3893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_236 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18188_ _03631_ net41 vssd1 vssd1 vccd1 vccd1 _03733_ sky130_fd_sc_hd__nor2_1
XFILLER_0_114_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_113_3757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold603 img_gen.tracker.frame\[24\] vssd1 vssd1 vccd1 vccd1 net2165 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_113_3768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_113_3779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17139_ ag2.body\[265\] net873 vssd1 vssd1 vccd1 vccd1 _02818_ sky130_fd_sc_hd__xnor2_1
Xhold614 control.body\[813\] vssd1 vssd1 vccd1 vccd1 net2176 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold625 _00237_ vssd1 vssd1 vccd1 vccd1 net2187 sky130_fd_sc_hd__dlygate4sd3_1
Xhold636 img_gen.updater.commands.rR1.rainbowRNG\[13\] vssd1 vssd1 vccd1 vccd1 net2198
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold647 control.body\[970\] vssd1 vssd1 vccd1 vccd1 net2209 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold658 control.body\[959\] vssd1 vssd1 vccd1 vccd1 net2220 sky130_fd_sc_hd__dlygate4sd3_1
X_20150_ clknet_leaf_96_clk _01094_ net1449 vssd1 vssd1 vccd1 vccd1 ag2.body\[244\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_122_291 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09961_ ag2.body\[86\] net1088 vssd1 vssd1 vccd1 vccd1 _04934_ sky130_fd_sc_hd__nand2_1
XANTENNA__19772__CLK clknet_leaf_127_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17707__B net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold669 _00640_ vssd1 vssd1 vccd1 vccd1 net2231 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_1407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkload26_A clknet_leaf_131_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20081_ clknet_leaf_77_clk _01025_ net1490 vssd1 vssd1 vccd1 vccd1 ag2.body\[319\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_102_1429 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09892_ ag2.body\[76\] net1143 vssd1 vssd1 vccd1 vccd1 _04865_ sky130_fd_sc_hd__nand2_1
XANTENNA__12877__B1 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15227__B net53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout191_A net192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14618__A1 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14618__B2 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17280__A2 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_0_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17442__B net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17568__B1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout456_A net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20588__1520 vssd1 vssd1 vccd1 vccd1 _20588__1520/HI net1520 sky130_fd_sc_hd__conb_1
XANTENNA__17032__A2 net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1198_A net1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19152__CLK clknet_leaf_52_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11852__A1 net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12586__B net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16058__B net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09241__A net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11490__B net1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16773__S net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_2779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout623_A net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09326_ net1587 _04337_ vssd1 vssd1 vccd1 vccd1 _01434_ sky130_fd_sc_hd__xor2_1
XFILLER_0_36_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11604__A1 net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_838 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13698__A net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09895__B net1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09257_ ssdec1.in\[3\] vssd1 vssd1 vccd1 vccd1 _04282_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout411_X net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17740__B1 _02491_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1153_X net1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09188_ ag2.body\[585\] vssd1 vssd1 vccd1 vccd1 _04213_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout992_A net995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10834__B net1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_1480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11907__A2 net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20417_ clknet_leaf_34_clk _01304_ net1357 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[53\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__17099__A2 net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13109__A1 net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16846__A2 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11150_ ag2.body\[604\] net1120 vssd1 vssd1 vccd1 vccd1 _06123_ sky130_fd_sc_hd__xor2_1
XFILLER_0_101_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20348_ clknet_leaf_139_clk _01239_ net1292 vssd1 vssd1 vccd1 vccd1 img_gen.updater.commands.rR1.rainbowRNG\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout780_X net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19211__RESET_B net1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout878_X net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10101_ net911 net919 net915 vssd1 vssd1 vccd1 vccd1 _05074_ sky130_fd_sc_hd__or3b_4
XFILLER_0_105_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11081_ ag2.body\[540\] net1132 vssd1 vssd1 vccd1 vccd1 _06054_ sky130_fd_sc_hd__or2_1
XFILLER_0_60_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20279_ clknet_leaf_35_clk control.divider.next_count\[0\] net1348 vssd1 vssd1 vccd1
+ vccd1 control.divider.count\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_41_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16059__B1 net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10032_ ag2.body\[505\] net1210 vssd1 vssd1 vccd1 vccd1 _05005_ sky130_fd_sc_hd__nand2_1
XANTENNA__17904__Y _03539_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14609__A1 net1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14609__B2 net822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15806__B1 _01641_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17633__A ag2.body\[164\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14840_ _08889_ _08895_ _08753_ vssd1 vssd1 vccd1 vccd1 _01511_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_51_1871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_51_1882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14771_ net976 _04024_ _04025_ net1030 _08926_ vssd1 vssd1 vccd1 vccd1 _08932_ sky130_fd_sc_hd__a221o_1
XANTENNA__17559__B1 net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11983_ img_gen.tracker.frame\[532\] net596 net541 img_gen.tracker.frame\[535\] vssd1
+ vssd1 vccd1 vccd1 _06955_ sky130_fd_sc_hd__o22a_1
XANTENNA__16249__A net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13832__A2 net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16510_ obsg2.obstacleArray\[6\] obsg2.obstacleArray\[7\] net456 vssd1 vssd1 vccd1
+ vccd1 _02189_ sky130_fd_sc_hd__mux2_1
X_13722_ net26 net25 vssd1 vssd1 vccd1 vccd1 toggle1.nextBlinkToggle\[1\] sky130_fd_sc_hd__and2b_1
XFILLER_0_98_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10934_ _05900_ _05902_ _05904_ _05906_ vssd1 vssd1 vccd1 vccd1 _05907_ sky130_fd_sc_hd__and4_2
X_17490_ _03165_ _03166_ _03168_ vssd1 vssd1 vccd1 vccd1 _03169_ sky130_fd_sc_hd__or3b_1
XFILLER_0_98_598 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16231__B1 net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12496__B net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13653_ _08009_ vssd1 vssd1 vccd1 vccd1 _08010_ sky130_fd_sc_hd__inv_2
X_16441_ _02116_ _02118_ _02119_ net365 vssd1 vssd1 vccd1 vccd1 _02120_ sky130_fd_sc_hd__a22o_1
X_10865_ _05752_ _05781_ _05812_ _05837_ vssd1 vssd1 vccd1 vccd1 _05838_ sky130_fd_sc_hd__and4_1
XANTENNA__16782__A1 net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_136_4458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12604_ net231 _07503_ _07504_ net1966 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[57\]
+ sky130_fd_sc_hd__a22o_1
X_16372_ _01896_ _02030_ _02049_ _02050_ _01895_ vssd1 vssd1 vccd1 vccd1 _02051_ sky130_fd_sc_hd__o221a_1
X_19160_ clknet_leaf_112_clk _00104_ net1403 vssd1 vssd1 vccd1 vccd1 toggle1.bcd_hundreds\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_136_4469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13584_ control.divider.count\[4\] _07958_ vssd1 vssd1 vccd1 vccd1 _07959_ sky130_fd_sc_hd__and2_1
XFILLER_0_82_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10796_ ag2.body\[38\] net1078 vssd1 vssd1 vccd1 vccd1 _05769_ sky130_fd_sc_hd__or2_1
XFILLER_0_27_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_45_1686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18111_ net44 _03689_ vssd1 vssd1 vccd1 vccd1 _03690_ sky130_fd_sc_hd__nor2_1
XFILLER_0_93_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15323_ control.body\[715\] net73 _01589_ net2548 vssd1 vssd1 vccd1 vccd1 _00621_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_45_1697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12535_ net2084 net652 _07465_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[27\]
+ sky130_fd_sc_hd__and3_1
XANTENNA__10584__X _05557_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19091_ clknet_leaf_0_clk img_gen.tracker.next_frame\[529\] net1239 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[529\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_129_1510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18042_ obsg2.obstacleArray\[33\] _03644_ net521 vssd1 vssd1 vccd1 vccd1 _01284_
+ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_10_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_1490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15254_ net2113 net109 net50 net2382 vssd1 vssd1 vccd1 vccd1 _00562_ sky130_fd_sc_hd__a22o_1
XFILLER_0_53_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19795__CLK clknet_leaf_124_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12466_ net611 net469 net561 _07312_ vssd1 vssd1 vccd1 vccd1 _07421_ sky130_fd_sc_hd__and4_1
XFILLER_0_53_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14205_ net843 ag2.body\[360\] ag2.body\[366\] net801 _08360_ vssd1 vssd1 vccd1 vccd1
+ _08366_ sky130_fd_sc_hd__a221o_1
XFILLER_0_22_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11417_ _06386_ _06387_ _06388_ _06389_ _06385_ vssd1 vssd1 vccd1 vccd1 _06390_ sky130_fd_sc_hd__a221o_1
X_15185_ control.body\[834\] net101 _01572_ net2484 vssd1 vssd1 vccd1 vccd1 _00500_
+ sky130_fd_sc_hd__a22o_1
X_12397_ net625 net588 _07292_ _07296_ vssd1 vssd1 vccd1 vccd1 _07361_ sky130_fd_sc_hd__and4_1
XANTENNA__10031__B1 net1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14136_ net972 ag2.body\[171\] vssd1 vssd1 vccd1 vccd1 _08297_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_91_3086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16837__A2 net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09972__B1 net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11348_ ag2.body\[443\] net1153 vssd1 vssd1 vccd1 vccd1 _06321_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_91_3097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19993_ clknet_leaf_66_clk _00937_ net1475 vssd1 vssd1 vccd1 vccd1 ag2.body\[407\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_103_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14848__A1 _08768_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14067_ net991 ag2.body\[209\] vssd1 vssd1 vccd1 vccd1 _08228_ sky130_fd_sc_hd__xnor2_1
X_18944_ clknet_leaf_139_clk img_gen.tracker.next_frame\[382\] net1290 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[382\] sky130_fd_sc_hd__dfrtp_1
X_11279_ _06241_ _06247_ _06248_ _06250_ vssd1 vssd1 vccd1 vccd1 _06252_ sky130_fd_sc_hd__or4_1
XANTENNA__10760__A net1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13018_ _07704_ net262 _07702_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[271\]
+ sky130_fd_sc_hd__mux2_1
X_18875_ clknet_leaf_13_clk img_gen.tracker.next_frame\[313\] net1282 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[313\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_1384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14567__A1_N net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17826_ net840 net224 vssd1 vssd1 vccd1 vccd1 _03490_ sky130_fd_sc_hd__nor2_1
XANTENNA__19175__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_106_3550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_3561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09613__X _04586_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17757_ _01742_ _03400_ _03402_ net349 net350 vssd1 vssd1 vccd1 vccd1 _03436_ sky130_fd_sc_hd__o2111a_1
XANTENNA__17262__B net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14969_ net2502 net157 net51 control.body\[1019\] vssd1 vssd1 vccd1 vccd1 _00309_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12687__A net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_3425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_3436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_3447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16708_ obsg2.obstacleArray\[79\] net500 net486 obsg2.obstacleArray\[78\] vssd1 vssd1
+ vccd1 vccd1 _02387_ sky130_fd_sc_hd__a22o_1
XFILLER_0_77_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17688_ ag2.body\[155\] net855 vssd1 vssd1 vccd1 vccd1 _03367_ sky130_fd_sc_hd__or2_1
XANTENNA__10919__B net1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_306 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15998__A net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19427_ clknet_leaf_107_clk _00371_ net1434 vssd1 vssd1 vccd1 vccd1 control.body\[961\]
+ sky130_fd_sc_hd__dfrtp_1
X_16639_ obsg2.obstacleArray\[52\] obsg2.obstacleArray\[53\] net444 vssd1 vssd1 vccd1
+ vccd1 _02318_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16593__S net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15576__A2 net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09996__A net1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_119_3944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19358_ clknet_leaf_101_clk _00302_ net1438 vssd1 vssd1 vccd1 vccd1 control.body\[1036\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_128_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_119_3955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_119_3966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09111_ ag2.body\[380\] vssd1 vssd1 vccd1 vccd1 _04136_ sky130_fd_sc_hd__inv_2
XFILLER_0_57_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18309_ track.nextHighScore\[1\] _03787_ net321 net323 vssd1 vssd1 vccd1 vccd1 _03805_
+ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_115_3819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19289_ clknet_leaf_98_clk net2271 net1446 vssd1 vssd1 vccd1 vccd1 control.body\[1111\]
+ sky130_fd_sc_hd__dfrtp_1
X_09042_ ag2.body\[207\] vssd1 vssd1 vccd1 vccd1 _04067_ sky130_fd_sc_hd__inv_2
XFILLER_0_44_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13311__A net225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10654__B net1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18278__A1 net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold400 img_gen.tracker.frame\[460\] vssd1 vssd1 vccd1 vccd1 net1962 sky130_fd_sc_hd__dlygate4sd3_1
Xhold411 img_gen.tracker.frame\[457\] vssd1 vssd1 vccd1 vccd1 net1973 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout204_A net218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold422 img_gen.tracker.frame\[157\] vssd1 vssd1 vccd1 vccd1 net1984 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10373__C net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20202_ clknet_leaf_55_clk _01146_ net1456 vssd1 vssd1 vccd1 vccd1 ag2.body\[184\]
+ sky130_fd_sc_hd__dfrtp_4
Xhold433 img_gen.tracker.frame\[151\] vssd1 vssd1 vccd1 vccd1 net1995 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09963__B1 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold444 img_gen.tracker.frame\[112\] vssd1 vssd1 vccd1 vccd1 net2006 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__16828__A2 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_2572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold455 img_gen.tracker.frame\[267\] vssd1 vssd1 vccd1 vccd1 net2017 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold466 img_gen.tracker.frame\[149\] vssd1 vssd1 vccd1 vccd1 net2028 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold477 img_gen.tracker.frame\[261\] vssd1 vssd1 vccd1 vccd1 net2039 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11770__B1 net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold488 img_gen.tracker.frame\[156\] vssd1 vssd1 vccd1 vccd1 net2050 sky130_fd_sc_hd__dlygate4sd3_1
X_09944_ net1048 control.body\[743\] vssd1 vssd1 vccd1 vccd1 _04917_ sky130_fd_sc_hd__xor2_1
Xfanout902 control.body_update.curr_length\[5\] vssd1 vssd1 vccd1 vccd1 net902 sky130_fd_sc_hd__clkbuf_4
X_20133_ clknet_leaf_80_clk _01077_ net1449 vssd1 vssd1 vccd1 vccd1 ag2.body\[259\]
+ sky130_fd_sc_hd__dfrtp_2
Xhold499 control.body\[753\] vssd1 vssd1 vccd1 vccd1 net2061 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout913 net915 vssd1 vssd1 vccd1 vccd1 net913 sky130_fd_sc_hd__buf_4
XANTENNA__15500__A2 net113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_2447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1113_A net1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_70_2458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout924 ag2.body\[6\] vssd1 vssd1 vccd1 vccd1 net924 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_70_2469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout935 net936 vssd1 vssd1 vccd1 vccd1 net935 sky130_fd_sc_hd__buf_4
X_20064_ clknet_leaf_72_clk _01008_ net1502 vssd1 vssd1 vccd1 vccd1 ag2.body\[334\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_102_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout946 net947 vssd1 vssd1 vccd1 vccd1 net946 sky130_fd_sc_hd__buf_4
Xfanout957 net958 vssd1 vssd1 vccd1 vccd1 net957 sky130_fd_sc_hd__clkbuf_4
X_09875_ ag2.body\[163\] net1154 vssd1 vssd1 vccd1 vccd1 _04848_ sky130_fd_sc_hd__or2_1
XANTENNA_input9_A nrst vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout968 obsg2.randCord\[4\] vssd1 vssd1 vccd1 vccd1 net968 sky130_fd_sc_hd__buf_4
XANTENNA__16768__S net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1100 control.body\[895\] vssd1 vssd1 vccd1 vccd1 net2662 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout573_A _06649_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout979 net980 vssd1 vssd1 vccd1 vccd1 net979 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_5_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_2966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_2977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout740_A net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout361_X net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_2988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1482_A net1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19668__CLK clknet_leaf_118_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout459_X net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_2387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout838_A net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09242__Y _04267_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_2398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_1300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10829__B net1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout626_X net626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1368_X net1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10650_ ag2.body\[280\] net1237 vssd1 vssd1 vccd1 vccd1 _05623_ sky130_fd_sc_hd__or2_1
XFILLER_0_48_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09309_ sound_gen.osc1.count\[7\] net272 _04319_ _04328_ vssd1 vssd1 vccd1 vccd1
+ _01442_ sky130_fd_sc_hd__a22o_1
XFILLER_0_64_955 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_4311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10581_ ag2.body\[185\] net1208 vssd1 vssd1 vccd1 vccd1 _05554_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_131_4322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_4333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11530__C_N _06497_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12320_ _07242_ _07286_ vssd1 vssd1 vccd1 vccd1 _07287_ sky130_fd_sc_hd__nand2_2
XFILLER_0_134_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_40_1550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout995_X net995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10564__B net1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12251_ img_gen.updater.commands.cmd_num\[0\] _07187_ _07219_ _07220_ vssd1 vssd1
+ vccd1 vccd1 _07221_ sky130_fd_sc_hd__o22a_2
X_11202_ control.body\[876\] net1131 vssd1 vssd1 vccd1 vccd1 _06175_ sky130_fd_sc_hd__nand2b_1
XANTENNA__16819__A2 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12182_ net1197 ag2.apple_cord\[1\] vssd1 vssd1 vccd1 vccd1 _07154_ sky130_fd_sc_hd__nand2_1
XFILLER_0_82_1185 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_129_4251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11761__B1 net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11133_ net1051 control.body\[871\] vssd1 vssd1 vccd1 vccd1 _06106_ sky130_fd_sc_hd__xnor2_1
XANTENNA__11676__A _06639_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_4262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17492__A2 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16990_ ag2.body\[88\] net739 net953 _04020_ vssd1 vssd1 vccd1 vccd1 _02669_ sky130_fd_sc_hd__a22o_1
XANTENNA__19198__CLK clknet_leaf_53_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_53_1933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13502__A1 net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_1490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09146__A ag2.body\[478\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11064_ ag2.body\[434\] net1176 vssd1 vssd1 vccd1 vccd1 _06037_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_125_4148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15941_ ag2.body\[163\] net195 _01653_ ag2.body\[155\] vssd1 vssd1 vccd1 vccd1 _01173_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_95_1502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_34_1354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_34_1365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10015_ ag2.body\[270\] net1091 vssd1 vssd1 vccd1 vccd1 _04988_ sky130_fd_sc_hd__xor2_1
X_18660_ clknet_leaf_5_clk img_gen.tracker.next_frame\[98\] net1276 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[98\] sky130_fd_sc_hd__dfrtp_1
X_15872_ ag2.body\[230\] net201 _01647_ ag2.body\[222\] vssd1 vssd1 vccd1 vccd1 _01112_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_30_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16452__B1 net367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18178__B net41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17611_ ag2.body\[605\] net946 vssd1 vssd1 vccd1 vccd1 _03290_ sky130_fd_sc_hd__xor2_1
X_14823_ net994 _04044_ ag2.body\[156\] net815 _01493_ vssd1 vssd1 vccd1 vccd1 _01494_
+ sky130_fd_sc_hd__a221o_1
XANTENNA__17082__B net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18591_ clknet_leaf_14_clk img_gen.tracker.next_frame\[29\] net1280 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[29\] sky130_fd_sc_hd__dfrtp_1
X_17542_ ag2.body\[322\] net866 vssd1 vssd1 vccd1 vccd1 _03221_ sky130_fd_sc_hd__xor2_1
XFILLER_0_114_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11966_ net560 _06937_ _06935_ vssd1 vssd1 vccd1 vccd1 _06938_ sky130_fd_sc_hd__a21o_1
X_14754_ net979 ag2.body\[42\] vssd1 vssd1 vccd1 vccd1 _08915_ sky130_fd_sc_hd__xor2_1
XFILLER_0_98_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10739__B net1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10917_ _05886_ _05887_ _05888_ _05889_ vssd1 vssd1 vccd1 vccd1 _05890_ sky130_fd_sc_hd__and4_2
X_13705_ _04283_ _08027_ _08043_ _08044_ _08045_ vssd1 vssd1 vccd1 vccd1 _08046_ sky130_fd_sc_hd__a221oi_1
XTAP_TAPCELL_ROW_47_1748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17473_ ag2.body\[133\] net953 vssd1 vssd1 vccd1 vccd1 _03152_ sky130_fd_sc_hd__nand2_1
X_14685_ net1032 _04020_ ag2.body\[95\] net794 vssd1 vssd1 vccd1 vccd1 _08846_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_47_1759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18194__A _01703_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11897_ img_gen.tracker.frame\[64\] net596 net541 img_gen.tracker.frame\[67\] _06868_
+ vssd1 vssd1 vccd1 vccd1 _06869_ sky130_fd_sc_hd__o221a_1
XFILLER_0_132_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19212_ clknet_leaf_57_clk _00156_ net1477 vssd1 vssd1 vccd1 vccd1 ag2.body\[75\]
+ sky130_fd_sc_hd__dfrtp_2
X_13636_ _07997_ _07998_ vssd1 vssd1 vccd1 vccd1 control.divider.next_count\[12\]
+ sky130_fd_sc_hd__nor2_1
X_16424_ _02074_ _02100_ _02076_ vssd1 vssd1 vccd1 vccd1 _02103_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_28_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10848_ ag2.body\[40\] net1219 vssd1 vssd1 vccd1 vccd1 _05821_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_15_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1499 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_15_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19143_ clknet_leaf_132_clk net1579 net1303 vssd1 vssd1 vccd1 vccd1 img_gen.control.detect4.Q\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_16355_ net420 _02033_ _02032_ net372 vssd1 vssd1 vccd1 vccd1 _02034_ sky130_fd_sc_hd__a211o_1
XFILLER_0_82_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13567_ _07933_ _07939_ _07944_ _07938_ vssd1 vssd1 vccd1 vccd1 _07946_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_26_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_97_3273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10755__A net1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10779_ _05740_ _05751_ _05633_ _05739_ vssd1 vssd1 vccd1 vccd1 _05752_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_82_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_843 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_3284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_3295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15306_ control.body\[733\] net75 _01586_ net2464 vssd1 vssd1 vccd1 vccd1 _00607_
+ sky130_fd_sc_hd__a22o_1
X_12518_ img_gen.tracker.frame\[20\] net649 _07455_ vssd1 vssd1 vccd1 vccd1 _07456_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_67_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16286_ obsg2.obstacleArray\[124\] obsg2.obstacleArray\[125\] net407 vssd1 vssd1
+ vccd1 vccd1 _01965_ sky130_fd_sc_hd__mux2_1
X_19074_ clknet_leaf_28_clk img_gen.tracker.next_frame\[512\] net1335 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[512\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_48_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_93_3148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13498_ net250 _07910_ _07911_ net1757 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[544\]
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_93_3159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18025_ net432 _01713_ net491 vssd1 vssd1 vccd1 vccd1 _03633_ sky130_fd_sc_hd__and3_1
X_12449_ img_gen.updater.commands.rR1.rainbowRNG\[7\] net248 _07377_ vssd1 vssd1 vccd1
+ vccd1 _07409_ sky130_fd_sc_hd__a21o_1
X_15237_ net2507 net98 _01578_ control.body\[776\] vssd1 vssd1 vccd1 vccd1 _00546_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12970__A net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15168_ control.body\[851\] net95 _01570_ control.body\[843\] vssd1 vssd1 vccd1 vccd1
+ _00485_ sky130_fd_sc_hd__a22o_1
XANTENNA__11752__B1 _06722_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14119_ _08273_ _08277_ _08278_ _08279_ vssd1 vssd1 vccd1 vccd1 _08280_ sky130_fd_sc_hd__or4_4
XANTENNA__17483__A2 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19976_ clknet_leaf_63_clk _00920_ net1470 vssd1 vssd1 vccd1 vccd1 ag2.body\[422\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_120_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout209 net210 vssd1 vssd1 vccd1 vccd1 net209 sky130_fd_sc_hd__buf_2
X_15099_ net2196 net148 _01563_ net2481 vssd1 vssd1 vccd1 vccd1 _00423_ sky130_fd_sc_hd__a22o_1
XFILLER_0_61_1269 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_3612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18927_ clknet_leaf_140_clk img_gen.tracker.next_frame\[365\] net1290 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[365\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_108_3623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18565__CLK clknet_leaf_15_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17235__A2 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09660_ control.body_update.curr_length\[6\] net902 net911 net906 vssd1 vssd1 vccd1
+ vccd1 _04633_ sky130_fd_sc_hd__nor4_1
XFILLER_0_59_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18858_ clknet_leaf_18_clk img_gen.tracker.next_frame\[296\] net1323 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[296\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_104_3509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17809_ net925 _08124_ vssd1 vssd1 vccd1 vccd1 _03477_ sky130_fd_sc_hd__nand2_1
X_09591_ net1107 control.body\[909\] vssd1 vssd1 vccd1 vccd1 _04564_ sky130_fd_sc_hd__xor2_1
XANTENNA__10489__X _05462_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18789_ clknet_leaf_13_clk img_gen.tracker.next_frame\[227\] net1284 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[227\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_136_1355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_2830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10649__B net1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkload93_A clknet_leaf_111_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19974__RESET_B net1470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12480__A1 net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_2240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_2251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout154_A net183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19903__RESET_B net1464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_1517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16210__A3 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_367 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10665__A net1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14137__A net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1063_A net1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_76_2634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09025_ ag2.body\[161\] vssd1 vssd1 vccd1 vccd1 _04050_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_76_2645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11991__B1 net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_2656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20461__RESET_B net1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16352__A obsg2.obstacleArray\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1230_A net1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_2509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_2055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19340__CLK clknet_leaf_103_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_2066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold230 img_gen.tracker.frame\[221\] vssd1 vssd1 vccd1 vccd1 net1792 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13695__B net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold241 img_gen.tracker.frame\[228\] vssd1 vssd1 vccd1 vccd1 net1803 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout690_A net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold252 img_gen.tracker.frame\[406\] vssd1 vssd1 vccd1 vccd1 net1814 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11743__B1 net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout788_A net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18908__CLK clknet_leaf_144_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold263 img_gen.tracker.frame\[452\] vssd1 vssd1 vccd1 vccd1 net1825 sky130_fd_sc_hd__dlygate4sd3_1
Xhold274 img_gen.tracker.frame\[76\] vssd1 vssd1 vccd1 vccd1 net1836 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09237__Y _04262_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16131__C1 net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold285 img_gen.tracker.frame\[56\] vssd1 vssd1 vccd1 vccd1 net1847 sky130_fd_sc_hd__dlygate4sd3_1
Xhold296 img_gen.tracker.frame\[305\] vssd1 vssd1 vccd1 vccd1 net1858 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1116_X net1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout710 net714 vssd1 vssd1 vccd1 vccd1 net710 sky130_fd_sc_hd__buf_4
Xfanout721 _04265_ vssd1 vssd1 vccd1 vccd1 net721 sky130_fd_sc_hd__buf_4
XFILLER_0_102_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout732 net733 vssd1 vssd1 vccd1 vccd1 net732 sky130_fd_sc_hd__clkbuf_4
X_20116_ clknet_leaf_80_clk _01060_ net1488 vssd1 vssd1 vccd1 vccd1 ag2.body\[274\]
+ sky130_fd_sc_hd__dfrtp_4
X_09927_ _04418_ _04896_ _04897_ _04899_ _04889_ vssd1 vssd1 vccd1 vccd1 _04900_ sky130_fd_sc_hd__o41a_1
XFILLER_0_121_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout743 net744 vssd1 vssd1 vccd1 vccd1 net743 sky130_fd_sc_hd__buf_4
XANTENNA_fanout955_A obsg2.randCord\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18279__A net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout754 _04232_ vssd1 vssd1 vccd1 vccd1 net754 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout576_X net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19490__CLK clknet_leaf_113_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout765 net766 vssd1 vssd1 vccd1 vccd1 net765 sky130_fd_sc_hd__buf_4
XANTENNA__17226__A2 net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout776 _04229_ vssd1 vssd1 vccd1 vccd1 net776 sky130_fd_sc_hd__clkbuf_4
X_20047_ clknet_leaf_68_clk _00991_ net1498 vssd1 vssd1 vccd1 vccd1 ag2.body\[349\]
+ sky130_fd_sc_hd__dfrtp_4
Xfanout787 net789 vssd1 vssd1 vccd1 vccd1 net787 sky130_fd_sc_hd__clkbuf_4
X_09858_ net907 _04470_ net641 vssd1 vssd1 vccd1 vccd1 _04831_ sky130_fd_sc_hd__a21oi_4
Xfanout798 net805 vssd1 vssd1 vccd1 vccd1 net798 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout67_A _08131_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11943__B net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09789_ net1181 control.body\[946\] vssd1 vssd1 vccd1 vccd1 _04762_ sky130_fd_sc_hd__xor2_1
XANTENNA_fanout743_X net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11820_ img_gen.tracker.frame\[389\] net601 net585 img_gen.tracker.frame\[395\] _06791_
+ vssd1 vssd1 vccd1 vccd1 _06792_ sky130_fd_sc_hd__o221a_1
XFILLER_0_96_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18187__B1 net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09467__A2 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_1439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_844 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11751_ net466 _06673_ _06722_ vssd1 vssd1 vccd1 vccd1 _06723_ sky130_fd_sc_hd__a21oi_1
XANTENNA__17934__B1 net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_80_clk clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_80_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_16_1558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10702_ ag2.body\[20\] net1128 vssd1 vssd1 vccd1 vccd1 _05675_ sky130_fd_sc_hd__nand2_1
X_14470_ net838 ag2.body\[265\] ag2.body\[266\] net828 _08624_ vssd1 vssd1 vccd1 vccd1
+ _08631_ sky130_fd_sc_hd__a221o_1
XFILLER_0_7_1394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_42_1601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11682_ img_gen.tracker.frame\[143\] net585 net546 img_gen.tracker.frame\[140\] _06653_
+ vssd1 vssd1 vccd1 vccd1 _06654_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_12_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13421_ net682 _07880_ vssd1 vssd1 vccd1 vccd1 _07881_ sky130_fd_sc_hd__nor2_1
XFILLER_0_138_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10633_ net1071 control.body\[670\] vssd1 vssd1 vccd1 vccd1 _05606_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_23_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14047__A net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16140_ _01721_ _01817_ vssd1 vssd1 vccd1 vccd1 _01819_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_88_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13352_ _07519_ net304 vssd1 vssd1 vccd1 vccd1 _07854_ sky130_fd_sc_hd__nor2_1
XFILLER_0_52_947 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10564_ ag2.body\[519\] net1059 vssd1 vssd1 vccd1 vccd1 _05537_ sky130_fd_sc_hd__and2b_1
XFILLER_0_88_1394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12303_ _07218_ _07221_ vssd1 vssd1 vccd1 vccd1 _07270_ sky130_fd_sc_hd__nand2b_1
XANTENNA__11982__B1 net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16071_ _01748_ _01749_ net375 vssd1 vssd1 vccd1 vccd1 _01750_ sky130_fd_sc_hd__mux2_1
XANTENNA__15173__B1 net63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13283_ net384 _07468_ vssd1 vssd1 vccd1 vccd1 _07827_ sky130_fd_sc_hd__nor2_2
X_10495_ ag2.body\[545\] net781 net1108 _04202_ vssd1 vssd1 vccd1 vccd1 _05468_ sky130_fd_sc_hd__o22a_1
X_15022_ net2651 net166 _01555_ net2236 vssd1 vssd1 vccd1 vccd1 _00354_ sky130_fd_sc_hd__a22o_1
X_12234_ _07187_ _07203_ vssd1 vssd1 vccd1 vccd1 _07204_ sky130_fd_sc_hd__nand2_1
XANTENNA__17077__B obsg2.randCord\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11734__B1 net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19830_ clknet_leaf_122_clk _00774_ net1407 vssd1 vssd1 vccd1 vccd1 ag2.body\[564\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__16122__C1 net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12165_ net559 _07133_ _07134_ _07136_ vssd1 vssd1 vccd1 vccd1 _07137_ sky130_fd_sc_hd__a22o_1
XFILLER_0_120_1112 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18526__RESET_B net1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11116_ net786 control.body\[1096\] _04257_ net1111 _06088_ vssd1 vssd1 vccd1 vccd1
+ _06089_ sky130_fd_sc_hd__o221a_1
X_19761_ clknet_leaf_130_clk _00705_ net1316 vssd1 vssd1 vccd1 vccd1 control.body\[639\]
+ sky130_fd_sc_hd__dfrtp_1
X_16973_ _02644_ _02647_ _02650_ _02651_ vssd1 vssd1 vccd1 vccd1 _02652_ sky130_fd_sc_hd__or4_2
X_12096_ img_gen.tracker.frame\[354\] net554 _07067_ net559 vssd1 vssd1 vccd1 vccd1
+ _07068_ sky130_fd_sc_hd__a211o_1
XANTENNA__12014__B _06985_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18712_ clknet_leaf_144_clk img_gen.tracker.next_frame\[150\] net1252 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[150\] sky130_fd_sc_hd__dfrtp_1
X_11047_ ag2.body\[389\] net1104 vssd1 vssd1 vccd1 vccd1 _06020_ sky130_fd_sc_hd__xor2_1
X_15924_ ag2.body\[179\] net136 _01654_ ag2.body\[171\] vssd1 vssd1 vccd1 vccd1 _01157_
+ sky130_fd_sc_hd__a22o_1
X_19692_ clknet_leaf_136_clk _00636_ net1302 vssd1 vssd1 vccd1 vccd1 control.body\[698\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16425__B1 _02102_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12949__B net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput9 nrst vssd1 vssd1 vccd1 vccd1 net9 sky130_fd_sc_hd__buf_1
X_18643_ clknet_leaf_141_clk img_gen.tracker.next_frame\[81\] net1295 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[81\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__09604__A net1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15855_ ag2.body\[247\] net176 _01645_ ag2.body\[239\] vssd1 vssd1 vccd1 vccd1 _01097_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_56_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14806_ _01473_ _01474_ _01476_ vssd1 vssd1 vccd1 vccd1 _01477_ sky130_fd_sc_hd__and3_1
X_18574_ clknet_leaf_14_clk img_gen.tracker.next_frame\[12\] net1279 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[12\] sky130_fd_sc_hd__dfrtp_1
X_15786_ ag2.body\[296\] net208 _01639_ ag2.body\[288\] vssd1 vssd1 vccd1 vccd1 _01034_
+ sky130_fd_sc_hd__a22o_1
X_12998_ net665 _07694_ vssd1 vssd1 vccd1 vccd1 _07695_ sky130_fd_sc_hd__nor2_1
XFILLER_0_8_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17525_ ag2.body\[486\] net938 vssd1 vssd1 vccd1 vccd1 _03204_ sky130_fd_sc_hd__xor2_1
XFILLER_0_8_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14737_ net1033 ag2.body\[333\] vssd1 vssd1 vccd1 vccd1 _08898_ sky130_fd_sc_hd__xor2_1
XANTENNA__11265__A2 _06226_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11949_ img_gen.tracker.frame\[103\] net547 net561 vssd1 vssd1 vccd1 vccd1 _06921_
+ sky130_fd_sc_hd__o21a_1
Xclkbuf_leaf_71_clk clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_71_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__16437__A net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_3335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_1241 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17456_ ag2.body\[435\] net717 net690 ag2.body\[439\] vssd1 vssd1 vccd1 vccd1 _03135_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_99_3346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_99_3357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14668_ net820 ag2.body\[523\] ag2.body\[525\] net809 _08820_ vssd1 vssd1 vccd1 vccd1
+ _08829_ sky130_fd_sc_hd__o221a_1
XANTENNA__19314__RESET_B net1435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16407_ _02084_ _02085_ vssd1 vssd1 vccd1 vccd1 _02086_ sky130_fd_sc_hd__and2_1
XFILLER_0_28_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13619_ control.divider.count\[6\] _07985_ net220 vssd1 vssd1 vccd1 vccd1 _07988_
+ sky130_fd_sc_hd__o21ai_1
X_17387_ ag2.body\[490\] net728 net935 _04179_ _03065_ vssd1 vssd1 vccd1 vccd1 _03066_
+ sky130_fd_sc_hd__a221o_1
XANTENNA__15951__A2 net196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14599_ net985 _04101_ ag2.body\[311\] net796 _08757_ vssd1 vssd1 vccd1 vccd1 _08760_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_116_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19126_ clknet_leaf_131_clk img_gen.tracker.next_frame\[564\] net1295 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[564\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__19363__CLK clknet_leaf_102_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16338_ obsg2.obstacleArray\[80\] obsg2.obstacleArray\[81\] net411 vssd1 vssd1 vccd1
+ vccd1 _02017_ sky130_fd_sc_hd__mux2_1
XFILLER_0_109_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19057_ clknet_leaf_10_clk img_gen.tracker.next_frame\[495\] net1273 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[495\] sky130_fd_sc_hd__dfrtp_1
X_16269_ obsg2.obstacleArray\[30\] obsg2.obstacleArray\[31\] net411 vssd1 vssd1 vccd1
+ vccd1 _01948_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18008_ net519 _03620_ vssd1 vssd1 vccd1 vccd1 _01274_ sky130_fd_sc_hd__nor2_1
XANTENNA__09918__B1 net1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11725__B1 net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17456__A2 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19959_ clknet_leaf_44_clk _00903_ net1381 vssd1 vssd1 vccd1 vccd1 ag2.body\[437\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__18099__A net44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09712_ _04682_ _04683_ _04684_ _04681_ vssd1 vssd1 vccd1 vccd1 _04685_ sky130_fd_sc_hd__a211o_1
XANTENNA__16111__S net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09514__A net1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09643_ net775 control.body\[1018\] control.body\[1016\] net787 vssd1 vssd1 vccd1
+ vccd1 _04616_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_74_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_65_2302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_2313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17731__A _01700_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15803__X _01641_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09574_ ag2.body\[200\] net785 net747 ag2.body\[207\] _04546_ vssd1 vssd1 vccd1 vccd1
+ _04547_ sky130_fd_sc_hd__a221o_1
XANTENNA__10012__X _04985_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18169__B1 net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_1016 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1180_A net1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12875__A net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_62_clk clknet_4_13__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_62_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_clkbuf_leaf_60_clk_A clknet_4_13__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1278_A net1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_1347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_2707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15942__A2 net195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_1358 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout703_A net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1066_X net1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_459 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_2117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_2128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20596_ net1528 vssd1 vssd1 vccd1 vccd1 gpio_oeb[8] sky130_fd_sc_hd__buf_2
XANTENNA_clkbuf_leaf_75_clk_A clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10767__A1 _04238_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11964__B1 net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18730__CLK clknet_leaf_141_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1233_X net1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14154__X _08315_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09008_ ag2.body\[128\] vssd1 vssd1 vccd1 vccd1 _04033_ sky130_fd_sc_hd__inv_2
XFILLER_0_14_671 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10280_ _04433_ _04446_ _04419_ vssd1 vssd1 vccd1 vccd1 _05253_ sky130_fd_sc_hd__o21ai_4
XANTENNA__14321__A1_N net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout693_X net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10842__B net1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17906__A _03533_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20105__Q ag2.body\[295\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1505 ag2.reset vssd1 vssd1 vccd1 vccd1 net1505 sky130_fd_sc_hd__buf_8
XTAP_TAPCELL_ROW_6_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1516 net1517 vssd1 vssd1 vccd1 vccd1 net1516 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout860_X net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_133_clk_A clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout958_X net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout540 net541 vssd1 vssd1 vccd1 vccd1 net540 sky130_fd_sc_hd__buf_2
XFILLER_0_121_1476 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout551 net552 vssd1 vssd1 vccd1 vccd1 net551 sky130_fd_sc_hd__clkbuf_4
XANTENNA__14130__A1 net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14130__B2 net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout562 net567 vssd1 vssd1 vccd1 vccd1 net562 sky130_fd_sc_hd__buf_2
X_13970_ ag2.body\[109\] net202 _08157_ ag2.body\[101\] vssd1 vssd1 vccd1 vccd1 _00190_
+ sky130_fd_sc_hd__a22o_1
Xfanout573 _06649_ vssd1 vssd1 vccd1 vccd1 net573 sky130_fd_sc_hd__buf_2
Xfanout584 net586 vssd1 vssd1 vccd1 vccd1 net584 sky130_fd_sc_hd__clkbuf_4
XANTENNA_clkbuf_leaf_13_clk_A clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09688__A2 _04655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout595 _06523_ vssd1 vssd1 vccd1 vccd1 net595 sky130_fd_sc_hd__buf_4
XANTENNA__12141__B1 net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1051 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11673__B _06644_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12921_ _07658_ net265 _07656_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[220\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15640_ ag2.body\[439\] net125 _01622_ ag2.body\[431\] vssd1 vssd1 vccd1 vccd1 _00905_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__14969__B1 net51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12852_ _06672_ _07538_ vssd1 vssd1 vccd1 vccd1 _07627_ sky130_fd_sc_hd__or2_1
XANTENNA__10289__B net1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11803_ net435 _06689_ _06719_ _06771_ _06774_ vssd1 vssd1 vccd1 vccd1 _06775_ sky130_fd_sc_hd__a32o_1
X_15571_ ag2.body\[489\] net135 _01615_ ag2.body\[481\] vssd1 vssd1 vccd1 vccd1 _00843_
+ sky130_fd_sc_hd__a22o_1
X_12783_ net286 _07593_ _07594_ net1823 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[146\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12444__A1 net1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_28_clk_A clknet_4_4__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12785__A net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12444__B2 net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11878__S0 net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_53_clk clknet_4_6__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_53_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_16_1344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17310_ ag2.body\[395\] net852 vssd1 vssd1 vccd1 vccd1 _02989_ sky130_fd_sc_hd__xor2_1
XFILLER_0_84_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14522_ _08676_ _08678_ _08679_ _08682_ vssd1 vssd1 vccd1 vccd1 _08683_ sky130_fd_sc_hd__or4_4
X_11734_ img_gen.tracker.frame\[26\] net618 net601 img_gen.tracker.frame\[29\] vssd1
+ vssd1 vccd1 vccd1 _06706_ sky130_fd_sc_hd__o22a_1
X_18290_ track.nextHighScore\[1\] net326 vssd1 vssd1 vccd1 vccd1 _03786_ sky130_fd_sc_hd__nor2_1
XFILLER_0_51_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17278__A1_N net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16900__A2_N net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17241_ ag2.body\[623\] net928 vssd1 vssd1 vccd1 vccd1 _02920_ sky130_fd_sc_hd__xnor2_1
X_14453_ net989 ag2.body\[433\] vssd1 vssd1 vccd1 vccd1 _08614_ sky130_fd_sc_hd__xor2_1
XANTENNA__20383__RESET_B net1374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11665_ net1147 _06636_ vssd1 vssd1 vccd1 vccd1 _06637_ sky130_fd_sc_hd__nand2_1
XANTENNA__16591__C1 net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20363__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10616_ ag2.body\[49\] net1198 vssd1 vssd1 vccd1 vccd1 _05589_ sky130_fd_sc_hd__xor2_1
XFILLER_0_36_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13404_ net284 net312 _07553_ _07873_ net1675 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[488\]
+ sky130_fd_sc_hd__a32o_1
X_17172_ _04161_ net882 net939 _04163_ _02850_ vssd1 vssd1 vccd1 vccd1 _02851_ sky130_fd_sc_hd__a221o_1
X_14384_ net1031 ag2.body\[301\] vssd1 vssd1 vccd1 vccd1 _08545_ sky130_fd_sc_hd__xor2_1
X_11596_ net505 _06567_ _06568_ vssd1 vssd1 vccd1 vccd1 _06569_ sky130_fd_sc_hd__or3_1
XFILLER_0_109_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11955__B1 net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16123_ net348 _01797_ _01801_ _01742_ vssd1 vssd1 vccd1 vccd1 _01802_ sky130_fd_sc_hd__o211a_1
XANTENNA__11688__X _06660_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13335_ net249 _07846_ _07847_ net1895 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[445\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__15146__B1 net50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10547_ ag2.body\[225\] net1206 vssd1 vssd1 vccd1 vccd1 _05520_ sky130_fd_sc_hd__nand2_1
XFILLER_0_84_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14064__X _08225_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16054_ net956 _01715_ vssd1 vssd1 vccd1 vccd1 _01733_ sky130_fd_sc_hd__nand2_1
X_13266_ net255 _07819_ _07820_ net1605 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[403\]
+ sky130_fd_sc_hd__a22o_1
X_10478_ net643 _04695_ _04572_ vssd1 vssd1 vccd1 vccd1 _05451_ sky130_fd_sc_hd__a21oi_2
XANTENNA__11707__B1 net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10752__B _05669_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12217_ img_gen.updater.commands.mode\[1\] _04391_ vssd1 vssd1 vccd1 vccd1 _07187_
+ sky130_fd_sc_hd__nor2_2
X_15005_ control.body\[994\] net152 _01552_ control.body\[986\] vssd1 vssd1 vccd1
+ vccd1 _00340_ sky130_fd_sc_hd__a22o_1
XANTENNA__17438__A2 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13197_ net675 _07788_ vssd1 vssd1 vccd1 vccd1 _07789_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_88_3003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_3014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19813_ clknet_leaf_124_clk _00757_ net1405 vssd1 vssd1 vccd1 vccd1 ag2.body\[579\]
+ sky130_fd_sc_hd__dfrtp_4
X_12148_ img_gen.tracker.frame\[444\] net614 net568 vssd1 vssd1 vccd1 vccd1 _07120_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_62_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10930__B2 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19744_ clknet_leaf_129_clk net2357 net1325 vssd1 vssd1 vccd1 vccd1 control.body\[654\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__15336__A _05283_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16956_ ag2.body\[294\] net700 net692 ag2.body\[295\] _02634_ vssd1 vssd1 vccd1 vccd1
+ _02635_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_10_Right_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12079_ net469 _07042_ _07045_ _06660_ vssd1 vssd1 vccd1 vccd1 _07051_ sky130_fd_sc_hd__a31o_1
XANTENNA__12132__B1 net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15907_ ag2.body\[197\] net132 _01651_ ag2.body\[189\] vssd1 vssd1 vccd1 vccd1 _01143_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11583__B net1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19675_ clknet_leaf_117_clk _00619_ net1384 vssd1 vssd1 vccd1 vccd1 control.body\[713\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11486__A2 _04469_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16887_ _02558_ _02563_ _02564_ _02565_ vssd1 vssd1 vccd1 vccd1 _02566_ sky130_fd_sc_hd__or4_1
XANTENNA__17071__B1 net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10694__B1 net1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_118 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18626_ clknet_leaf_0_clk img_gen.tracker.next_frame\[64\] net1243 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[64\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__17610__A2 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11891__C1 net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15838_ _05698_ net59 vssd1 vssd1 vccd1 vccd1 _01644_ sky130_fd_sc_hd__nor2_4
XANTENNA__18603__CLK clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10199__B net1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19729__CLK clknet_leaf_132_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_1325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1179 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18557_ clknet_leaf_43_clk _00083_ net1373 vssd1 vssd1 vccd1 vccd1 control.fsm.temp\[2\]
+ sky130_fd_sc_hd__dfstp_1
X_15769_ ag2.body\[313\] net209 _01637_ ag2.body\[305\] vssd1 vssd1 vccd1 vccd1 _01019_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_38_1591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_44_clk clknet_4_7__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_44_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_47_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18166__A3 _03705_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17508_ _03183_ _03186_ vssd1 vssd1 vccd1 vccd1 _03187_ sky130_fd_sc_hd__or2_1
XFILLER_0_74_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09290_ sound_gen.osc1.count\[2\] _04308_ vssd1 vssd1 vccd1 vccd1 _04310_ sky130_fd_sc_hd__or2_1
XANTENNA__16177__A2 net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18488_ net1516 net1510 vssd1 vssd1 vccd1 vccd1 _00019_ sky130_fd_sc_hd__or2_1
XFILLER_0_111_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10997__B2 ag2.body\[342\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17439_ _04041_ net856 net953 _04043_ vssd1 vssd1 vccd1 vccd1 _03118_ sky130_fd_sc_hd__o22a_1
XFILLER_0_118_949 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_14 _03446_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18753__CLK clknet_leaf_144_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13303__B _07483_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_25 net1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_36 _08924_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10646__C _05587_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20450_ clknet_leaf_41_clk _01337_ net1371 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[86\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__13935__B2 ag2.body\[70\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19109_ clknet_leaf_0_clk img_gen.tracker.next_frame\[547\] net1245 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[547\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15137__B1 net50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20381_ clknet_leaf_40_clk _01268_ net1374 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[17\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__17677__A2 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_1106 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout117_A net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19109__CLK clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16885__B1 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_676 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10007__X _04980_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1026_A net1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13973__B net60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout486_A net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14150__A net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12123__B1 net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09244__A net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11493__B net1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout653_A net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11108__A_N net1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_106_Right_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1395_A net1404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17601__A2 net733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09626_ net910 net905 net914 vssd1 vssd1 vccd1 vccd1 _04599_ sky130_fd_sc_hd__nand3_4
XFILLER_0_74_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12876__Y _07639_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17180__B net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09557_ net1072 control.body\[726\] vssd1 vssd1 vccd1 vccd1 _04530_ sky130_fd_sc_hd__xor2_1
XANTENNA__09898__B net1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout820_A net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1183_X net1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_35_clk clknet_4_5__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_35_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout539_X net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout918_A net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13053__X _07720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_825 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__20386__CLK clknet_leaf_43_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11634__C1 net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09488_ ag2.body\[372\] net1138 vssd1 vssd1 vccd1 vccd1 _04461_ sky130_fd_sc_hd__xor2_1
XANTENNA__16168__A2 net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_869 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14179__A1 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14179__B2 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15376__B1 _01594_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16573__C1 _02228_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout706_X net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18292__A track.nextHighScore\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13926__A1 ag2.body\[70\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11450_ net1161 control.body\[955\] vssd1 vssd1 vccd1 vccd1 _06423_ sky130_fd_sc_hd__xor2_1
XANTENNA__13926__B2 ag2.body\[62\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_338 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10401_ _05362_ _05363_ _05369_ _05370_ _05373_ vssd1 vssd1 vccd1 vccd1 _05374_ sky130_fd_sc_hd__a221o_1
XANTENNA__10204__A3 _05176_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16325__C1 net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11381_ net1220 control.body\[640\] vssd1 vssd1 vccd1 vccd1 _06354_ sky130_fd_sc_hd__nand2_1
XANTENNA__10853__A net1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20579_ clknet_leaf_107_clk _01436_ _00043_ vssd1 vssd1 vccd1 vccd1 sound_gen.osc1.count\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_13120_ net291 _07750_ _07751_ net1591 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[326\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_81_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10332_ _04600_ _05304_ vssd1 vssd1 vccd1 vccd1 _05305_ sky130_fd_sc_hd__nor2_1
XFILLER_0_132_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11668__B net1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10572__B net1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13051_ net268 _07718_ _07719_ net1711 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[289\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__17636__A ag2.body\[162\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10263_ _05211_ _05222_ _05223_ _05235_ vssd1 vssd1 vccd1 vccd1 _05236_ sky130_fd_sc_hd__a2bb2oi_1
XFILLER_0_63_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16540__A net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12002_ img_gen.tracker.frame\[433\] net613 net597 img_gen.tracker.frame\[436\] vssd1
+ vssd1 vccd1 vccd1 _06974_ sky130_fd_sc_hd__o22a_1
XANTENNA__13883__B net56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1302 net1310 vssd1 vssd1 vccd1 vccd1 net1302 sky130_fd_sc_hd__clkbuf_4
X_10194_ ag2.body\[119\] net1065 vssd1 vssd1 vccd1 vccd1 _05167_ sky130_fd_sc_hd__or2_1
Xfanout1313 net1314 vssd1 vssd1 vccd1 vccd1 net1313 sky130_fd_sc_hd__clkbuf_4
Xfanout1324 net1333 vssd1 vssd1 vccd1 vccd1 net1324 sky130_fd_sc_hd__clkbuf_4
X_16810_ _02487_ _02488_ vssd1 vssd1 vccd1 vccd1 _02489_ sky130_fd_sc_hd__nand2_1
Xfanout1335 net1337 vssd1 vssd1 vccd1 vccd1 net1335 sky130_fd_sc_hd__clkbuf_4
XANTENNA__14103__A1 net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1346 net1357 vssd1 vssd1 vccd1 vccd1 net1346 sky130_fd_sc_hd__clkbuf_4
XANTENNA__14103__B2 net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17790_ net1016 _03463_ vssd1 vssd1 vccd1 vccd1 _03466_ sky130_fd_sc_hd__and2_1
Xfanout1357 net1505 vssd1 vssd1 vccd1 vccd1 net1357 sky130_fd_sc_hd__buf_4
Xfanout370 _01908_ vssd1 vssd1 vccd1 vccd1 net370 sky130_fd_sc_hd__buf_2
XFILLER_0_17_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18626__CLK clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1368 net1369 vssd1 vssd1 vccd1 vccd1 net1368 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12499__B net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1379 net1383 vssd1 vssd1 vccd1 vccd1 net1379 sky130_fd_sc_hd__clkbuf_4
Xfanout381 _01706_ vssd1 vssd1 vccd1 vccd1 net381 sky130_fd_sc_hd__buf_2
Xfanout392 net393 vssd1 vssd1 vccd1 vccd1 net392 sky130_fd_sc_hd__buf_4
X_16741_ obsg2.obstacleArray\[36\] net490 net481 obsg2.obstacleArray\[37\] vssd1 vssd1
+ vccd1 vccd1 _02420_ sky130_fd_sc_hd__a22o_1
X_13953_ ag2.body\[94\] net191 _08155_ ag2.body\[86\] vssd1 vssd1 vccd1 vccd1 _00175_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_57_1422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11468__A2 _04599_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17053__B1 net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19460_ clknet_leaf_109_clk _00404_ net1417 vssd1 vssd1 vccd1 vccd1 control.body\[930\]
+ sky130_fd_sc_hd__dfrtp_1
X_12904_ net245 _07650_ _07651_ net1753 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[210\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_57_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16672_ obsg2.obstacleArray\[30\] obsg2.obstacleArray\[31\] net447 vssd1 vssd1 vccd1
+ vccd1 _02351_ sky130_fd_sc_hd__mux2_1
X_13884_ ag2.body\[32\] net115 _08148_ ag2.body\[24\] vssd1 vssd1 vccd1 vccd1 _00113_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__14406__A2 ag2.body\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18186__B net41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18411_ _03839_ _03899_ _03900_ vssd1 vssd1 vccd1 vccd1 _03901_ sky130_fd_sc_hd__a21o_1
XFILLER_0_134_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15623_ _06314_ net56 vssd1 vssd1 vccd1 vccd1 _01621_ sky130_fd_sc_hd__nor2_2
XANTENNA__17090__B net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12835_ _07431_ _07618_ vssd1 vssd1 vccd1 vccd1 _07619_ sky130_fd_sc_hd__nor2_1
X_19391_ clknet_leaf_102_clk _00335_ net1428 vssd1 vssd1 vccd1 vccd1 control.body\[1005\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__18776__CLK clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_26_clk clknet_4_4__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_26_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_130_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_1644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18342_ _04642_ _08026_ _03827_ vssd1 vssd1 vccd1 vccd1 _03838_ sky130_fd_sc_hd__and3_1
XANTENNA__11625__C1 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15554_ ag2.body\[507\] net186 _01612_ ag2.body\[499\] vssd1 vssd1 vccd1 vccd1 _00829_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_57_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12766_ net284 _07585_ _07586_ net1879 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[137\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__10747__B net1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14505_ net981 _04056_ ag2.body\[183\] net792 vssd1 vssd1 vccd1 vccd1 _08666_ sky130_fd_sc_hd__a22o_1
X_18273_ net516 _03775_ vssd1 vssd1 vccd1 vccd1 _01384_ sky130_fd_sc_hd__nor2_1
XANTENNA__15367__B1 _01593_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11717_ _06668_ net386 _06688_ vssd1 vssd1 vccd1 vccd1 _06689_ sky130_fd_sc_hd__or3_1
XANTENNA__15906__A2 net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12697_ net344 net329 _07433_ vssd1 vssd1 vccd1 vccd1 _07553_ sky130_fd_sc_hd__and3_2
X_15485_ ag2.body\[573\] net112 _01605_ ag2.body\[565\] vssd1 vssd1 vccd1 vccd1 _00767_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_51_1098 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17224_ _04104_ net876 net934 _04108_ vssd1 vssd1 vccd1 vccd1 _02903_ sky130_fd_sc_hd__o22a_1
XANTENNA__13917__A1 ag2.body\[62\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14436_ net987 ag2.body\[17\] vssd1 vssd1 vccd1 vccd1 _08597_ sky130_fd_sc_hd__xor2_1
X_11648_ _06465_ _06484_ _06620_ _06619_ vssd1 vssd1 vccd1 vccd1 _06621_ sky130_fd_sc_hd__a31o_1
XFILLER_0_25_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14590__A1 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17155_ ag2.body\[610\] net722 net928 _04221_ _02833_ vssd1 vssd1 vccd1 vccd1 _02834_
+ sky130_fd_sc_hd__a221o_1
X_11579_ _06550_ _06551_ net507 vssd1 vssd1 vccd1 vccd1 _06552_ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14590__B2 net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16316__C1 net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14367_ net817 ag2.body\[603\] ag2.body\[607\] net790 _08526_ vssd1 vssd1 vccd1 vccd1
+ _08528_ sky130_fd_sc_hd__a221o_1
XFILLER_0_3_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold807 control.body\[657\] vssd1 vssd1 vccd1 vccd1 net2369 sky130_fd_sc_hd__dlygate4sd3_1
X_16106_ net349 _01780_ _01784_ _01743_ vssd1 vssd1 vccd1 vccd1 _01785_ sky130_fd_sc_hd__o211a_1
XFILLER_0_12_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold818 control.body\[956\] vssd1 vssd1 vccd1 vccd1 net2380 sky130_fd_sc_hd__dlygate4sd3_1
X_13318_ _07494_ _07807_ net645 vssd1 vssd1 vccd1 vccd1 _07841_ sky130_fd_sc_hd__o21a_1
XFILLER_0_64_1448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14298_ ag2.body\[220\] net816 net984 _04069_ vssd1 vssd1 vccd1 vccd1 _08459_ sky130_fd_sc_hd__a2bb2o_1
X_17086_ ag2.body\[198\] net938 vssd1 vssd1 vccd1 vccd1 _02765_ sky130_fd_sc_hd__xnor2_1
Xhold829 control.body\[828\] vssd1 vssd1 vccd1 vccd1 net2391 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10482__B net1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19401__CLK clknet_leaf_102_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16037_ _01684_ _01687_ vssd1 vssd1 vccd1 vccd1 _01716_ sky130_fd_sc_hd__nand2_1
X_13249_ net227 _07811_ vssd1 vssd1 vccd1 vccd1 _07812_ sky130_fd_sc_hd__nor2_1
XANTENNA__16450__A net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14522__X _08683_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_111_3696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16619__B1 net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_877 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18084__A2 _03539_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17988_ _03540_ _03545_ _03553_ vssd1 vssd1 vccd1 vccd1 _03606_ sky130_fd_sc_hd__or3_1
XANTENNA__19551__CLK clknet_leaf_115_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19727_ clknet_leaf_132_clk _00671_ net1304 vssd1 vssd1 vccd1 vccd1 control.body\[669\]
+ sky130_fd_sc_hd__dfrtp_1
X_16939_ ag2.body\[525\] net951 vssd1 vssd1 vccd1 vccd1 _02618_ sky130_fd_sc_hd__xor2_1
XANTENNA__13853__B1 _08134_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09521__A1 net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19658_ clknet_leaf_119_clk _00602_ net1390 vssd1 vssd1 vccd1 vccd1 control.body\[728\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09999__A net1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10003__A net1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17595__A1 net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18096__B _03679_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09411_ img_gen.updater.commands.mode\[2\] img_gen.updater.commands.mode\[0\] vssd1
+ vssd1 vccd1 vccd1 _04391_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_36_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18609_ clknet_leaf_17_clk img_gen.tracker.next_frame\[47\] net1318 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[47\] sky130_fd_sc_hd__dfrtp_1
X_19589_ clknet_leaf_118_clk _00533_ net1386 vssd1 vssd1 vccd1 vccd1 control.body\[803\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09809__C1 _04739_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_460 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_17_clk clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_17_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_90_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09342_ sound_gen.osc1.stayCount\[7\] _04345_ vssd1 vssd1 vccd1 vccd1 _04346_ sky130_fd_sc_hd__and2_1
XANTENNA__13314__A net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_110 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10657__B net1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11092__B1 net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09273_ sound_gen.osc1.stayCount\[18\] sound_gen.osc1.stayCount\[16\] _04288_ vssd1
+ vssd1 vccd1 vccd1 _04296_ sky130_fd_sc_hd__o21a_1
XFILLER_0_5_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15358__B1 _01592_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11631__A2 net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout234_A net236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20502_ clknet_leaf_22_clk _01389_ net1359 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[138\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_99_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_1594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14581__A1 net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20433_ clknet_leaf_22_clk _01320_ net1358 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[69\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_71_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout401_A net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16307__C1 net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14581__B2 net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14145__A net996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1143_A ag2.x\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09239__A net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20364_ clknet_leaf_50_clk _01251_ net1370 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__11488__B net1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14333__A1 net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14333__B2 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20295_ clknet_leaf_36_clk control.divider.next_count\[16\] net1349 vssd1 vssd1 vccd1
+ vccd1 control.divider.count\[16\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout1310_A net1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1029_X net1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14799__B ag2.body\[294\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17175__B net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout391_X net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout770_A net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12895__A1 net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout489_X net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout868_A net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13048__X _07718_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08988_ ag2.body\[83\] vssd1 vssd1 vccd1 vccd1 _04013_ sky130_fd_sc_hd__inv_2
XFILLER_0_138_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13208__B _07639_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10950_ ag2.body\[173\] net1105 vssd1 vssd1 vccd1 vccd1 _05923_ sky130_fd_sc_hd__xor2_1
XANTENNA__19070__RESET_B net1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09702__A ag2.body\[70\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09609_ net1169 control.body\[634\] vssd1 vssd1 vccd1 vccd1 _04582_ sky130_fd_sc_hd__xor2_1
XANTENNA_fanout823_X net823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10881_ _05850_ _05851_ _05852_ _05853_ vssd1 vssd1 vccd1 vccd1 _05854_ sky130_fd_sc_hd__or4_1
XANTENNA__11870__A2 net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11607__C1 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12620_ net333 _07511_ vssd1 vssd1 vccd1 vccd1 _07512_ sky130_fd_sc_hd__nand2_1
XFILLER_0_136_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12551_ img_gen.tracker.frame\[35\] net652 _07473_ vssd1 vssd1 vccd1 vccd1 _07474_
+ sky130_fd_sc_hd__and3_1
XANTENNA__17889__A2 _03519_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14607__X _08768_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11502_ net1199 net1225 vssd1 vssd1 vccd1 vccd1 _06475_ sky130_fd_sc_hd__and2b_2
XFILLER_0_108_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_705 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15270_ control.body\[765\] net108 _01582_ net2381 vssd1 vssd1 vccd1 vccd1 _00575_
+ sky130_fd_sc_hd__a22o_1
X_12482_ net334 _07433_ vssd1 vssd1 vccd1 vccd1 _07434_ sky130_fd_sc_hd__nand2_1
XANTENNA__10854__Y _05827_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_134_4397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_850 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14221_ net982 ag2.body\[394\] vssd1 vssd1 vccd1 vccd1 _08382_ sky130_fd_sc_hd__xnor2_1
X_11433_ ag2.body\[398\] net1088 vssd1 vssd1 vccd1 vccd1 _06406_ sky130_fd_sc_hd__xor2_1
XANTENNA__14572__A1 net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19424__CLK clknet_leaf_111_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14572__B2 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14055__A net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14152_ net811 ag2.body\[596\] ag2.body\[597\] net806 _08312_ vssd1 vssd1 vccd1 vccd1
+ _08313_ sky130_fd_sc_hd__a221o_1
X_11364_ net783 control.body\[808\] _04243_ net1049 _06336_ vssd1 vssd1 vccd1 vccd1
+ _06337_ sky130_fd_sc_hd__a221o_1
XFILLER_0_46_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10315_ ag2.body\[614\] net1073 vssd1 vssd1 vccd1 vccd1 _05288_ sky130_fd_sc_hd__xor2_1
X_13103_ _07744_ net258 _07742_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[316\]
+ sky130_fd_sc_hd__mux2_1
X_18960_ clknet_leaf_7_clk img_gen.tracker.next_frame\[398\] net1266 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[398\] sky130_fd_sc_hd__dfrtp_1
X_14083_ net831 ag2.body\[562\] ag2.body\[566\] net799 vssd1 vssd1 vccd1 vccd1 _08244_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_123_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11295_ net1046 control.body\[687\] vssd1 vssd1 vccd1 vccd1 _06268_ sky130_fd_sc_hd__xor2_1
X_17911_ _03535_ _03544_ vssd1 vssd1 vccd1 vccd1 _03546_ sky130_fd_sc_hd__nor2_1
XANTENNA__19574__CLK clknet_leaf_118_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13034_ img_gen.tracker.frame\[280\] net649 vssd1 vssd1 vccd1 vccd1 _07712_ sky130_fd_sc_hd__and2_1
XANTENNA__14875__A2 net182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10246_ ag2.body\[323\] net1165 vssd1 vssd1 vccd1 vccd1 _05219_ sky130_fd_sc_hd__or2_1
XFILLER_0_119_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18891_ clknet_leaf_26_clk img_gen.tracker.next_frame\[329\] net1342 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[329\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_101_1622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1110 net1112 vssd1 vssd1 vccd1 vccd1 net1110 sky130_fd_sc_hd__clkbuf_4
XANTENNA__19840__RESET_B net1414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1121 net1122 vssd1 vssd1 vccd1 vccd1 net1121 sky130_fd_sc_hd__buf_4
X_17842_ img_gen.updater.commands.rR1.rainbowRNG\[3\] img_gen.updater.commands.rR1.rainbowRNG\[2\]
+ img_gen.updater.commands.rR1.rainbowRNG\[1\] img_gen.updater.commands.rR1.rainbowRNG\[0\]
+ vssd1 vssd1 vccd1 vccd1 _03498_ sky130_fd_sc_hd__and4_1
Xfanout1132 net1143 vssd1 vssd1 vccd1 vccd1 net1132 sky130_fd_sc_hd__buf_4
XANTENNA__10897__B1 _04573_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10177_ ag2.body\[421\] net1105 vssd1 vssd1 vccd1 vccd1 _05150_ sky130_fd_sc_hd__xor2_1
XFILLER_0_121_1070 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1143 ag2.x\[0\] vssd1 vssd1 vccd1 vccd1 net1143 sky130_fd_sc_hd__buf_4
Xfanout1154 net1155 vssd1 vssd1 vccd1 vccd1 net1154 sky130_fd_sc_hd__buf_4
XANTENNA__19158__RESET_B net1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20551__CLK clknet_leaf_105_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1165 net1166 vssd1 vssd1 vccd1 vccd1 net1165 sky130_fd_sc_hd__clkbuf_4
Xfanout1176 net1177 vssd1 vssd1 vccd1 vccd1 net1176 sky130_fd_sc_hd__buf_4
X_17773_ _03448_ _03449_ _03450_ _03451_ vssd1 vssd1 vccd1 vccd1 _03452_ sky130_fd_sc_hd__and4_1
XANTENNA__12099__C1 net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1187 net1188 vssd1 vssd1 vccd1 vccd1 net1187 sky130_fd_sc_hd__buf_4
X_14985_ control.body\[1008\] net151 _01549_ control.body\[1000\] vssd1 vssd1 vccd1
+ vccd1 _00322_ sky130_fd_sc_hd__a22o_1
XANTENNA__18197__A net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1198 net1199 vssd1 vssd1 vccd1 vccd1 net1198 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_135_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19512_ clknet_leaf_121_clk _00456_ net1402 vssd1 vssd1 vccd1 vccd1 control.body\[886\]
+ sky130_fd_sc_hd__dfrtp_1
X_16724_ _02397_ _02402_ net380 vssd1 vssd1 vccd1 vccd1 _02403_ sky130_fd_sc_hd__mux2_1
X_13936_ ag2.body\[79\] net185 _08153_ ag2.body\[71\] vssd1 vssd1 vccd1 vccd1 _00160_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_18_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19443_ clknet_leaf_109_clk _00387_ net1420 vssd1 vssd1 vccd1 vccd1 control.body\[945\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09612__A _04574_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16655_ obsg2.obstacleArray\[10\] obsg2.obstacleArray\[11\] net446 vssd1 vssd1 vccd1
+ vccd1 _02334_ sky130_fd_sc_hd__mux2_1
XFILLER_0_76_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10758__A net1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11861__A2 net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13867_ _04422_ _04519_ _04432_ vssd1 vssd1 vccd1 vccd1 _08141_ sky130_fd_sc_hd__a21bo_2
XFILLER_0_85_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13134__A net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15606_ _05885_ net63 vssd1 vssd1 vccd1 vccd1 _01620_ sky130_fd_sc_hd__and2_4
XFILLER_0_130_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12818_ net669 _07610_ vssd1 vssd1 vccd1 vccd1 _07611_ sky130_fd_sc_hd__nor2_1
XFILLER_0_9_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19374_ clknet_leaf_102_clk _00318_ net1426 vssd1 vssd1 vccd1 vccd1 control.body\[1020\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13063__A1 net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16586_ obsg2.obstacleArray\[65\] net451 net396 _02264_ vssd1 vssd1 vccd1 vccd1 _02265_
+ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_100_3364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_3375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13798_ _04275_ _08102_ _08096_ vssd1 vssd1 vccd1 vccd1 _00073_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_84_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11074__B1 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_100_3386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18325_ net906 _04641_ _03820_ _08036_ vssd1 vssd1 vccd1 vccd1 _03821_ sky130_fd_sc_hd__a31o_1
X_15537_ ag2.body\[523\] net160 _01611_ ag2.body\[515\] vssd1 vssd1 vccd1 vccd1 _00813_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_70_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12810__A1 net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12749_ net329 _07471_ vssd1 vssd1 vccd1 vccd1 _07578_ sky130_fd_sc_hd__nand2_2
XFILLER_0_44_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18256_ _03696_ net35 vssd1 vssd1 vccd1 vccd1 _03767_ sky130_fd_sc_hd__nor2_1
XFILLER_0_127_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15468_ ag2.body\[590\] net90 _01603_ ag2.body\[582\] vssd1 vssd1 vccd1 vccd1 _00752_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_4_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17207_ ag2.body\[54\] net937 vssd1 vssd1 vccd1 vccd1 _02886_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_117_3883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14419_ _08576_ _08577_ _08578_ _08579_ vssd1 vssd1 vccd1 vccd1 _08580_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_117_3894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18187_ obsg2.obstacleArray\[90\] _03732_ net531 vssd1 vssd1 vccd1 vccd1 _01341_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_4_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15399_ net2625 net82 _01581_ control.body\[632\] vssd1 vssd1 vccd1 vccd1 _00690_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_114_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_113_3758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17138_ ag2.body\[271\] net933 vssd1 vssd1 vccd1 vccd1 _02817_ sky130_fd_sc_hd__xor2_1
Xhold604 img_gen.updater.commands.rR1.rainbowRNG\[9\] vssd1 vssd1 vccd1 vccd1 net2166
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_128_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_113_3769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold615 img_gen.updater.commands.rR1.rainbowRNG\[4\] vssd1 vssd1 vccd1 vccd1 net2177
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold626 control.body\[653\] vssd1 vssd1 vccd1 vccd1 net2188 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__19928__RESET_B net1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold637 control.body\[1095\] vssd1 vssd1 vccd1 vccd1 net2199 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap356 _08050_ vssd1 vssd1 vccd1 vccd1 net356 sky130_fd_sc_hd__clkbuf_2
Xhold648 control.body\[654\] vssd1 vssd1 vccd1 vccd1 net2210 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09960_ ag2.body\[83\] net772 net1068 _04015_ _04932_ vssd1 vssd1 vccd1 vccd1 _04933_
+ sky130_fd_sc_hd__a221o_1
X_17069_ ag2.body\[29\] net946 vssd1 vssd1 vccd1 vccd1 _02748_ sky130_fd_sc_hd__xor2_1
Xhold659 control.body\[1069\] vssd1 vssd1 vccd1 vccd1 net2221 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14252__X _08413_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_6_clk clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_6_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_111_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20080_ clknet_leaf_77_clk _01024_ net1492 vssd1 vssd1 vccd1 vccd1 ag2.body\[318\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_106_1599 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09891_ ag2.body\[79\] net1065 vssd1 vssd1 vccd1 vccd1 _04864_ sky130_fd_sc_hd__xor2_1
XANTENNA__12877__A1 _07425_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16068__A1 net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10940__B net1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10352__A2 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14618__A2 ag2.body\[59\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout184_A net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09522__A net1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout351_A _01703_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1093_A ag2.x\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10767__B1_N _05517_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout449_A net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_931 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09325_ sound_gen.dac1.dacCount\[6\] sound_gen.dac1.dacCount\[5\] _04336_ vssd1 vssd1
+ vccd1 vccd1 _04337_ sky130_fd_sc_hd__and3_1
XFILLER_0_34_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_400 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1260_A net1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout616_A net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout237_X net237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09256_ ssdec1.in\[0\] vssd1 vssd1 vccd1 vccd1 _04281_ sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_4_10__f_clk_A clknet_3_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16074__B net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11499__A net1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09187_ ag2.body\[580\] vssd1 vssd1 vccd1 vccd1 _04212_ sky130_fd_sc_hd__inv_2
XFILLER_0_133_546 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20416_ clknet_leaf_35_clk _01303_ net1350 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[52\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_107_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19597__CLK clknet_leaf_118_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout985_A net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20347_ clknet_leaf_139_clk _01238_ net1292 vssd1 vssd1 vccd1 vccd1 img_gen.updater.commands.rR1.rainbowRNG\[7\]
+ sky130_fd_sc_hd__dfrtp_2
X_10100_ net911 net919 net922 vssd1 vssd1 vccd1 vccd1 _05073_ sky130_fd_sc_hd__or3_1
XANTENNA_fanout97_A net100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11946__B net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11080_ ag2.body\[540\] net1132 vssd1 vssd1 vccd1 vccd1 _06053_ sky130_fd_sc_hd__nand2_1
X_20278_ clknet_leaf_36_clk net1571 net1347 vssd1 vssd1 vccd1 vccd1 control.button1.Q\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_101_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12868__A1 net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout773_X net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10031_ _04184_ net1233 net1089 _04186_ vssd1 vssd1 vccd1 vccd1 _05004_ sky130_fd_sc_hd__a22o_1
XANTENNA__17256__B1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13219__A net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09416__B net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_127_4190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19251__RESET_B net1482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10343__A2 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout940_X net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17633__B net961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17008__B1 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_4076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_123_4087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15434__A _05287_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14770_ net1022 ag2.body\[102\] vssd1 vssd1 vccd1 vccd1 _08931_ sky130_fd_sc_hd__nand2_1
XANTENNA__12096__A2 net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11982_ img_gen.tracker.frame\[541\] net613 net596 img_gen.tracker.frame\[544\] _06953_
+ vssd1 vssd1 vccd1 vccd1 _06954_ sky130_fd_sc_hd__o221a_1
XANTENNA_fanout52_X net52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09432__A ag2.body\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13721_ net26 net25 vssd1 vssd1 vccd1 vccd1 toggle1.nextBlinkToggle\[0\] sky130_fd_sc_hd__nor2_1
XANTENNA__17920__Y _03554_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10933_ net769 control.body\[1035\] control.body\[1039\] net745 _05905_ vssd1 vssd1
+ vccd1 vccd1 _05906_ sky130_fd_sc_hd__o221a_1
XFILLER_0_93_1496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11843__A2 net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16231__A1 net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12496__C net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16440_ obsg2.obstacleArray\[92\] obsg2.obstacleArray\[93\] obsg2.obstacleArray\[94\]
+ obsg2.obstacleArray\[95\] net454 net398 vssd1 vssd1 vccd1 vccd1 _02119_ sky130_fd_sc_hd__mux4_1
X_13652_ control.divider.count\[18\] control.divider.count\[17\] _08005_ vssd1 vssd1
+ vccd1 vccd1 _08009_ sky130_fd_sc_hd__and3_1
XFILLER_0_85_238 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10864_ _05813_ _05819_ _05824_ _05836_ vssd1 vssd1 vccd1 vccd1 _05837_ sky130_fd_sc_hd__o31a_1
XFILLER_0_131_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18464__B net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12603_ net667 _07503_ vssd1 vssd1 vccd1 vccd1 _07504_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_136_4459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16371_ _01930_ _01947_ _01896_ vssd1 vssd1 vccd1 vccd1 _02050_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_137_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13583_ control.divider.count\[2\] control.divider.count\[3\] control.divider.count\[1\]
+ control.divider.count\[0\] vssd1 vssd1 vccd1 vccd1 _07958_ sky130_fd_sc_hd__and4_1
X_10795_ ag2.body\[38\] net1078 vssd1 vssd1 vccd1 vccd1 _05768_ sky130_fd_sc_hd__nand2_1
XANTENNA__14793__B2 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18110_ net353 _03624_ vssd1 vssd1 vccd1 vccd1 _03689_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_45_1687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15322_ control.body\[714\] net73 _01589_ net2350 vssd1 vssd1 vccd1 vccd1 _00620_
+ sky130_fd_sc_hd__a22o_1
X_19090_ clknet_leaf_146_clk img_gen.tracker.next_frame\[528\] net1240 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[528\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_45_1698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12534_ net313 _07464_ vssd1 vssd1 vccd1 vccd1 _07465_ sky130_fd_sc_hd__or2_1
XFILLER_0_124_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18041_ net42 _03643_ vssd1 vssd1 vccd1 vccd1 _03644_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_10_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15253_ net2372 net97 _01579_ control.body\[775\] vssd1 vssd1 vccd1 vccd1 _00561_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_10_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12465_ net290 _07419_ _07420_ net1746 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[2\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11359__A1 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11359__B2 net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14204_ net1009 ag2.body\[367\] vssd1 vssd1 vccd1 vccd1 _08365_ sky130_fd_sc_hd__xor2_1
XFILLER_0_112_719 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11416_ net1051 control.body\[855\] vssd1 vssd1 vccd1 vccd1 _06389_ sky130_fd_sc_hd__nand2_1
X_12396_ img_gen.updater.commands.rR1.rainbowRNG\[3\] net248 net241 _07337_ vssd1
+ vssd1 vccd1 vccd1 _07360_ sky130_fd_sc_hd__a211o_1
X_15184_ net2363 net101 _01572_ control.body\[825\] vssd1 vssd1 vccd1 vccd1 _00499_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_22_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12020__A2 net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16298__A1 net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11347_ ag2.body\[446\] net1079 vssd1 vssd1 vccd1 vccd1 _06320_ sky130_fd_sc_hd__xor2_1
X_14135_ net972 ag2.body\[171\] vssd1 vssd1 vccd1 vccd1 _08296_ sky130_fd_sc_hd__nand2_1
XANTENNA__18964__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19992_ clknet_leaf_65_clk _00936_ net1474 vssd1 vssd1 vccd1 vccd1 ag2.body\[406\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_91_3087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_1598 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16204__S net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_3098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11278_ _06242_ _06243_ _06245_ _06246_ vssd1 vssd1 vccd1 vccd1 _06251_ sky130_fd_sc_hd__a22o_1
X_14066_ net976 ag2.body\[211\] vssd1 vssd1 vccd1 vccd1 _08227_ sky130_fd_sc_hd__xor2_1
X_18943_ clknet_leaf_143_clk img_gen.tracker.next_frame\[381\] net1290 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[381\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__11856__B net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17247__B1 net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13017_ img_gen.tracker.frame\[271\] net657 vssd1 vssd1 vccd1 vccd1 _07704_ sky130_fd_sc_hd__and2_1
X_10229_ ag2.body\[560\] net1228 vssd1 vssd1 vccd1 vccd1 _05202_ sky130_fd_sc_hd__xor2_1
X_18874_ clknet_leaf_13_clk img_gen.tracker.next_frame\[312\] net1284 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[312\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__12033__A net1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17825_ _03962_ ag2.appleSet _01535_ vssd1 vssd1 vccd1 vccd1 _03489_ sky130_fd_sc_hd__a21bo_1
Xhold1 obsmode.sOBSMODE.sync vssd1 vssd1 vccd1 vccd1 net1563 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__17543__B net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_3551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_3562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17756_ _02481_ _03434_ vssd1 vssd1 vccd1 vccd1 _03435_ sky130_fd_sc_hd__nand2_1
XANTENNA__12087__A2 net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14968_ net2278 net152 net51 control.body\[1018\] vssd1 vssd1 vccd1 vccd1 _00308_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_102_3426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12687__B net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_3437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16707_ obsg2.obstacleArray\[72\] net490 net481 obsg2.obstacleArray\[73\] _02385_
+ vssd1 vssd1 vccd1 vccd1 _02386_ sky130_fd_sc_hd__a221o_1
X_13919_ _04669_ net61 vssd1 vssd1 vccd1 vccd1 _08152_ sky130_fd_sc_hd__nor2_2
X_17687_ ag2.body\[155\] net855 vssd1 vssd1 vccd1 vccd1 _03366_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_102_3448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11834__A2 net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14899_ net2275 net178 _01540_ control.body\[1084\] vssd1 vssd1 vccd1 vccd1 _00246_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_72_1558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19426_ clknet_leaf_111_clk _00370_ net1422 vssd1 vssd1 vccd1 vccd1 control.body\[960\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_134_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16638_ _02310_ _02312_ _02316_ _02228_ vssd1 vssd1 vccd1 vccd1 _02317_ sky130_fd_sc_hd__o211a_1
XFILLER_0_9_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13036__A1 net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_8_Right_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19357_ clknet_leaf_101_clk _00301_ net1438 vssd1 vssd1 vccd1 vccd1 control.body\[1035\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16569_ net395 _02247_ _02246_ net361 vssd1 vssd1 vccd1 vccd1 _02248_ sky130_fd_sc_hd__a211o_1
XFILLER_0_31_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_3945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16175__A _01728_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_119_3956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09110_ ag2.body\[379\] vssd1 vssd1 vccd1 vccd1 _04135_ sky130_fd_sc_hd__inv_2
XANTENNA__11598__A1 _06485_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_119_3967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18308_ _03799_ _03803_ _03797_ vssd1 vssd1 vccd1 vccd1 _03804_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_61_2190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19288_ clknet_leaf_98_clk net2394 net1446 vssd1 vssd1 vccd1 vccd1 control.body\[1110\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19259__Q ag2.body\[122\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09041_ ag2.body\[206\] vssd1 vssd1 vccd1 vccd1 _04066_ sky130_fd_sc_hd__inv_2
X_18239_ obsg2.obstacleArray\[116\] _03758_ net526 vssd1 vssd1 vccd1 vccd1 _01367_
+ sky130_fd_sc_hd__o21a_1
XANTENNA__14536__A1 net975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14536__B2 net1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18278__A2 net48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold401 img_gen.tracker.frame\[202\] vssd1 vssd1 vccd1 vccd1 net1963 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1020 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold412 img_gen.tracker.frame\[529\] vssd1 vssd1 vccd1 vccd1 net1974 sky130_fd_sc_hd__dlygate4sd3_1
X_20201_ clknet_leaf_54_clk _01145_ net1454 vssd1 vssd1 vccd1 vccd1 ag2.body\[199\]
+ sky130_fd_sc_hd__dfrtp_4
Xhold423 img_gen.tracker.frame\[205\] vssd1 vssd1 vccd1 vccd1 net1985 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__17486__B1 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold434 img_gen.tracker.frame\[155\] vssd1 vssd1 vccd1 vccd1 net1996 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10373__D net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold445 img_gen.tracker.frame\[64\] vssd1 vssd1 vccd1 vccd1 net2007 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_2573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold456 img_gen.tracker.frame\[468\] vssd1 vssd1 vccd1 vccd1 net2018 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold467 img_gen.tracker.frame\[314\] vssd1 vssd1 vccd1 vccd1 net2029 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20132_ clknet_leaf_80_clk _01076_ net1485 vssd1 vssd1 vccd1 vccd1 ag2.body\[258\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__09517__A net1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold478 img_gen.tracker.frame\[425\] vssd1 vssd1 vccd1 vccd1 net2040 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09943_ _04911_ _04912_ _04914_ _04915_ vssd1 vssd1 vccd1 vccd1 _04916_ sky130_fd_sc_hd__or4_2
Xhold489 img_gen.tracker.frame\[542\] vssd1 vssd1 vccd1 vccd1 net2051 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout903 control.body_update.curr_length\[5\] vssd1 vssd1 vccd1 vccd1 net903 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_70_2448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_39_Right_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout914 net915 vssd1 vssd1 vccd1 vccd1 net914 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_70_2459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout925 net926 vssd1 vssd1 vccd1 vccd1 net925 sky130_fd_sc_hd__clkbuf_4
Xfanout936 obsg2.randCord\[7\] vssd1 vssd1 vccd1 vccd1 net936 sky130_fd_sc_hd__buf_4
XANTENNA_fanout399_A net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20063_ clknet_leaf_73_clk _01007_ net1500 vssd1 vssd1 vccd1 vccd1 ag2.body\[333\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__17429__A2_N net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09874_ ag2.body\[167\] net1057 vssd1 vssd1 vccd1 vccd1 _04847_ sky130_fd_sc_hd__xor2_1
Xfanout947 net950 vssd1 vssd1 vccd1 vccd1 net947 sky130_fd_sc_hd__clkbuf_8
Xfanout958 net968 vssd1 vssd1 vccd1 vccd1 net958 sky130_fd_sc_hd__buf_4
Xfanout969 obsg2.obstacleFlag vssd1 vssd1 vccd1 vccd1 net969 sky130_fd_sc_hd__buf_2
Xhold1101 control.body\[946\] vssd1 vssd1 vccd1 vccd1 net2663 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1106_A ag2.x\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17453__B net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout187_X net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout566_A net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_2967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09479__B1 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_2978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13275__A1 net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_2989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10089__A1 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10089__B2 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_2388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11825__A2 net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_2399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout733_A _04263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout354_X net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10398__A net1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1475_A net1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1096_X net1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1470 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18837__CLK clknet_leaf_142_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16764__A2 net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_48_Right_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout521_X net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout900_A net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout619_X net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1263_X net1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09308_ sound_gen.osc1.count\[7\] _04327_ vssd1 vssd1 vccd1 vccd1 _04328_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_35_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10580_ ag2.body\[191\] net1057 vssd1 vssd1 vccd1 vccd1 _05553_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_131_4312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_1328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_131_4323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17909__A net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09239_ net860 vssd1 vssd1 vccd1 vccd1 _04264_ sky130_fd_sc_hd__inv_2
XFILLER_0_17_872 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18987__CLK clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_1551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_4_9__f_clk_A clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12250_ _07188_ _07214_ _07204_ vssd1 vssd1 vccd1 vccd1 _07220_ sky130_fd_sc_hd__o21a_1
XANTENNA__12002__A2 net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout988_X net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11201_ control.body\[878\] net1076 vssd1 vssd1 vccd1 vccd1 _06174_ sky130_fd_sc_hd__nand2b_1
XANTENNA__17477__B1 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09954__A1 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09954__B2 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12181_ net1197 ag2.apple_cord\[1\] vssd1 vssd1 vccd1 vccd1 _07153_ sky130_fd_sc_hd__or2_1
XANTENNA__10861__A net1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20621__1546 vssd1 vssd1 vccd1 vccd1 _20621__1546/HI net1546 sky130_fd_sc_hd__conb_1
XPHY_EDGE_ROW_57_Right_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11132_ _06103_ _06104_ net637 vssd1 vssd1 vccd1 vccd1 _06105_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_129_4252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_4263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10580__B net1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold990 control.body\[714\] vssd1 vssd1 vccd1 vccd1 net2552 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_38_1480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11063_ ag2.body\[435\] net1154 vssd1 vssd1 vccd1 vccd1 _06036_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_125_4127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15940_ ag2.body\[162\] net196 _01653_ ag2.body\[154\] vssd1 vssd1 vccd1 vccd1 _01172_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_25_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_1491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_34_1355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10014_ ag2.body\[265\] net1212 vssd1 vssd1 vccd1 vccd1 _04987_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_34_1366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15871_ ag2.body\[229\] net160 _01647_ net2290 vssd1 vssd1 vccd1 vccd1 _01111_ sky130_fd_sc_hd__a22o_1
XANTENNA__16452__A1 net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17610_ net703 net696 _01814_ _03288_ _03287_ vssd1 vssd1 vccd1 vccd1 _03289_ sky130_fd_sc_hd__a41o_1
X_14822_ net839 ag2.body\[153\] ag2.body\[158\] net802 vssd1 vssd1 vccd1 vccd1 _01493_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_95_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12069__A2 net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13266__A1 net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18590_ clknet_leaf_13_clk img_gen.tracker.next_frame\[28\] net1278 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[28\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_99_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17541_ _04111_ net966 net702 ag2.body\[326\] vssd1 vssd1 vccd1 vccd1 _03220_ sky130_fd_sc_hd__o22a_1
X_14753_ _08907_ _08911_ _08912_ _08913_ vssd1 vssd1 vccd1 vccd1 _08914_ sky130_fd_sc_hd__or4_1
X_11965_ img_gen.tracker.frame\[484\] net600 net584 img_gen.tracker.frame\[490\] _06936_
+ vssd1 vssd1 vccd1 vccd1 _06937_ sky130_fd_sc_hd__o221a_1
XPHY_EDGE_ROW_66_Right_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_1375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13704_ track.highScore\[4\] _08026_ vssd1 vssd1 vccd1 vccd1 _08045_ sky130_fd_sc_hd__nor2_1
XFILLER_0_135_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10916_ ag2.body\[462\] net1079 vssd1 vssd1 vccd1 vccd1 _05889_ sky130_fd_sc_hd__xnor2_1
XANTENNA__13018__A1 net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17472_ _03145_ _03147_ _03150_ vssd1 vssd1 vccd1 vccd1 _03151_ sky130_fd_sc_hd__or3_1
X_14684_ net844 ag2.body\[88\] _04021_ net1021 _08843_ vssd1 vssd1 vccd1 vccd1 _08845_
+ sky130_fd_sc_hd__o221a_1
XANTENNA__16755__A2 net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11896_ net1215 net1190 img_gen.tracker.frame\[61\] vssd1 vssd1 vccd1 vccd1 _06868_
+ sky130_fd_sc_hd__or3_1
XANTENNA__19762__CLK clknet_leaf_127_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19211_ clknet_leaf_85_clk _00155_ net1483 vssd1 vssd1 vccd1 vccd1 ag2.body\[74\]
+ sky130_fd_sc_hd__dfrtp_2
X_16423_ net363 _02090_ _02094_ _02101_ vssd1 vssd1 vccd1 vccd1 _02102_ sky130_fd_sc_hd__a31o_1
XFILLER_0_132_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13635_ control.divider.count\[12\] _07995_ net222 vssd1 vssd1 vccd1 vccd1 _07998_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_89_1318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10847_ ag2.body\[40\] net1219 vssd1 vssd1 vccd1 vccd1 _05820_ sky130_fd_sc_hd__nand2_1
XANTENNA__14508__A net1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19142_ clknet_leaf_138_clk net1583 net1292 vssd1 vssd1 vccd1 vccd1 img_gen.control.detect4.Q\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_16354_ obsg2.obstacleArray\[4\] obsg2.obstacleArray\[5\] net409 vssd1 vssd1 vccd1
+ vccd1 _02033_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_15_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13566_ _07944_ vssd1 vssd1 vccd1 vccd1 _07945_ sky130_fd_sc_hd__inv_2
XFILLER_0_109_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17825__B1_N _01535_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10778_ _05745_ _05750_ vssd1 vssd1 vccd1 vccd1 _05751_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_97_3274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14518__A1 net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_97_3285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15305_ control.body\[732\] net77 _01586_ net2412 vssd1 vssd1 vccd1 vccd1 _00606_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_109_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_3296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19073_ clknet_leaf_29_clk img_gen.tracker.next_frame\[511\] net1335 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[511\] sky130_fd_sc_hd__dfrtp_1
X_12517_ net1937 net650 _07455_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[19\]
+ sky130_fd_sc_hd__and3_1
X_16285_ obsg2.obstacleArray\[126\] obsg2.obstacleArray\[127\] net407 vssd1 vssd1
+ vccd1 vccd1 _01964_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_855 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14518__B2 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13497_ net230 _07910_ _07911_ net1607 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[543\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_67_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_3149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18024_ obsg2.obstacleArray\[27\] _03632_ net531 vssd1 vssd1 vccd1 vccd1 _01278_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_2_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15236_ _05223_ net63 vssd1 vssd1 vccd1 vccd1 _01578_ sky130_fd_sc_hd__and2_2
XFILLER_0_124_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12448_ _07282_ _07396_ _07408_ _07300_ vssd1 vssd1 vccd1 vccd1 net31 sky130_fd_sc_hd__a22o_1
XFILLER_0_1_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_75_Right_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17468__B1 net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09945__A1 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15167_ control.body\[850\] net102 _01570_ net2286 vssd1 vssd1 vccd1 vccd1 _00484_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_22_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09945__B2 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12379_ img_gen.updater.commands.count\[2\] _07190_ _07342_ img_gen.updater.commands.count\[12\]
+ vssd1 vssd1 vccd1 vccd1 _07344_ sky130_fd_sc_hd__or4bb_1
XANTENNA__14243__A net1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11752__A1 net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14118_ net979 ag2.body\[570\] vssd1 vssd1 vccd1 vccd1 _08279_ sky130_fd_sc_hd__xor2_1
X_19975_ clknet_leaf_62_clk _00919_ net1478 vssd1 vssd1 vccd1 vccd1 ag2.body\[421\]
+ sky130_fd_sc_hd__dfrtp_4
X_15098_ net2604 net148 _01563_ net2153 vssd1 vssd1 vccd1 vccd1 _00422_ sky130_fd_sc_hd__a22o_1
XANTENNA__10490__B net1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_3602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14049_ net819 ag2.body\[187\] ag2.body\[188\] net811 vssd1 vssd1 vccd1 vccd1 _08210_
+ sky130_fd_sc_hd__a22o_1
X_18926_ clknet_leaf_139_clk img_gen.tracker.next_frame\[364\] net1290 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[364\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_43_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_3613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_3624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09624__X _04597_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17273__B net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19292__CLK clknet_leaf_98_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18857_ clknet_leaf_18_clk img_gen.tracker.next_frame\[295\] net1319 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[295\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_136_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17808_ _03474_ _03476_ _03970_ vssd1 vssd1 vccd1 vccd1 _01219_ sky130_fd_sc_hd__mux2_1
X_09590_ net1058 control.body\[911\] vssd1 vssd1 vccd1 vccd1 _04563_ sky130_fd_sc_hd__xor2_1
XFILLER_0_94_1057 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13257__A1 net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18788_ clknet_leaf_12_clk img_gen.tracker.next_frame\[226\] net1285 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[226\] sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_84_Right_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_19_Left_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_1188 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_1079 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17739_ _02844_ _02849_ _03414_ _03415_ _03417_ vssd1 vssd1 vccd1 vccd1 _03418_ sky130_fd_sc_hd__o2111a_1
XTAP_TAPCELL_ROW_82_2820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_2831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_2230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_2241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12480__A2 _07425_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_2252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09800__A net1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19409_ clknet_leaf_103_clk _00353_ net1428 vssd1 vssd1 vccd1 vccd1 control.body\[991\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14757__A1 net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16210__A4 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14757__B2 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10946__A _05909_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11541__S net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout147_A net154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09633__B1 _04605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12209__Y _07181_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14509__A1 net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11440__B1 _04772_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14509__B2 net1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15706__B1 _01629_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout314_A net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_28_Left_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09024_ ag2.body\[160\] vssd1 vssd1 vccd1 vccd1 _04049_ sky130_fd_sc_hd__inv_2
XFILLER_0_116_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1056_A net1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_93_Right_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_76_2635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_76_2646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16352__B net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_57_2056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17459__B1 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold220 img_gen.tracker.frame\[375\] vssd1 vssd1 vccd1 vccd1 net1782 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_2067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold231 img_gen.tracker.frame\[122\] vssd1 vssd1 vccd1 vccd1 net1793 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1223_A net1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold242 img_gen.tracker.frame\[72\] vssd1 vssd1 vccd1 vccd1 net1804 sky130_fd_sc_hd__dlygate4sd3_1
Xhold253 img_gen.tracker.frame\[273\] vssd1 vssd1 vccd1 vccd1 net1815 sky130_fd_sc_hd__dlygate4sd3_1
Xhold264 img_gen.tracker.frame\[172\] vssd1 vssd1 vccd1 vccd1 net1826 sky130_fd_sc_hd__dlygate4sd3_1
Xhold275 img_gen.tracker.frame\[66\] vssd1 vssd1 vccd1 vccd1 net1837 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16779__S net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout700 net702 vssd1 vssd1 vccd1 vccd1 net700 sky130_fd_sc_hd__buf_4
XANTENNA_fanout683_A net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold286 img_gen.tracker.frame\[531\] vssd1 vssd1 vccd1 vccd1 net1848 sky130_fd_sc_hd__dlygate4sd3_1
Xhold297 img_gen.tracker.frame\[386\] vssd1 vssd1 vccd1 vccd1 net1859 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20115_ clknet_leaf_80_clk _01059_ net1488 vssd1 vssd1 vccd1 vccd1 ag2.body\[273\]
+ sky130_fd_sc_hd__dfrtp_4
Xfanout711 net712 vssd1 vssd1 vccd1 vccd1 net711 sky130_fd_sc_hd__clkbuf_4
X_09926_ _04107_ net1091 net747 ag2.body\[319\] _04898_ vssd1 vssd1 vccd1 vccd1 _04899_
+ sky130_fd_sc_hd__a221o_1
Xfanout722 net723 vssd1 vssd1 vccd1 vccd1 net722 sky130_fd_sc_hd__clkbuf_4
Xfanout733 _04263_ vssd1 vssd1 vccd1 vccd1 net733 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout1011_X net1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout744 _04234_ vssd1 vssd1 vccd1 vccd1 net744 sky130_fd_sc_hd__buf_4
XANTENNA_fanout1109_X net1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout755 net756 vssd1 vssd1 vccd1 vccd1 net755 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_77_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20046_ clknet_leaf_68_clk _00990_ net1498 vssd1 vssd1 vccd1 vccd1 ag2.body\[348\]
+ sky130_fd_sc_hd__dfrtp_4
Xfanout766 _04231_ vssd1 vssd1 vccd1 vccd1 net766 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout850_A net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09857_ _04824_ _04825_ _04826_ _04829_ vssd1 vssd1 vccd1 vccd1 _04830_ sky130_fd_sc_hd__or4_2
Xfanout777 net778 vssd1 vssd1 vccd1 vccd1 net777 sky130_fd_sc_hd__buf_4
XANTENNA__17183__B net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout788 net789 vssd1 vssd1 vccd1 vccd1 net788 sky130_fd_sc_hd__buf_4
XANTENNA_fanout471_X net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout948_A net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout799 net805 vssd1 vssd1 vccd1 vccd1 net799 sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_37_Left_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_1244 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09788_ _04754_ _04755_ _04760_ vssd1 vssd1 vccd1 vccd1 _04761_ sky130_fd_sc_hd__a21o_1
XANTENNA__16985__A2 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_1299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout736_X net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1478_X net1478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15712__A _06041_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_856 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_4510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11750_ net1046 _06721_ vssd1 vssd1 vccd1 vccd1 _06722_ sky130_fd_sc_hd__and2_1
XANTENNA__16737__A2 net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10701_ ag2.body\[20\] net1128 vssd1 vssd1 vccd1 vccd1 _05674_ sky130_fd_sc_hd__or2_1
XANTENNA__10856__A net1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11681_ img_gen.tracker.frame\[134\] net619 net601 img_gen.tracker.frame\[137\] vssd1
+ vssd1 vccd1 vccd1 _06653_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_42_1602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11304__X _06277_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_1613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13420_ _07564_ net303 vssd1 vssd1 vccd1 vccd1 _07880_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_23_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10632_ _05601_ _05602_ _05603_ _05604_ vssd1 vssd1 vccd1 vccd1 _05605_ sky130_fd_sc_hd__a22o_1
XANTENNA__10575__B net1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_46_Left_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17639__A ag2.body\[163\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13351_ net274 _07852_ _07853_ net2054 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[455\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_36_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10563_ net1059 ag2.body\[519\] vssd1 vssd1 vccd1 vccd1 _05536_ sky130_fd_sc_hd__and2b_1
XFILLER_0_134_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19165__CLK clknet_leaf_52_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19613__RESET_B net1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_959 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12302_ _07218_ _07221_ vssd1 vssd1 vccd1 vccd1 _07269_ sky130_fd_sc_hd__and2b_1
X_16070_ obsg2.obstacleArray\[120\] obsg2.obstacleArray\[121\] net424 vssd1 vssd1
+ vccd1 vccd1 _01749_ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15173__A1 _06180_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10494_ ag2.body\[548\] net762 net1101 _04202_ vssd1 vssd1 vccd1 vccd1 _05467_ sky130_fd_sc_hd__a22o_1
X_13282_ net280 _07825_ _07826_ net1615 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[413\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12790__B net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09927__A1 _04418_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11687__A net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15021_ _05476_ net66 vssd1 vssd1 vccd1 vccd1 _01555_ sky130_fd_sc_hd__and2_2
XFILLER_0_133_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12233_ img_gen.updater.commands.cmd_num\[1\] _04273_ img_gen.updater.commands.cmd_num\[3\]
+ img_gen.updater.commands.cmd_num\[4\] vssd1 vssd1 vccd1 vccd1 _07203_ sky130_fd_sc_hd__or4_1
XFILLER_0_60_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10591__A net1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11195__C1 net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12164_ img_gen.tracker.frame\[399\] net600 net545 img_gen.tracker.frame\[402\] _07135_
+ vssd1 vssd1 vccd1 vccd1 _07136_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_36_1428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11115_ net1062 control.body\[1103\] vssd1 vssd1 vccd1 vccd1 _06088_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_120_1124 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16972_ ag2.body\[411\] net718 net691 ag2.body\[415\] _02646_ vssd1 vssd1 vccd1 vccd1
+ _02651_ sky130_fd_sc_hd__a221o_1
XFILLER_0_100_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_9_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12095_ img_gen.tracker.frame\[348\] net627 net609 img_gen.tracker.frame\[351\] _07066_
+ vssd1 vssd1 vccd1 vccd1 _07067_ sky130_fd_sc_hd__a221o_1
X_19760_ clknet_leaf_130_clk _00704_ net1316 vssd1 vssd1 vccd1 vccd1 control.body\[638\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_55_Left_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11046_ ag2.body\[385\] net1209 vssd1 vssd1 vccd1 vccd1 _06019_ sky130_fd_sc_hd__xnor2_1
X_15923_ ag2.body\[178\] net124 _01654_ ag2.body\[170\] vssd1 vssd1 vccd1 vccd1 _01156_
+ sky130_fd_sc_hd__a22o_1
X_18711_ clknet_leaf_144_clk img_gen.tracker.next_frame\[149\] net1255 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[149\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_127_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17093__B net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19691_ clknet_leaf_136_clk _00635_ net1302 vssd1 vssd1 vccd1 vccd1 control.body\[697\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__20292__CLK clknet_leaf_37_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15606__B net63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16425__A1 _02057_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11593__S0 net1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17622__B1 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18642_ clknet_leaf_131_clk img_gen.tracker.next_frame\[80\] net1314 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[80\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__13239__A1 net238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15854_ ag2.body\[246\] net174 _01645_ ag2.body\[238\] vssd1 vssd1 vccd1 vccd1 _01096_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_56_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14805_ net844 ag2.body\[288\] ag2.body\[290\] net830 _01475_ vssd1 vssd1 vccd1 vccd1
+ _01476_ sky130_fd_sc_hd__o221a_1
X_18573_ clknet_leaf_15_clk img_gen.tracker.next_frame\[11\] net1312 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[11\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15785_ _05909_ net60 vssd1 vssd1 vccd1 vccd1 _01639_ sky130_fd_sc_hd__nor2_2
XANTENNA__10102__Y _05075_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12997_ net337 net332 _07515_ vssd1 vssd1 vccd1 vccd1 _07694_ sky130_fd_sc_hd__and3_1
X_17524_ _04174_ net862 net962 _04176_ _03202_ vssd1 vssd1 vccd1 vccd1 _03203_ sky130_fd_sc_hd__a221o_1
XFILLER_0_118_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14736_ net1041 _04116_ ag2.body\[335\] net796 _08896_ vssd1 vssd1 vccd1 vccd1 _08897_
+ sky130_fd_sc_hd__a221o_1
X_11948_ img_gen.tracker.frame\[124\] net602 net561 _06919_ vssd1 vssd1 vccd1 vccd1
+ _06920_ sky130_fd_sc_hd__o211a_1
XANTENNA__16728__A2 net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17455_ _03130_ _03131_ _03132_ _03133_ vssd1 vssd1 vccd1 vccd1 _03134_ sky130_fd_sc_hd__nand4_1
XTAP_TAPCELL_ROW_99_3336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11670__B1 net1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_3347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14667_ _08821_ _08822_ _08825_ _08827_ vssd1 vssd1 vccd1 vccd1 _08828_ sky130_fd_sc_hd__a211o_1
XFILLER_0_131_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11879_ img_gen.tracker.frame\[4\] net606 net551 img_gen.tracker.frame\[7\] net566
+ vssd1 vssd1 vccd1 vccd1 _06851_ sky130_fd_sc_hd__o221a_1
X_16406_ net354 _02055_ vssd1 vssd1 vccd1 vccd1 _02085_ sky130_fd_sc_hd__or2_1
X_13618_ control.divider.count\[6\] _07985_ vssd1 vssd1 vccd1 vccd1 _07987_ sky130_fd_sc_hd__and2_1
X_17386_ ag2.body\[493\] net953 vssd1 vssd1 vccd1 vccd1 _03065_ sky130_fd_sc_hd__xor2_1
XANTENNA__19508__CLK clknet_leaf_113_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12214__A2 _07181_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14598_ net816 ag2.body\[308\] ag2.body\[310\] net803 _08756_ vssd1 vssd1 vccd1 vccd1
+ _08759_ sky130_fd_sc_hd__a221o_1
XFILLER_0_32_1383 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19125_ clknet_leaf_141_clk img_gen.tracker.next_frame\[563\] net1294 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[563\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_55_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16337_ net419 _02015_ _02014_ net372 vssd1 vssd1 vccd1 vccd1 _02016_ sky130_fd_sc_hd__a211o_1
XFILLER_0_67_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13549_ ssdec1.in\[1\] _04281_ vssd1 vssd1 vccd1 vccd1 _07931_ sky130_fd_sc_hd__or2_1
XANTENNA__12981__A net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17153__A2 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11973__A1 net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19056_ clknet_leaf_8_clk img_gen.tracker.next_frame\[494\] net1273 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[494\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16268_ _01918_ _01938_ _01946_ _01927_ _01916_ vssd1 vssd1 vccd1 vccd1 _01947_ sky130_fd_sc_hd__o32a_1
XFILLER_0_113_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18007_ net38 _03619_ obsg2.obstacleArray\[23\] vssd1 vssd1 vccd1 vccd1 _03620_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_2_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15219_ control.body\[800\] net95 _01576_ net2543 vssd1 vssd1 vccd1 vccd1 _00530_
+ sky130_fd_sc_hd__a22o_1
X_16199_ net348 _01877_ _01874_ _01742_ vssd1 vssd1 vccd1 vccd1 _01878_ sky130_fd_sc_hd__o211a_1
X_19958_ clknet_leaf_45_clk _00902_ net1382 vssd1 vssd1 vccd1 vccd1 ag2.body\[436\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__13478__A1 net250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18099__B _03681_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09711_ ag2.body\[245\] net1111 vssd1 vssd1 vccd1 vccd1 _04684_ sky130_fd_sc_hd__xor2_1
X_18909_ clknet_leaf_144_clk img_gen.tracker.next_frame\[347\] net1251 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[347\] sky130_fd_sc_hd__dfrtp_1
X_19889_ clknet_leaf_83_clk _00833_ net1480 vssd1 vssd1 vccd1 vccd1 ag2.body\[511\]
+ sky130_fd_sc_hd__dfrtp_4
X_09642_ net1084 control.body\[1022\] vssd1 vssd1 vccd1 vccd1 _04615_ sky130_fd_sc_hd__xor2_1
XFILLER_0_78_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_65_2303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_2314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17731__B _01818_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09573_ _04062_ net1233 net781 ag2.body\[201\] vssd1 vssd1 vccd1 vccd1 _04546_ sky130_fd_sc_hd__a22o_1
XFILLER_0_117_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout264_A net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_856 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16719__A2 net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20620__1545 vssd1 vssd1 vccd1 vccd1 _20620__1545/HI net1545 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_19_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12875__B net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout431_A _01734_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1173_A net1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14148__A net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout529_A net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12205__A2 _06825_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13402__A1 net238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_2708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13953__A2 net191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_59_2118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20595_ net1527 vssd1 vssd1 vccd1 vccd1 gpio_oeb[7] sky130_fd_sc_hd__buf_2
XFILLER_0_89_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12891__A _07443_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17144__A2 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_2129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1059_X net1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11037__A_N net1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17178__B net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16082__B net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout898_A net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09007_ ag2.body\[127\] vssd1 vssd1 vccd1 vccd1 _04032_ sky130_fd_sc_hd__inv_2
XFILLER_0_42_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17893__S obsg2.obstacleCount\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10519__A2 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1226_X net1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11716__A1 net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11300__A net1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_176 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout686_X net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1506 net1508 vssd1 vssd1 vccd1 vccd1 net1506 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_44_1298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_6_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13469__A1 net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1517 net1 vssd1 vssd1 vccd1 vccd1 net1517 sky130_fd_sc_hd__clkbuf_2
Xfanout530 net534 vssd1 vssd1 vccd1 vccd1 net530 sky130_fd_sc_hd__buf_2
XFILLER_0_22_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout541 net543 vssd1 vssd1 vccd1 vccd1 net541 sky130_fd_sc_hd__clkbuf_4
X_09909_ _04878_ _04879_ _04880_ _04881_ _04877_ vssd1 vssd1 vccd1 vccd1 _04882_ sky130_fd_sc_hd__a221o_1
XFILLER_0_121_1488 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout552 net553 vssd1 vssd1 vccd1 vccd1 net552 sky130_fd_sc_hd__clkbuf_4
Xfanout563 net567 vssd1 vssd1 vccd1 vccd1 net563 sky130_fd_sc_hd__buf_2
XANTENNA_fanout853_X net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout574 net575 vssd1 vssd1 vccd1 vccd1 net574 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_96_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09688__A3 _04660_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout585 net586 vssd1 vssd1 vccd1 vccd1 net585 sky130_fd_sc_hd__clkbuf_4
XANTENNA__17604__B1 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20029_ clknet_leaf_67_clk _00973_ net1473 vssd1 vssd1 vccd1 vccd1 ag2.body\[363\]
+ sky130_fd_sc_hd__dfrtp_4
Xfanout596 net598 vssd1 vssd1 vccd1 vccd1 net596 sky130_fd_sc_hd__clkbuf_4
X_12920_ img_gen.tracker.frame\[220\] net660 vssd1 vssd1 vccd1 vccd1 _07658_ sky130_fd_sc_hd__and2_1
XANTENNA__10203__X _05176_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10152__B1 net1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14418__B1 ag2.body\[534\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12851_ net287 _07625_ _07626_ net1790 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[182\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_38_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_48_1800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15630__A2 net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_17_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11802_ net387 _06772_ _06773_ net438 vssd1 vssd1 vccd1 vccd1 _06774_ sky130_fd_sc_hd__o31a_1
X_15570_ ag2.body\[488\] net135 _01615_ ag2.body\[480\] vssd1 vssd1 vccd1 vccd1 _00842_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_90_1241 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12782_ net261 _07593_ _07594_ net1695 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[145\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__09845__B1 _04817_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11878__S1 net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14521_ _08675_ _08681_ _08677_ _08680_ vssd1 vssd1 vccd1 vccd1 _08682_ sky130_fd_sc_hd__or4b_1
X_11733_ net474 _06703_ _06704_ _06696_ _06691_ vssd1 vssd1 vccd1 vccd1 _06705_ sky130_fd_sc_hd__o221a_1
XANTENNA__15918__B1 _01652_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14058__A net996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17240_ ag2.body\[617\] net730 net710 ag2.body\[620\] vssd1 vssd1 vccd1 vccd1 _02919_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_132_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14452_ _08603_ _08612_ _08606_ _08611_ vssd1 vssd1 vccd1 vccd1 _08613_ sky130_fd_sc_hd__or4b_1
XFILLER_0_33_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11664_ net1119 net1097 vssd1 vssd1 vccd1 vccd1 _06636_ sky130_fd_sc_hd__xor2_4
XFILLER_0_138_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_94_3200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10207__A1 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18555__CLK clknet_leaf_43_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13403_ net259 net312 _07553_ _07873_ net1919 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[487\]
+ sky130_fd_sc_hd__a32o_1
X_17171_ ag2.body\[458\] net860 vssd1 vssd1 vccd1 vccd1 _02850_ sky130_fd_sc_hd__xor2_1
XANTENNA__10207__B2 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10615_ net634 _04758_ vssd1 vssd1 vccd1 vccd1 _05588_ sky130_fd_sc_hd__nor2_1
XFILLER_0_135_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14383_ net816 ag2.body\[300\] ag2.body\[302\] net804 _08543_ vssd1 vssd1 vccd1 vccd1
+ _08544_ sky130_fd_sc_hd__a221o_1
XFILLER_0_107_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11595_ obsg2.obstacleArray\[11\] net633 net509 obsg2.obstacleArray\[15\] net1123
+ vssd1 vssd1 vccd1 vccd1 _06568_ sky130_fd_sc_hd__o221a_1
XFILLER_0_25_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19800__CLK clknet_leaf_127_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11955__A1 net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16122_ net376 _01800_ _01799_ net346 vssd1 vssd1 vccd1 vccd1 _01801_ sky130_fd_sc_hd__a211o_1
X_13334_ net228 _07846_ _07847_ net1802 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[444\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__15146__A1 _04421_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10546_ ag2.body\[228\] net1136 vssd1 vssd1 vccd1 vccd1 _05519_ sky130_fd_sc_hd__or2_1
XFILLER_0_121_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16053_ _01720_ _01730_ vssd1 vssd1 vccd1 vccd1 _01732_ sky130_fd_sc_hd__nand2b_2
X_13265_ net234 _07819_ _07820_ net1842 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[402\]
+ sky130_fd_sc_hd__a22o_1
X_10477_ net904 _04446_ net896 vssd1 vssd1 vccd1 vccd1 _05450_ sky130_fd_sc_hd__o21ai_1
XANTENNA__11210__A net1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15004_ control.body\[993\] net153 _01552_ control.body\[985\] vssd1 vssd1 vccd1
+ vccd1 _00339_ sky130_fd_sc_hd__a22o_1
XANTENNA__10752__C _05696_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12216_ img_gen.control.current\[1\] img_gen.control.current\[0\] _07185_ _07186_
+ vssd1 vssd1 vccd1 vccd1 img_gen.control.next\[1\] sky130_fd_sc_hd__o22a_1
X_13196_ net383 _07618_ vssd1 vssd1 vccd1 vccd1 _07788_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_63_Left_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13836__S net1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16646__B2 net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_3004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19812_ clknet_leaf_125_clk _00756_ net1410 vssd1 vssd1 vccd1 vccd1 ag2.body\[578\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_88_3015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12147_ _07099_ _07105_ _07111_ _07118_ net472 net437 vssd1 vssd1 vccd1 vccd1 _07119_
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_40_1641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_1517 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_1439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09615__A net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19743_ clknet_leaf_129_clk _00687_ net1325 vssd1 vssd1 vccd1 vccd1 control.body\[653\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__15336__B net52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16955_ ag2.body\[289\] net875 vssd1 vssd1 vccd1 vccd1 _02634_ sky130_fd_sc_hd__xor2_1
X_12078_ _07047_ _07049_ net572 vssd1 vssd1 vccd1 vccd1 _07050_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13137__A net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15906_ ag2.body\[196\] net132 _01651_ ag2.body\[188\] vssd1 vssd1 vccd1 vccd1 _01142_
+ sky130_fd_sc_hd__a22o_1
X_11029_ net1061 control.body\[1047\] vssd1 vssd1 vccd1 vccd1 _06002_ sky130_fd_sc_hd__nand2_1
X_16886_ _02557_ _02559_ _02560_ _02561_ vssd1 vssd1 vccd1 vccd1 _02565_ sky130_fd_sc_hd__or4_1
XFILLER_0_2_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19674_ clknet_leaf_136_clk _00618_ net1384 vssd1 vssd1 vccd1 vccd1 control.body\[712\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__15623__Y _01621_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18625_ clknet_leaf_0_clk img_gen.tracker.next_frame\[63\] net1248 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[63\] sky130_fd_sc_hd__dfrtp_1
X_15837_ ag2.body\[263\] net175 net49 ag2.body\[255\] vssd1 vssd1 vccd1 vccd1 _01081_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_56_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14458__A1_N net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_1570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18556_ clknet_leaf_43_clk _00082_ net1372 vssd1 vssd1 vccd1 vccd1 control.fsm.temp\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_133_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15768_ ag2.body\[312\] net209 _01637_ ag2.body\[304\] vssd1 vssd1 vccd1 vccd1 _01018_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_133_1359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16167__B net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_72_Left_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18020__B1 net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14719_ net846 ag2.body\[336\] ag2.body\[337\] net839 _08872_ vssd1 vssd1 vccd1 vccd1
+ _08880_ sky130_fd_sc_hd__a221o_1
XFILLER_0_75_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17507_ _03178_ _03179_ _03181_ _03185_ vssd1 vssd1 vccd1 vccd1 _03186_ sky130_fd_sc_hd__or4_1
X_18487_ net1514 net1508 vssd1 vssd1 vccd1 vccd1 _00018_ sky130_fd_sc_hd__or2_1
X_15699_ ag2.body\[380\] net140 _01628_ ag2.body\[372\] vssd1 vssd1 vccd1 vccd1 _00958_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_131_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10997__A2 net1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17438_ ag2.body\[144\] net741 net701 ag2.body\[150\] vssd1 vssd1 vccd1 vccd1 _03117_
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_129_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_15 _03446_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_26 _03442_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_37 _08924_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10646__D _05618_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17369_ ag2.body\[3\] _03047_ vssd1 vssd1 vccd1 vccd1 _03048_ sky130_fd_sc_hd__and2_1
XFILLER_0_127_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19108_ clknet_leaf_0_clk img_gen.tracker.next_frame\[546\] net1239 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[546\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_127_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20380_ clknet_leaf_40_clk _01267_ net1374 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[16\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_28_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19039_ clknet_leaf_6_clk img_gen.tracker.next_frame\[477\] net1267 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[477\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_63_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13699__A1 net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_81_Left_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11120__A net1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16637__A1 net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17834__A0 net1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_174 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14431__A net1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1019_A ag2.randCord\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09525__A net1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_105_clk_X clknet_leaf_105_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14976__A_N _04607_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10023__X _04996_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16496__S0 net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09625_ _04587_ _04597_ _04536_ _04570_ _04585_ vssd1 vssd1 vccd1 vccd1 _04598_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_39_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12886__A _07439_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout646_A net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15612__A2 net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1608 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15262__A _04416_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09556_ _04526_ _04527_ _04528_ vssd1 vssd1 vccd1 vccd1 _04529_ sky130_fd_sc_hd__a21o_1
XFILLER_0_66_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18578__CLK clknet_leaf_15_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11634__B1 net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_837 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout813_A _03969_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_906 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09487_ ag2.body\[369\] net1208 vssd1 vssd1 vccd1 vccd1 _04460_ sky130_fd_sc_hd__xor2_1
XANTENNA_fanout434_X net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1176_X net1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_1608 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11014__B net1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout601_X net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14606__A net994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17117__A2 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10400_ _05360_ _05361_ _05371_ _05372_ vssd1 vssd1 vccd1 vccd1 _05373_ sky130_fd_sc_hd__or4_1
XFILLER_0_117_994 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11380_ ag2.body\[474\] net774 _06352_ vssd1 vssd1 vccd1 vccd1 _06353_ sky130_fd_sc_hd__o21ai_1
X_20578_ clknet_leaf_107_clk _01435_ _00042_ vssd1 vssd1 vccd1 vccd1 sound_gen.osc1.count\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_10331_ net899 _04979_ net636 vssd1 vssd1 vccd1 vccd1 _05304_ sky130_fd_sc_hd__a21o_1
XANTENNA__16380__X _02059_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11030__A net1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10262_ _05231_ _05232_ _05234_ vssd1 vssd1 vccd1 vccd1 _05235_ sky130_fd_sc_hd__and3_1
X_13050_ net246 _07718_ _07719_ net1865 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[288\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__17636__B net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout970_X net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12001_ img_gen.tracker.frame\[451\] net540 _06972_ net568 vssd1 vssd1 vccd1 vccd1
+ _06973_ sky130_fd_sc_hd__o211a_1
XANTENNA__16628__B2 net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10193_ ag2.body\[119\] net1065 vssd1 vssd1 vccd1 vccd1 _05166_ sky130_fd_sc_hd__nand2_1
Xfanout1303 net1306 vssd1 vssd1 vccd1 vccd1 net1303 sky130_fd_sc_hd__clkbuf_4
XANTENNA__14341__A net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1314 net1324 vssd1 vssd1 vccd1 vccd1 net1314 sky130_fd_sc_hd__clkbuf_2
Xfanout1325 net1327 vssd1 vssd1 vccd1 vccd1 net1325 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10912__A2 _04980_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1336 net1337 vssd1 vssd1 vccd1 vccd1 net1336 sky130_fd_sc_hd__clkbuf_4
Xfanout1347 net1348 vssd1 vssd1 vccd1 vccd1 net1347 sky130_fd_sc_hd__clkbuf_4
Xfanout360 _02223_ vssd1 vssd1 vccd1 vccd1 net360 sky130_fd_sc_hd__clkbuf_4
Xfanout1358 net1359 vssd1 vssd1 vccd1 vccd1 net1358 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_108_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout371 _01907_ vssd1 vssd1 vccd1 vccd1 net371 sky130_fd_sc_hd__buf_4
Xfanout1369 net1370 vssd1 vssd1 vccd1 vccd1 net1369 sky130_fd_sc_hd__buf_2
X_16740_ _02416_ _02418_ net495 vssd1 vssd1 vccd1 vccd1 _02419_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout382 _06822_ vssd1 vssd1 vccd1 vccd1 net382 sky130_fd_sc_hd__buf_4
Xfanout393 _02217_ vssd1 vssd1 vccd1 vccd1 net393 sky130_fd_sc_hd__buf_2
X_13952_ ag2.body\[93\] net190 _08155_ ag2.body\[85\] vssd1 vssd1 vccd1 vccd1 _00174_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_57_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12665__A2 _07536_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11468__A3 _04982_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09722__X _04695_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12903_ net680 _07650_ vssd1 vssd1 vccd1 vccd1 _07651_ sky130_fd_sc_hd__nor2_1
X_16671_ obsg2.obstacleArray\[28\] obsg2.obstacleArray\[29\] net447 vssd1 vssd1 vccd1
+ vccd1 _02350_ sky130_fd_sc_hd__mux2_1
XANTENNA__11873__B1 net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15443__Y _01601_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13883_ _05670_ net56 vssd1 vssd1 vccd1 vccd1 _08148_ sky130_fd_sc_hd__nor2_2
X_15622_ ag2.body\[455\] net124 _01613_ ag2.body\[447\] vssd1 vssd1 vccd1 vccd1 _00889_
+ sky130_fd_sc_hd__a22o_1
X_18410_ _03839_ _03890_ vssd1 vssd1 vccd1 vccd1 _03900_ sky130_fd_sc_hd__nor2_1
XFILLER_0_97_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12834_ _06671_ _07526_ vssd1 vssd1 vccd1 vccd1 _07618_ sky130_fd_sc_hd__nand2_1
X_19390_ clknet_leaf_102_clk _00334_ net1426 vssd1 vssd1 vccd1 vccd1 control.body\[1004\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_33_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18341_ _03826_ _03836_ _03825_ vssd1 vssd1 vccd1 vccd1 _03837_ sky130_fd_sc_hd__a21o_1
XANTENNA__11625__B1 net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15553_ ag2.body\[506\] net186 _01612_ ag2.body\[498\] vssd1 vssd1 vccd1 vccd1 _00828_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_5_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12765_ net256 _07585_ _07586_ net1600 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[136\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_90_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14504_ net999 ag2.body\[176\] vssd1 vssd1 vccd1 vccd1 _08665_ sky130_fd_sc_hd__xor2_1
X_18272_ net319 _03567_ obsg2.obstacleArray\[133\] vssd1 vssd1 vccd1 vccd1 _03775_
+ sky130_fd_sc_hd__a21oi_1
X_11716_ net473 _06681_ _06687_ _06660_ vssd1 vssd1 vccd1 vccd1 _06688_ sky130_fd_sc_hd__o211a_1
XFILLER_0_70_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15484_ ag2.body\[572\] net111 _01605_ ag2.body\[564\] vssd1 vssd1 vccd1 vccd1 _00766_
+ sky130_fd_sc_hd__a22o_1
X_12696_ net283 net310 _07551_ _07552_ net1593 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[101\]
+ sky130_fd_sc_hd__a32o_1
X_17223_ _02898_ _02900_ _02901_ _02899_ vssd1 vssd1 vccd1 vccd1 _02902_ sky130_fd_sc_hd__or4b_1
X_14435_ net980 ag2.body\[18\] vssd1 vssd1 vccd1 vccd1 _08596_ sky130_fd_sc_hd__xor2_1
X_11647_ obsg2.obstacleArray\[136\] obsg2.obstacleArray\[137\] obsg2.obstacleArray\[138\]
+ obsg2.obstacleArray\[139\] net1124 net507 vssd1 vssd1 vccd1 vccd1 _06620_ sky130_fd_sc_hd__mux4_1
XANTENNA__17108__A2 net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18305__A1 track.nextHighScore\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14516__A net1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13420__A _07564_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17154_ net698 ag2.body\[614\] _04220_ net848 vssd1 vssd1 vccd1 vccd1 _02833_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__12050__B1 net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14366_ net1034 ag2.body\[604\] vssd1 vssd1 vccd1 vccd1 _08527_ sky130_fd_sc_hd__xnor2_1
X_11578_ obsg2.obstacleArray\[83\] obsg2.obstacleArray\[87\] net514 vssd1 vssd1 vccd1
+ vccd1 _06551_ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16105_ net378 _01783_ _01782_ net347 vssd1 vssd1 vccd1 vccd1 _01784_ sky130_fd_sc_hd__a211o_1
XFILLER_0_3_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13317_ net275 _07839_ _07840_ net1943 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[434\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_29_1547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold808 control.body\[879\] vssd1 vssd1 vccd1 vccd1 net2370 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17085_ ag2.body\[192\] net738 net849 _04061_ vssd1 vssd1 vccd1 vccd1 _02764_ sky130_fd_sc_hd__o22a_1
X_10529_ net1107 control.body\[917\] vssd1 vssd1 vccd1 vccd1 _05502_ sky130_fd_sc_hd__nand2_1
Xhold819 control.body\[757\] vssd1 vssd1 vccd1 vccd1 net2381 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14297_ net976 ag2.body\[219\] vssd1 vssd1 vccd1 vccd1 _08458_ sky130_fd_sc_hd__xor2_1
XFILLER_0_29_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16036_ net870 net860 net850 net882 vssd1 vssd1 vccd1 vccd1 _01715_ sky130_fd_sc_hd__nor4b_1
XFILLER_0_21_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13248_ net2053 net648 _07811_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[394\]
+ sky130_fd_sc_hd__and3_1
XANTENNA__17546__B net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_111_3697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18084__A3 net38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13179_ net277 _07778_ _07779_ net1833 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[356\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11561__C1 net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16095__A2 net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17987_ obsg2.obstacleArray\[17\] _03605_ net531 vssd1 vssd1 vccd1 vccd1 _01268_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_97_1247 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12105__A1 net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11539__S0 net1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19726_ clknet_leaf_129_clk net2397 net1329 vssd1 vssd1 vccd1 vccd1 control.body\[668\]
+ sky130_fd_sc_hd__dfrtp_1
X_16938_ ag2.body\[520\] net740 net711 ag2.body\[524\] _02616_ vssd1 vssd1 vccd1 vccd1
+ _02617_ sky130_fd_sc_hd__o221ai_1
XFILLER_0_79_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14397__A1_N net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_74_clk_A clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18241__B1 net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10667__A1 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09521__A2 _04493_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10667__B2 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19657_ clknet_leaf_133_clk _00601_ net1308 vssd1 vssd1 vccd1 vccd1 control.body\[743\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11864__B1 net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16869_ ag2.body\[464\] net880 vssd1 vssd1 vccd1 vccd1 _02548_ sky130_fd_sc_hd__xor2_1
XANTENNA__18720__CLK clknet_leaf_142_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09410_ img_gen.updater.commands.mode\[2\] img_gen.updater.commands.mode\[0\] vssd1
+ vssd1 vccd1 vccd1 _04390_ sky130_fd_sc_hd__and2b_1
X_18608_ clknet_leaf_17_clk img_gen.tracker.next_frame\[46\] net1319 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[46\] sky130_fd_sc_hd__dfrtp_1
X_19588_ clknet_leaf_118_clk _00532_ net1386 vssd1 vssd1 vccd1 vccd1 control.body\[802\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09809__B1 _04781_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10938__B net1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14802__B1 ag2.body\[295\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09341_ sound_gen.osc1.stayCount\[6\] sound_gen.osc1.stayCount\[5\] _04344_ vssd1
+ vssd1 vccd1 vccd1 _04345_ sky130_fd_sc_hd__and3_1
X_18539_ clknet_leaf_136_clk _00065_ net1301 vssd1 vssd1 vccd1 vccd1 img_gen.updater.commands.count\[8\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_90_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11115__A net1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_89_clk_A clknet_4_9__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11092__A1 _06041_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11092__B2 _05303_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09272_ sound_gen.osc1.stayCount\[15\] net535 _04292_ _04293_ _04294_ vssd1 vssd1
+ vccd1 vccd1 _04295_ sky130_fd_sc_hd__o221a_1
XFILLER_0_114_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16555__B1 net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_132_clk_A clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20501_ clknet_leaf_23_clk _01388_ net1362 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[137\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_1_1538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13908__A2 net90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16117__S net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14426__A net980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_1641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20432_ clknet_leaf_23_clk _01319_ net1359 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[68\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_126_780 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_12_clk_A clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10673__B net1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19226__CLK clknet_leaf_75_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12592__A1 net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20363_ clknet_leaf_21_clk _00003_ net1361 vssd1 vssd1 vccd1 vccd1 obsg2.obsNeeded\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_101_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1136_A net1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20294_ clknet_leaf_37_clk control.divider.next_count\[15\] net1349 vssd1 vssd1 vccd1
+ vccd1 control.divider.count\[15\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout596_A net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_27_clk_A clknet_4_4__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19376__CLK clknet_leaf_93_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08987_ ag2.body\[81\] vssd1 vssd1 vccd1 vccd1 _04012_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout763_A net765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout384_X net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15263__Y _01581_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11855__B1 net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17191__B net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout930_A net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout551_X net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1293_X net1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13505__A net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09608_ net1219 control.body\[632\] vssd1 vssd1 vccd1 vccd1 _04581_ sky130_fd_sc_hd__xor2_1
XFILLER_0_97_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09702__B net1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10880_ ag2.body\[528\] net1231 vssd1 vssd1 vccd1 vccd1 _05853_ sky130_fd_sc_hd__xor2_1
XANTENNA_fanout42_A net43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10848__B net1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11607__B1 net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09539_ _04507_ _04510_ _04511_ _04509_ vssd1 vssd1 vccd1 vccd1 _04512_ sky130_fd_sc_hd__or4b_2
XFILLER_0_17_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout816_X net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12550_ net2105 net649 _07473_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[34\]
+ sky130_fd_sc_hd__and3_1
XANTENNA__16546__B1 net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11501_ net1225 net1197 vssd1 vssd1 vccd1 vccd1 _06474_ sky130_fd_sc_hd__or2_1
XFILLER_0_81_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12481_ net469 net561 net556 _07312_ vssd1 vssd1 vccd1 vccd1 _07433_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_134_4398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14220_ net1028 ag2.body\[397\] vssd1 vssd1 vccd1 vccd1 _08381_ sky130_fd_sc_hd__xnor2_1
X_11432_ ag2.body\[392\] net1234 vssd1 vssd1 vccd1 vccd1 _06405_ sky130_fd_sc_hd__xor2_1
XFILLER_0_80_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11679__B net1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_430 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12583__A1 net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16849__B2 net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14151_ net806 ag2.body\[597\] ag2.body\[594\] net824 vssd1 vssd1 vccd1 vccd1 _08312_
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_132_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11363_ net1119 control.body\[812\] vssd1 vssd1 vccd1 vccd1 _06336_ sky130_fd_sc_hd__xor2_1
XFILLER_0_21_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13102_ img_gen.tracker.frame\[316\] net652 vssd1 vssd1 vccd1 vccd1 _07744_ sky130_fd_sc_hd__and2_1
X_10314_ _04421_ _04571_ net643 vssd1 vssd1 vccd1 vccd1 _05287_ sky130_fd_sc_hd__o21ai_2
X_14082_ net841 ag2.body\[560\] _04208_ net1035 _08237_ vssd1 vssd1 vccd1 vccd1 _08243_
+ sky130_fd_sc_hd__o221a_1
X_11294_ net742 _04859_ _06266_ _06253_ _06240_ vssd1 vssd1 vccd1 vccd1 _06267_ sky130_fd_sc_hd__o32a_2
XFILLER_0_120_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17910_ _03535_ _03544_ vssd1 vssd1 vccd1 vccd1 _03545_ sky130_fd_sc_hd__or2_2
XFILLER_0_24_1433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13033_ net238 _07710_ _07711_ net1737 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[279\]
+ sky130_fd_sc_hd__a22o_1
X_10245_ ag2.body\[323\] net1165 vssd1 vssd1 vccd1 vccd1 _05218_ sky130_fd_sc_hd__nand2_1
X_18890_ clknet_leaf_26_clk img_gen.tracker.next_frame\[328\] net1342 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[328\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__11543__C1 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1100 net1101 vssd1 vssd1 vccd1 vccd1 net1100 sky130_fd_sc_hd__buf_2
XFILLER_0_28_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1111 net1112 vssd1 vssd1 vccd1 vccd1 net1111 sky130_fd_sc_hd__clkbuf_4
X_10176_ ag2.body\[418\] net1178 vssd1 vssd1 vccd1 vccd1 _05149_ sky130_fd_sc_hd__xor2_1
Xfanout1122 ag2.x\[0\] vssd1 vssd1 vccd1 vccd1 net1122 sky130_fd_sc_hd__buf_2
X_17841_ ag2.apple_cord\[7\] net224 _03497_ net686 vssd1 vssd1 vccd1 vccd1 _01230_
+ sky130_fd_sc_hd__a211o_1
Xfanout1133 net1134 vssd1 vssd1 vccd1 vccd1 net1133 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_121_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1144 net1156 vssd1 vssd1 vccd1 vccd1 net1144 sky130_fd_sc_hd__buf_4
XFILLER_0_121_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1155 net1156 vssd1 vssd1 vccd1 vccd1 net1155 sky130_fd_sc_hd__clkbuf_4
Xfanout1166 ag2.y\[3\] vssd1 vssd1 vccd1 vccd1 net1166 sky130_fd_sc_hd__buf_4
X_17772_ _03124_ _03129_ _02556_ _02622_ vssd1 vssd1 vccd1 vccd1 _03451_ sky130_fd_sc_hd__o211a_1
Xfanout1177 net1178 vssd1 vssd1 vccd1 vccd1 net1177 sky130_fd_sc_hd__buf_4
XANTENNA__10104__A net1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14984_ net2120 net158 _01550_ net2203 vssd1 vssd1 vccd1 vccd1 _00321_ sky130_fd_sc_hd__a22o_1
Xfanout190 net191 vssd1 vssd1 vccd1 vccd1 net190 sky130_fd_sc_hd__clkbuf_2
Xfanout1188 net1189 vssd1 vssd1 vccd1 vccd1 net1188 sky130_fd_sc_hd__buf_4
Xfanout1199 net1200 vssd1 vssd1 vccd1 vccd1 net1199 sky130_fd_sc_hd__buf_4
X_19511_ clknet_leaf_121_clk _00455_ net1402 vssd1 vssd1 vccd1 vccd1 control.body\[885\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_135_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09503__A2 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16723_ _02399_ _02401_ net499 vssd1 vssd1 vccd1 vccd1 _02402_ sky130_fd_sc_hd__mux2_1
X_13935_ ag2.body\[78\] net185 _08153_ ag2.body\[70\] vssd1 vssd1 vccd1 vccd1 _00159_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11846__B1 net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19198__RESET_B net1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkload5_A clknet_4_11__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13415__A _07561_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16654_ net362 _02328_ _02332_ net358 vssd1 vssd1 vccd1 vccd1 _02333_ sky130_fd_sc_hd__o211a_1
X_19442_ clknet_leaf_109_clk _00386_ net1420 vssd1 vssd1 vccd1 vccd1 control.body\[944\]
+ sky130_fd_sc_hd__dfrtp_1
X_13866_ _08031_ _08035_ vssd1 vssd1 vccd1 vccd1 _08140_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_104_3490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15605_ ag2.body\[471\] net121 _01619_ ag2.body\[463\] vssd1 vssd1 vccd1 vccd1 _00873_
+ sky130_fd_sc_hd__a22o_1
X_12817_ net341 net327 net308 _07515_ vssd1 vssd1 vccd1 vccd1 _07610_ sky130_fd_sc_hd__and4_1
X_16585_ obsg2.obstacleArray\[64\] net446 vssd1 vssd1 vccd1 vccd1 _02264_ sky130_fd_sc_hd__or2_1
X_19373_ clknet_leaf_102_clk _00317_ net1436 vssd1 vssd1 vccd1 vccd1 control.body\[1019\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14260__A1 net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13797_ _08098_ _08101_ _08102_ vssd1 vssd1 vccd1 vccd1 _00072_ sky130_fd_sc_hd__and3_1
XFILLER_0_130_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14260__B2 net1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_100_3365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_100_3376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_100_3387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18324_ _04236_ _08028_ vssd1 vssd1 vccd1 vccd1 _03820_ sky130_fd_sc_hd__nor2_1
X_15536_ ag2.body\[522\] net160 _01611_ ag2.body\[514\] vssd1 vssd1 vccd1 vccd1 _00812_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_84_453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12748_ net284 _07576_ _07577_ net1775 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[128\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_45_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19249__CLK clknet_leaf_75_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16445__B net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18255_ net526 _03766_ vssd1 vssd1 vccd1 vccd1 _01375_ sky130_fd_sc_hd__and2_1
X_15467_ ag2.body\[589\] net89 _01603_ ag2.body\[581\] vssd1 vssd1 vccd1 vccd1 _00751_
+ sky130_fd_sc_hd__a22o_1
X_12679_ net289 _07543_ _07544_ net1796 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[92\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_114_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17206_ ag2.body\[54\] net937 vssd1 vssd1 vccd1 vccd1 _02885_ sky130_fd_sc_hd__nand2_1
XFILLER_0_114_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14418_ net991 _04193_ ag2.body\[534\] net804 vssd1 vssd1 vccd1 vccd1 _08579_ sky130_fd_sc_hd__a22o_1
X_18186_ _03628_ net41 vssd1 vssd1 vccd1 vccd1 _03732_ sky130_fd_sc_hd__nor2_1
XFILLER_0_114_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12023__B1 net557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11589__B _06561_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_117_3884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15398_ net2624 net80 _01596_ net2259 vssd1 vssd1 vccd1 vccd1 _00689_ sky130_fd_sc_hd__a22o_1
XANTENNA__20226__CLK clknet_leaf_66_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_117_3895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10493__B net1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11377__A2 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_884 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17137_ ag2.body\[267\] net854 vssd1 vssd1 vccd1 vccd1 _02816_ sky130_fd_sc_hd__xor2_1
X_14349_ net1018 ag2.body\[406\] vssd1 vssd1 vccd1 vccd1 _08510_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_113_3759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold605 control.body\[1053\] vssd1 vssd1 vccd1 vccd1 net2167 sky130_fd_sc_hd__dlygate4sd3_1
Xhold616 control.body\[1089\] vssd1 vssd1 vccd1 vccd1 net2178 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold627 obsg2.arraySet vssd1 vssd1 vccd1 vccd1 net2189 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__19399__CLK clknet_leaf_102_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09627__X _04600_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold638 _00241_ vssd1 vssd1 vccd1 vccd1 net2200 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xmax_cap357 _02228_ vssd1 vssd1 vccd1 vccd1 net357 sky130_fd_sc_hd__buf_4
X_17068_ _02743_ _02744_ _02745_ _02746_ vssd1 vssd1 vccd1 vccd1 _02747_ sky130_fd_sc_hd__a22o_1
Xhold649 control.body\[664\] vssd1 vssd1 vccd1 vccd1 net2211 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17276__B net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xmax_cap368 _01911_ vssd1 vssd1 vccd1 vccd1 net368 sky130_fd_sc_hd__buf_4
X_16019_ _01695_ _01697_ vssd1 vssd1 vccd1 vccd1 _01698_ sky130_fd_sc_hd__nand2_2
XFILLER_0_100_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09890_ net894 _04861_ vssd1 vssd1 vccd1 vccd1 _04863_ sky130_fd_sc_hd__nor2_2
XANTENNA__12877__A2 _07638_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13309__B net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1006 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16400__S net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09803__A net1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19709_ clknet_leaf_134_clk _00653_ net1307 vssd1 vssd1 vccd1 vccd1 control.body\[683\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_75_1331 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11837__B1 net550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15524__B net65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15028__B1 _01555_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16225__C1 net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12586__D _07312_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20455__RESET_B net1356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1086_A net1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09324_ sound_gen.dac1.dacCount\[4\] sound_gen.dac1.dacCount\[3\] _04335_ vssd1 vssd1
+ vccd1 vccd1 _04336_ sky130_fd_sc_hd__and3_1
XFILLER_0_90_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09255_ img_gen.updater.commands.rR1.rainbowRNG\[0\] vssd1 vssd1 vccd1 vccd1 _04280_
+ sky130_fd_sc_hd__inv_2
XANTENNA_fanout511_A net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout132_X net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14156__A net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout609_A net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13060__A net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18616__CLK clknet_leaf_144_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11499__B net1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09186_ ag2.body\[579\] vssd1 vssd1 vccd1 vccd1 _04211_ sky130_fd_sc_hd__inv_2
XFILLER_0_133_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_575 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12565__A1 net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20415_ clknet_leaf_39_clk _01302_ net1352 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[51\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA_fanout1041_X net1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1139_X net1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20346_ clknet_leaf_139_clk _01237_ net1292 vssd1 vssd1 vccd1 vccd1 img_gen.updater.commands.rR1.rainbowRNG\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__17186__B net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16700__B1 net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout880_A net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16090__B net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18766__CLK clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout978_A ag2.randCord\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13059__X _07723_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout599_X net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20277_ clknet_leaf_36_clk net2 net1347 vssd1 vssd1 vccd1 vccd1 control.button1.Q\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_102_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10328__B1 _05287_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10030_ ag2.body\[507\] net771 net756 ag2.body\[509\] vssd1 vssd1 vccd1 vccd1 _05003_
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_60_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout766_X net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_4191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18205__B1 net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15434__B net52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_4088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout933_X net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11981_ img_gen.tracker.frame\[550\] net579 vssd1 vssd1 vccd1 vccd1 _06953_ sky130_fd_sc_hd__or2_1
XANTENNA__10859__A net1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15019__B1 _01553_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17559__A2 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13720_ _08053_ vssd1 vssd1 vccd1 vccd1 track.nextHighScore\[7\] sky130_fd_sc_hd__inv_2
XFILLER_0_58_1584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17930__A net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09432__B net1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10932_ net775 control.body\[1034\] control.body\[1038\] net750 vssd1 vssd1 vccd1
+ vccd1 _05905_ sky130_fd_sc_hd__o22a_1
XANTENNA_fanout45_X net45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_1459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13651_ _08007_ _08008_ vssd1 vssd1 vccd1 vccd1 control.divider.next_count\[17\]
+ sky130_fd_sc_hd__nor2_1
XANTENNA__15721__Y _01631_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12496__D net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10863_ _05827_ _05831_ _05835_ vssd1 vssd1 vccd1 vccd1 _05836_ sky130_fd_sc_hd__or3_1
XANTENNA__17154__A1_N net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12602_ _07431_ _07502_ vssd1 vssd1 vccd1 vccd1 _07503_ sky130_fd_sc_hd__nor2_1
XFILLER_0_112_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16370_ _01918_ _01955_ _01963_ _02048_ _01929_ vssd1 vssd1 vccd1 vccd1 _02049_ sky130_fd_sc_hd__o311a_1
X_13582_ control.divider.count\[2\] control.divider.count\[1\] control.divider.count\[0\]
+ vssd1 vssd1 vccd1 vccd1 _07957_ sky130_fd_sc_hd__nand3_1
XANTENNA__16519__B1 _02057_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10794_ ag2.body\[36\] net1128 vssd1 vssd1 vccd1 vccd1 _05767_ sky130_fd_sc_hd__or2_1
XFILLER_0_81_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15321_ control.body\[713\] net73 _01589_ net2343 vssd1 vssd1 vccd1 vccd1 _00619_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_45_1688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12533_ net338 net330 _07463_ vssd1 vssd1 vccd1 vccd1 _07464_ sky130_fd_sc_hd__or3_1
XFILLER_0_87_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10594__A net1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14066__A net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11042__X _06015_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18040_ _03542_ net301 vssd1 vssd1 vccd1 vccd1 _03643_ sky130_fd_sc_hd__nand2_1
XFILLER_0_19_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15252_ net2287 net96 _01579_ net2524 vssd1 vssd1 vccd1 vccd1 _00560_ sky130_fd_sc_hd__a22o_1
XANTENNA__12005__B1 net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15742__A1 ag2.body\[337\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19541__CLK clknet_leaf_118_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12464_ net1631 _07420_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[1\] sky130_fd_sc_hd__and2_1
XFILLER_0_53_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_1500 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14203_ net973 ag2.body\[363\] vssd1 vssd1 vccd1 vccd1 _08364_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_10_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11415_ net1051 control.body\[855\] vssd1 vssd1 vccd1 vccd1 _06388_ sky130_fd_sc_hd__or2_1
XANTENNA__11202__B net1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15183_ net2207 net101 _01572_ control.body\[824\] vssd1 vssd1 vccd1 vccd1 _00498_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__09421__A1 ag2.goodColl vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12395_ _07282_ _07349_ _07359_ _07300_ vssd1 vssd1 vccd1 vccd1 net27 sky130_fd_sc_hd__a22o_1
XANTENNA__10567__B1 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14134_ net1027 ag2.body\[173\] vssd1 vssd1 vccd1 vccd1 _08295_ sky130_fd_sc_hd__xor2_1
XANTENNA__10031__A2 net1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11346_ _06315_ _06316_ _06317_ _06318_ vssd1 vssd1 vccd1 vccd1 _06319_ sky130_fd_sc_hd__or4_1
XANTENNA__17096__B net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09972__A2 _04427_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19991_ clknet_leaf_64_clk _00935_ net1474 vssd1 vssd1 vccd1 vccd1 ag2.body\[405\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_91_3088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_91_3099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11629__S net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14065_ _08211_ _08214_ _08225_ vssd1 vssd1 vccd1 vccd1 _08226_ sky130_fd_sc_hd__o21a_1
X_18942_ clknet_leaf_139_clk img_gen.tracker.next_frame\[380\] net1288 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[380\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_120_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11277_ ag2.body\[121\] net1211 vssd1 vssd1 vccd1 vccd1 _06250_ sky130_fd_sc_hd__xor2_1
X_13016_ net240 _07702_ _07703_ net1933 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[270\]
+ sky130_fd_sc_hd__a22o_1
X_10228_ ag2.body\[565\] net1101 vssd1 vssd1 vccd1 vccd1 _05201_ sky130_fd_sc_hd__xor2_1
X_18873_ clknet_leaf_22_clk img_gen.tracker.next_frame\[311\] net1358 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[311\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__15258__B1 net50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12033__B net1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17824_ net1514 net1508 vssd1 vssd1 vccd1 vccd1 _00004_ sky130_fd_sc_hd__or2_1
Xhold2 control.button4.Q\[1\] vssd1 vssd1 vccd1 vccd1 net1564 sky130_fd_sc_hd__dlygate4sd3_1
X_10159_ _05124_ _05128_ _05129_ _05131_ vssd1 vssd1 vccd1 vccd1 _05132_ sky130_fd_sc_hd__or4_1
XFILLER_0_101_1486 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_106_3541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_106_3552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11819__B1 net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_3563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17755_ _03045_ _03418_ _03426_ _03433_ vssd1 vssd1 vccd1 vccd1 _03434_ sky130_fd_sc_hd__and4_2
X_14967_ control.body\[1025\] net157 net51 control.body\[1017\] vssd1 vssd1 vccd1
+ vccd1 _00307_ sky130_fd_sc_hd__a22o_1
XANTENNA__14481__A1 net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14481__B2 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_3427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16706_ obsg2.obstacleArray\[75\] net500 net486 obsg2.obstacleArray\[74\] vssd1 vssd1
+ vccd1 vccd1 _02385_ sky130_fd_sc_hd__a22o_1
XFILLER_0_77_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17840__A net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_3438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13918_ ag2.body\[63\] net129 _08151_ ag2.body\[55\] vssd1 vssd1 vccd1 vccd1 _00144_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__16758__B1 net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_3449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17686_ _03361_ _03362_ _03364_ vssd1 vssd1 vccd1 vccd1 _03365_ sky130_fd_sc_hd__or3b_1
XFILLER_0_72_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14898_ net2186 net177 _01540_ net2313 vssd1 vssd1 vccd1 vccd1 _00245_ sky130_fd_sc_hd__a22o_1
XFILLER_0_134_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19425_ clknet_leaf_108_clk _00369_ net1434 vssd1 vssd1 vccd1 vccd1 control.body\[975\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16637_ net395 _02315_ _02314_ net361 vssd1 vssd1 vccd1 vccd1 _02316_ sky130_fd_sc_hd__a211o_1
X_13849_ ag2.body\[13\] net116 _08133_ net926 vssd1 vssd1 vccd1 vccd1 _00093_ sky130_fd_sc_hd__a22o_1
XFILLER_0_29_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16456__A _02057_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1201 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18639__CLK clknet_leaf_131_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13799__B net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19356_ clknet_leaf_102_clk _00300_ net1429 vssd1 vssd1 vccd1 vccd1 control.body\[1034\]
+ sky130_fd_sc_hd__dfrtp_1
X_16568_ obsg2.obstacleArray\[120\] obsg2.obstacleArray\[121\] net444 vssd1 vssd1
+ vccd1 vccd1 _02247_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_80_2770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_1600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_119_3946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12795__A1 net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_119_3957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18307_ net323 _03801_ _03800_ vssd1 vssd1 vccd1 vccd1 _03803_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_112_1571 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15519_ ag2.body\[539\] net156 _01609_ ag2.body\[531\] vssd1 vssd1 vccd1 vccd1 _00797_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_61_2180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16499_ obsg2.obstacleArray\[20\] obsg2.obstacleArray\[21\] obsg2.obstacleArray\[22\]
+ obsg2.obstacleArray\[23\] net458 net399 vssd1 vssd1 vccd1 vccd1 _02178_ sky130_fd_sc_hd__mux4_1
XFILLER_0_73_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19287_ clknet_leaf_98_clk _00231_ net1446 vssd1 vssd1 vccd1 vccd1 control.body\[1109\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_61_2191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09040_ ag2.body\[205\] vssd1 vssd1 vccd1 vccd1 _04065_ sky130_fd_sc_hd__inv_2
XFILLER_0_2_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18238_ _03679_ net35 vssd1 vssd1 vccd1 vccd1 _03758_ sky130_fd_sc_hd__nor2_1
XFILLER_0_115_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15733__B2 ag2.body\[337\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16930__B1 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16903__B net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18789__CLK clknet_leaf_13_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18169_ obsg2.obstacleArray\[81\] _03723_ net533 vssd1 vssd1 vccd1 vccd1 _01332_
+ sky130_fd_sc_hd__o21a_1
XANTENNA__14704__A net1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10009__A net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold402 img_gen.tracker.frame\[234\] vssd1 vssd1 vccd1 vccd1 net1964 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold413 img_gen.tracker.frame\[276\] vssd1 vssd1 vccd1 vccd1 net1975 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20200_ clknet_leaf_88_clk _01144_ net1454 vssd1 vssd1 vccd1 vccd1 ag2.body\[198\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_29_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold424 img_gen.tracker.frame\[213\] vssd1 vssd1 vccd1 vccd1 net1986 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09963__A2 net1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold435 img_gen.tracker.frame\[473\] vssd1 vssd1 vccd1 vccd1 net1997 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10951__B net1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold446 img_gen.tracker.frame\[299\] vssd1 vssd1 vccd1 vccd1 net2008 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_74_2574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold457 img_gen.tracker.frame\[378\] vssd1 vssd1 vccd1 vccd1 net2019 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20131_ clknet_leaf_81_clk _01075_ net1485 vssd1 vssd1 vccd1 vccd1 ag2.body\[257\]
+ sky130_fd_sc_hd__dfrtp_4
Xhold468 img_gen.tracker.frame\[260\] vssd1 vssd1 vccd1 vccd1 net2030 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11770__A2 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09942_ _03985_ net1054 _04908_ _04909_ _04910_ vssd1 vssd1 vccd1 vccd1 _04915_ sky130_fd_sc_hd__a2111o_1
Xhold479 img_gen.tracker.frame\[494\] vssd1 vssd1 vccd1 vccd1 net2041 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout904 net905 vssd1 vssd1 vccd1 vccd1 net904 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_70_2449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout915 net916 vssd1 vssd1 vccd1 vccd1 net915 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_42_1352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout926 ag2.body\[5\] vssd1 vssd1 vccd1 vccd1 net926 sky130_fd_sc_hd__buf_2
X_20062_ clknet_leaf_73_clk _01006_ net1501 vssd1 vssd1 vccd1 vccd1 ag2.body\[332\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_96_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout937 net941 vssd1 vssd1 vccd1 vccd1 net937 sky130_fd_sc_hd__buf_4
X_09873_ _04822_ _04830_ _04832_ _04845_ vssd1 vssd1 vccd1 vccd1 _04846_ sky130_fd_sc_hd__o22a_1
Xfanout948 net950 vssd1 vssd1 vccd1 vccd1 net948 sky130_fd_sc_hd__buf_4
Xfanout959 net961 vssd1 vssd1 vccd1 vccd1 net959 sky130_fd_sc_hd__buf_4
XANTENNA__16130__S net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1001_A net1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11782__B net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_2968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_87_2979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14472__A1 net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19414__CLK clknet_leaf_111_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14472__B2 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout559_A net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_2389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16749__B1 net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_1482 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14224__A1 net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout347_X net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1370_A net1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout726_A net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14224__B2 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1468_A net1478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11038__A1 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1089_X net1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09307_ sound_gen.osc1.count\[6\] _04325_ vssd1 vssd1 vccd1 vccd1 _04327_ sky130_fd_sc_hd__nand2_1
XANTENNA__17749__X _03428_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout514_X net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_4313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10923__A2_N net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_4324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_1408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09238_ net869 vssd1 vssd1 vccd1 vccd1 _04263_ sky130_fd_sc_hd__clkinv_4
XANTENNA__20541__CLK clknet_leaf_105_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_1530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_20_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17909__B _03533_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_20_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_1552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16813__B net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11022__B net1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09169_ ag2.body\[530\] vssd1 vssd1 vccd1 vccd1 _04194_ sky130_fd_sc_hd__inv_2
XANTENNA__14614__A net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11200_ net918 net921 net913 net909 vssd1 vssd1 vccd1 vccd1 _06173_ sky130_fd_sc_hd__o211a_2
X_12180_ net1174 ag2.apple_cord\[2\] vssd1 vssd1 vccd1 vccd1 _07152_ sky130_fd_sc_hd__xor2_1
XANTENNA_fanout883_X net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11131_ net1100 control.body\[869\] vssd1 vssd1 vccd1 vccd1 _06104_ sky130_fd_sc_hd__or2_1
XFILLER_0_124_1464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20329_ clknet_leaf_112_clk track.current_collision net1424 vssd1 vssd1 vccd1 vccd1
+ track.last_collision sky130_fd_sc_hd__dfrtp_1
XANTENNA__14151__A1_N net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_4253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_4264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold980 control.body\[672\] vssd1 vssd1 vccd1 vccd1 net2542 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_120_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold991 control.body\[1072\] vssd1 vssd1 vccd1 vccd1 net2553 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11062_ ag2.body\[438\] net1079 vssd1 vssd1 vccd1 vccd1 _06035_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_125_4128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_125_4139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_34_1356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10013_ _04981_ _04985_ vssd1 vssd1 vccd1 vccd1 _04986_ sky130_fd_sc_hd__nor2_2
X_15870_ ag2.body\[228\] net201 _01647_ ag2.body\[220\] vssd1 vssd1 vccd1 vccd1 _01110_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_34_1367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10721__B1 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14821_ net1013 ag2.body\[159\] vssd1 vssd1 vccd1 vccd1 _01492_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09443__A net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15164__B net63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13236__Y _07807_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_320 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10589__A net1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17540_ ag2.body\[320\] net741 net702 ag2.body\[326\] vssd1 vssd1 vccd1 vccd1 _03219_
+ sky130_fd_sc_hd__a22o_1
X_14752_ net975 ag2.body\[107\] vssd1 vssd1 vccd1 vccd1 _08913_ sky130_fd_sc_hd__xor2_1
X_11964_ img_gen.tracker.frame\[481\] net616 net546 img_gen.tracker.frame\[487\] vssd1
+ vssd1 vccd1 vccd1 _06936_ sky130_fd_sc_hd__o22a_1
XFILLER_0_98_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__20071__CLK clknet_leaf_73_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13703_ track.highScore\[3\] _04642_ _08026_ track.highScore\[4\] vssd1 vssd1 vccd1
+ vccd1 _08044_ sky130_fd_sc_hd__a22oi_1
X_10915_ ag2.body\[463\] net1055 vssd1 vssd1 vccd1 vccd1 _05888_ sky130_fd_sc_hd__xnor2_1
X_17471_ _03148_ _03149_ vssd1 vssd1 vccd1 vccd1 _03150_ sky130_fd_sc_hd__nand2_1
X_14683_ net808 ag2.body\[93\] ag2.body\[94\] net804 vssd1 vssd1 vccd1 vccd1 _08844_
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_6_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11895_ net472 _06866_ vssd1 vssd1 vccd1 vccd1 _06867_ sky130_fd_sc_hd__nand2_1
XANTENNA__10101__B net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14348__X _08509_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19210_ clknet_leaf_85_clk _00154_ net1463 vssd1 vssd1 vccd1 vccd1 ag2.body\[73\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_54_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18194__C _03703_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13634_ control.divider.count\[12\] _07995_ vssd1 vssd1 vccd1 vccd1 _07997_ sky130_fd_sc_hd__and2_1
X_16422_ _02075_ _02083_ _02057_ vssd1 vssd1 vccd1 vccd1 _02101_ sky130_fd_sc_hd__a21bo_1
X_10846_ _05814_ _05816_ _05817_ _05818_ vssd1 vssd1 vccd1 vccd1 _05819_ sky130_fd_sc_hd__or4_1
XFILLER_0_67_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_15_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16353_ obsg2.obstacleArray\[7\] net414 _02031_ net416 vssd1 vssd1 vccd1 vccd1 _02032_
+ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_15_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19141_ clknet_leaf_139_clk net1570 net1289 vssd1 vssd1 vccd1 vccd1 img_gen.control.button5.Q\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_13565_ ssdec1.in\[2\] ssdec1.in\[3\] vssd1 vssd1 vccd1 vccd1 _07944_ sky130_fd_sc_hd__nand2_1
XFILLER_0_26_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_1576 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10777_ _05746_ _05747_ _05748_ _05749_ vssd1 vssd1 vccd1 vccd1 _05750_ sky130_fd_sc_hd__or4_1
XANTENNA__18931__CLK clknet_leaf_141_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17165__B1 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11213__A net1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15304_ net2386 net75 _01586_ net2418 vssd1 vssd1 vccd1 vccd1 _00605_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_97_3275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19072_ clknet_leaf_28_clk img_gen.tracker.next_frame\[510\] net1335 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[510\] sky130_fd_sc_hd__dfrtp_1
X_12516_ net2082 net650 _07455_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[18\]
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_114_3810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16284_ net372 _01962_ _01959_ _01911_ vssd1 vssd1 vccd1 vccd1 _01963_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_97_3286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_1320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13496_ net664 _07910_ vssd1 vssd1 vccd1 vccd1 _07911_ sky130_fd_sc_hd__nor2_1
XFILLER_0_48_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16912__B1 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_867 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18023_ net45 _03631_ vssd1 vssd1 vccd1 vccd1 _03632_ sky130_fd_sc_hd__nor2_1
X_15235_ control.body\[799\] net96 _01577_ net2267 vssd1 vssd1 vccd1 vccd1 _00545_
+ sky130_fd_sc_hd__a22o_1
X_12447_ img_gen.updater.commands.rR1.rainbowRNG\[14\] _07319_ _07338_ _07397_ _07407_
+ vssd1 vssd1 vccd1 vccd1 _07408_ sky130_fd_sc_hd__a221o_1
XFILLER_0_65_1330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_max_cap357_A _02228_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14524__A net1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09618__A net1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15166_ control.body\[849\] net103 _01570_ net2435 vssd1 vssd1 vccd1 vccd1 _00483_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11867__B net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12378_ img_gen.updater.commands.count\[7\] _07211_ _07341_ vssd1 vssd1 vccd1 vccd1
+ _07343_ sky130_fd_sc_hd__a21o_1
XFILLER_0_26_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10771__B net1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11070__A2_N net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14117_ net832 ag2.body\[569\] ag2.body\[575\] net791 _08274_ vssd1 vssd1 vccd1 vccd1
+ _08278_ sky130_fd_sc_hd__o221ai_1
XFILLER_0_107_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17835__A net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11329_ net1217 control.body\[656\] vssd1 vssd1 vccd1 vccd1 _06302_ sky130_fd_sc_hd__xor2_1
X_19974_ clknet_leaf_63_clk _00918_ net1470 vssd1 vssd1 vccd1 vccd1 ag2.body\[420\]
+ sky130_fd_sc_hd__dfrtp_4
X_15097_ net2603 net145 _01563_ net2154 vssd1 vssd1 vccd1 vccd1 _00421_ sky130_fd_sc_hd__a22o_1
XFILLER_0_5_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14048_ net817 ag2.body\[187\] ag2.body\[188\] net811 _08207_ vssd1 vssd1 vccd1 vccd1
+ _08209_ sky130_fd_sc_hd__o221a_1
X_18925_ clknet_leaf_140_clk img_gen.tracker.next_frame\[363\] net1290 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[363\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__17554__B net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_3603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_1559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_108_3614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_3625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12701__A1 net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11883__A net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18856_ clknet_leaf_18_clk img_gen.tracker.next_frame\[294\] net1322 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[294\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__10712__B1 net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19142__RESET_B net1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17807_ _08110_ net56 vssd1 vssd1 vccd1 vccd1 _03476_ sky130_fd_sc_hd__nor2_1
XANTENNA__17640__B2 net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14454__A1 net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18787_ clknet_leaf_13_clk img_gen.tracker.next_frame\[225\] net1284 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[225\] sky130_fd_sc_hd__dfrtp_1
X_15999_ net930 _01676_ vssd1 vssd1 vccd1 vccd1 _01678_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_55_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14454__B2 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17738_ _02632_ _02633_ _02642_ _03416_ _02601_ vssd1 vssd1 vccd1 vccd1 _03417_ sky130_fd_sc_hd__o311a_1
XTAP_TAPCELL_ROW_82_2810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19587__CLK clknet_leaf_118_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_2821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18196__A2 _03703_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_2832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17669_ ag2.body\[454\] net939 vssd1 vssd1 vccd1 vccd1 _03348_ sky130_fd_sc_hd__xor2_1
XANTENNA__14206__A1 net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_2231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14206__B2 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15403__B1 _01581_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_2242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10011__B _04791_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_63_2253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19408_ clknet_leaf_103_clk _00352_ net1429 vssd1 vssd1 vccd1 vccd1 control.body\[990\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__20564__CLK clknet_leaf_43_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19339_ clknet_leaf_100_clk _00283_ net1443 vssd1 vssd1 vccd1 vccd1 control.body\[1049\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_50_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17569__X _03248_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11123__A net1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09023_ ag2.body\[158\] vssd1 vssd1 vccd1 vccd1 _04048_ sky130_fd_sc_hd__inv_2
XFILLER_0_116_889 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_2636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11991__A2 net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_2647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14434__A net1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout307_A _07445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1049_A net1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14390__B1 ag2.body\[303\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold210 img_gen.tracker.frame\[458\] vssd1 vssd1 vccd1 vccd1 net1772 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_4_1__f_clk_X clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_2057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11777__B net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_2068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold221 img_gen.tracker.frame\[497\] vssd1 vssd1 vccd1 vccd1 net1783 sky130_fd_sc_hd__dlygate4sd3_1
Xhold232 img_gen.tracker.frame\[415\] vssd1 vssd1 vccd1 vccd1 net1794 sky130_fd_sc_hd__dlygate4sd3_1
Xhold243 img_gen.tracker.frame\[308\] vssd1 vssd1 vccd1 vccd1 net1805 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11743__A2 net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold254 img_gen.tracker.frame\[351\] vssd1 vssd1 vccd1 vccd1 net1816 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__16131__A1 net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold265 img_gen.tracker.frame\[89\] vssd1 vssd1 vccd1 vccd1 net1827 sky130_fd_sc_hd__dlygate4sd3_1
Xhold276 img_gen.tracker.frame\[119\] vssd1 vssd1 vccd1 vccd1 net1838 sky130_fd_sc_hd__dlygate4sd3_1
Xhold287 img_gen.tracker.frame\[173\] vssd1 vssd1 vccd1 vccd1 net1849 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1216_A net1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout701 net702 vssd1 vssd1 vccd1 vccd1 net701 sky130_fd_sc_hd__buf_4
X_09925_ ag2.body\[317\] net1116 vssd1 vssd1 vccd1 vccd1 _04898_ sky130_fd_sc_hd__xor2_1
Xfanout712 net714 vssd1 vssd1 vccd1 vccd1 net712 sky130_fd_sc_hd__buf_2
Xhold298 img_gen.tracker.frame\[516\] vssd1 vssd1 vccd1 vccd1 net1860 sky130_fd_sc_hd__dlygate4sd3_1
X_20114_ clknet_leaf_80_clk _01058_ net1487 vssd1 vssd1 vccd1 vccd1 ag2.body\[272\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__16209__B_N net860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout723 net725 vssd1 vssd1 vccd1 vccd1 net723 sky130_fd_sc_hd__buf_4
XANTENNA__17464__B net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14693__A1 net993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout734 net736 vssd1 vssd1 vccd1 vccd1 net734 sky130_fd_sc_hd__buf_4
XANTENNA__14693__B2 net1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout676_A net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout745 net746 vssd1 vssd1 vccd1 vccd1 net745 sky130_fd_sc_hd__buf_4
X_20045_ clknet_leaf_68_clk _00989_ net1495 vssd1 vssd1 vccd1 vccd1 ag2.body\[347\]
+ sky130_fd_sc_hd__dfrtp_4
Xfanout756 net757 vssd1 vssd1 vccd1 vccd1 net756 sky130_fd_sc_hd__buf_4
X_09856_ _04772_ _04828_ vssd1 vssd1 vccd1 vccd1 _04829_ sky130_fd_sc_hd__nand2_1
Xfanout767 net768 vssd1 vssd1 vccd1 vccd1 net767 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout1004_X net1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout778 net782 vssd1 vssd1 vccd1 vccd1 net778 sky130_fd_sc_hd__clkbuf_8
Xfanout789 _04227_ vssd1 vssd1 vccd1 vccd1 net789 sky130_fd_sc_hd__buf_4
XFILLER_0_77_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09787_ net1204 control.body\[945\] vssd1 vssd1 vccd1 vccd1 _04760_ sky130_fd_sc_hd__xor2_1
XANTENNA_fanout843_A net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout464_X net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15642__B1 _01623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_137_4500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout631_X net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10696__X _05669_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15712__B net67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_137_4511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17395__B1 net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18954__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout729_X net729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10700_ ag2.body\[23\] net1054 vssd1 vssd1 vccd1 vccd1 _05673_ sky130_fd_sc_hd__or2_1
XANTENNA__09710__B net1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15945__A1 ag2.body\[167\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11680_ net1225 net1199 vssd1 vssd1 vccd1 vccd1 _06652_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_138_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_1603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12759__A1 net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10631_ net1192 control.body\[665\] vssd1 vssd1 vccd1 vccd1 _05604_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_27_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_23_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_119 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_23_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13350_ net249 _07852_ _07853_ net1953 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[454\]
+ sky130_fd_sc_hd__a22o_1
X_10562_ ag2.body\[514\] net775 _05533_ _05534_ vssd1 vssd1 vccd1 vccd1 _05535_ sky130_fd_sc_hd__a211o_1
XANTENNA__17639__B net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_101_Left_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12301_ _07221_ _07267_ vssd1 vssd1 vccd1 vccd1 _07268_ sky130_fd_sc_hd__and2_1
XANTENNA__11982__A2 net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13281_ net255 _07825_ _07826_ net1915 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[412\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__16370__A1 _01918_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10493_ ag2.body\[551\] net1059 vssd1 vssd1 vccd1 vccd1 _05466_ sky130_fd_sc_hd__xnor2_1
XANTENNA__14344__A net1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15020_ _04551_ net59 vssd1 vssd1 vccd1 vccd1 _01554_ sky130_fd_sc_hd__nor2_4
XFILLER_0_122_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12232_ _07195_ _07201_ img_gen.updater.commands.cmd_num\[3\] _07188_ vssd1 vssd1
+ vccd1 vccd1 _07202_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_27_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11687__B net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14920__A2 net171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11734__A2 net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16122__A1 net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12163_ img_gen.tracker.frame\[396\] net617 vssd1 vssd1 vccd1 vccd1 _07135_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_36_1418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_1429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11114_ _06080_ _06084_ _06085_ _06086_ vssd1 vssd1 vccd1 vccd1 _06087_ sky130_fd_sc_hd__and4_4
XTAP_TAPCELL_ROW_9_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16971_ _02648_ _02643_ _02645_ _02649_ vssd1 vssd1 vccd1 vccd1 _02650_ sky130_fd_sc_hd__or4bb_1
X_12094_ net1215 net1190 img_gen.tracker.frame\[357\] vssd1 vssd1 vccd1 vccd1 _07066_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_120_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14684__A1 net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14684__B2 net1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18710_ clknet_leaf_143_clk img_gen.tracker.next_frame\[148\] net1255 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[148\] sky130_fd_sc_hd__dfrtp_1
X_15922_ ag2.body\[177\] net124 _01654_ ag2.body\[169\] vssd1 vssd1 vccd1 vccd1 _01155_
+ sky130_fd_sc_hd__a22o_1
X_11045_ _05884_ _05908_ _05936_ _06017_ vssd1 vssd1 vccd1 vccd1 _06018_ sky130_fd_sc_hd__or4_1
X_19690_ clknet_leaf_136_clk _00634_ net1300 vssd1 vssd1 vccd1 vccd1 control.body\[696\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_36_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16425__A2 _02103_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18641_ clknet_leaf_131_clk img_gen.tracker.next_frame\[79\] net1314 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[79\] sky130_fd_sc_hd__dfrtp_1
X_15853_ ag2.body\[245\] net174 _01645_ ag2.body\[237\] vssd1 vssd1 vccd1 vccd1 _01095_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_56_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14804_ net830 ag2.body\[290\] ag2.body\[291\] net823 vssd1 vssd1 vccd1 vccd1 _01475_
+ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__11208__A _04446_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__20587__CLK clknet_leaf_105_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18572_ clknet_leaf_15_clk img_gen.tracker.next_frame\[10\] net1312 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[10\] sky130_fd_sc_hd__dfrtp_1
X_15784_ ag2.body\[311\] net210 _01638_ ag2.body\[303\] vssd1 vssd1 vccd1 vccd1 _01033_
+ sky130_fd_sc_hd__a22o_1
X_12996_ net279 _07691_ _07692_ net2030 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[260\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__14987__A2 net154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20140__RESET_B net1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_4_12__f_clk_X clknet_4_12__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17523_ ag2.body\[482\] net724 net717 ag2.body\[483\] vssd1 vssd1 vccd1 vccd1 _03202_
+ sky130_fd_sc_hd__a22o_1
X_14735_ net1004 ag2.body\[328\] vssd1 vssd1 vccd1 vccd1 _08896_ sky130_fd_sc_hd__xor2_1
X_11947_ img_gen.tracker.frame\[130\] net585 net547 img_gen.tracker.frame\[127\] _06918_
+ vssd1 vssd1 vccd1 vccd1 _06919_ sky130_fd_sc_hd__o221a_1
XFILLER_0_74_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17454_ ag2.body\[436\] net960 vssd1 vssd1 vccd1 vccd1 _03133_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_15_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11670__A1 net1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14666_ net820 ag2.body\[523\] ag2.body\[525\] net809 _08826_ vssd1 vssd1 vccd1 vccd1
+ _08827_ sky130_fd_sc_hd__a221o_1
XFILLER_0_129_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_3337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11878_ _06831_ _06837_ _06844_ _06849_ net468 net438 vssd1 vssd1 vccd1 vccd1 _06850_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__15936__B2 ag2.body\[166\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_3348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13617_ _07985_ _07986_ vssd1 vssd1 vccd1 vccd1 control.divider.next_count\[5\] sky130_fd_sc_hd__nor2_1
XFILLER_0_117_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16405_ net354 _02055_ vssd1 vssd1 vccd1 vccd1 _02084_ sky130_fd_sc_hd__nand2_1
X_10829_ ag2.body\[305\] net1212 vssd1 vssd1 vccd1 vccd1 _05802_ sky130_fd_sc_hd__xor2_1
X_14597_ net845 ag2.body\[304\] ag2.body\[310\] net803 _08755_ vssd1 vssd1 vccd1 vccd1
+ _08758_ sky130_fd_sc_hd__o221ai_1
X_17385_ _03059_ _03060_ _03062_ _03063_ vssd1 vssd1 vccd1 vccd1 _03064_ sky130_fd_sc_hd__a22o_1
XFILLER_0_138_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17428__A2_N net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19124_ clknet_leaf_141_clk img_gen.tracker.next_frame\[562\] net1294 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[562\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_32_1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16336_ obsg2.obstacleArray\[84\] obsg2.obstacleArray\[85\] net411 vssd1 vssd1 vccd1
+ vccd1 _02015_ sky130_fd_sc_hd__mux2_1
X_13548_ net2069 net659 _07929_ _07930_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[575\]
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_43_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16267_ net371 _01941_ _01945_ net368 vssd1 vssd1 vccd1 vccd1 _01946_ sky130_fd_sc_hd__o211a_1
X_19055_ clknet_leaf_8_clk img_gen.tracker.next_frame\[493\] net1273 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[493\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_124_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13479_ net276 _07902_ _07903_ net1982 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[533\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__10782__A net1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14254__A net1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18006_ net345 net299 _03573_ vssd1 vssd1 vccd1 vccd1 _03619_ sky130_fd_sc_hd__and3_1
XFILLER_0_112_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15218_ _04587_ net53 vssd1 vssd1 vccd1 vccd1 _01576_ sky130_fd_sc_hd__nor2_2
XANTENNA__09918__A2 net1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16198_ _01875_ _01876_ net377 vssd1 vssd1 vccd1 vccd1 _01877_ sky130_fd_sc_hd__mux2_1
XANTENNA__11186__B1 net1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_71_2500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11725__A2 net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12922__A1 net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15149_ control.body\[866\] net105 _01568_ control.body\[858\] vssd1 vssd1 vccd1
+ vccd1 _00468_ sky130_fd_sc_hd__a22o_1
XFILLER_0_22_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18827__CLK clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19957_ clknet_leaf_45_clk _00901_ net1381 vssd1 vssd1 vccd1 vccd1 ag2.body\[435\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_103_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17284__B net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20299__RESET_B net1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09710_ ag2.body\[242\] net1182 vssd1 vssd1 vccd1 vccd1 _04683_ sky130_fd_sc_hd__or2_1
X_18908_ clknet_leaf_144_clk img_gen.tracker.next_frame\[346\] net1251 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[346\] sky130_fd_sc_hd__dfrtp_1
X_19888_ clknet_leaf_87_clk _00832_ net1460 vssd1 vssd1 vccd1 vccd1 ag2.body\[510\]
+ sky130_fd_sc_hd__dfrtp_4
X_09641_ net893 _04602_ _04492_ vssd1 vssd1 vccd1 vccd1 _04614_ sky130_fd_sc_hd__o21ai_2
X_18839_ clknet_leaf_4_clk img_gen.tracker.next_frame\[277\] net1277 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[277\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_69_2440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15624__B1 _01621_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15372__X _01594_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_2304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09572_ _04065_ net1114 net1064 _04067_ _04544_ vssd1 vssd1 vccd1 vccd1 _04545_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_65_2315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_312 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09811__A net1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12989__A1 net254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14429__A net997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout257_A net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13333__A net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09530__B _04494_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10676__B net1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17129__B1 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout424_A net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12205__A3 _06986_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_78_2709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1166_A ag2.y\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_2108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20594_ net1526 vssd1 vssd1 vccd1 vccd1 gpio_oeb[6] sky130_fd_sc_hd__buf_2
XANTENNA__10963__Y _05936_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_2119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12891__B _07639_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11964__A2 net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14164__A net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1333_A net1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_372 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09006_ ag2.body\[126\] vssd1 vssd1 vccd1 vccd1 _04031_ sky130_fd_sc_hd__inv_2
XANTENNA__13166__A1 net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout793_A net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17301__B1 net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1500_A net1502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1121_X net1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1219_X net1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09545__X _04518_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout960_A net961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1507 net1508 vssd1 vssd1 vccd1 vccd1 net1507 sky130_fd_sc_hd__buf_1
Xfanout520 net528 vssd1 vssd1 vccd1 vccd1 net520 sky130_fd_sc_hd__buf_2
XANTENNA__14666__A1 net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout531 net533 vssd1 vssd1 vccd1 vccd1 net531 sky130_fd_sc_hd__clkbuf_4
XANTENNA__14666__B2 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1591 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout542 net543 vssd1 vssd1 vccd1 vccd1 net542 sky130_fd_sc_hd__clkbuf_4
XANTENNA__17762__X _03441_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09908_ ag2.body\[132\] net1141 vssd1 vssd1 vccd1 vccd1 _04881_ sky130_fd_sc_hd__or2_1
Xfanout553 _06652_ vssd1 vssd1 vccd1 vccd1 net553 sky130_fd_sc_hd__buf_2
Xfanout564 net567 vssd1 vssd1 vccd1 vccd1 net564 sky130_fd_sc_hd__buf_2
Xfanout575 _06649_ vssd1 vssd1 vccd1 vccd1 net575 sky130_fd_sc_hd__clkbuf_4
Xfanout586 net592 vssd1 vssd1 vccd1 vccd1 net586 sky130_fd_sc_hd__buf_2
XANTENNA__12141__A2 net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20028_ clknet_leaf_67_clk _00972_ net1477 vssd1 vssd1 vccd1 vccd1 ag2.body\[362\]
+ sky130_fd_sc_hd__dfrtp_4
X_09839_ net1204 control.body\[921\] vssd1 vssd1 vccd1 vccd1 _04812_ sky130_fd_sc_hd__nand2_1
Xfanout597 net598 vssd1 vssd1 vccd1 vccd1 net597 sky130_fd_sc_hd__buf_2
XFILLER_0_96_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout846_X net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14418__A1 net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14418__B2 net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11028__A net1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12850_ net261 _07625_ _07626_ net2023 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[181\]
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_48_1801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_29_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11801_ net468 _06735_ _06730_ net466 vssd1 vssd1 vccd1 vccd1 _06773_ sky130_fd_sc_hd__o211a_1
XFILLER_0_68_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11970__B net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12781_ net239 _07593_ _07594_ net2057 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[144\]
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_29_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14339__A net1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14520_ net1003 _04103_ ag2.body\[317\] net810 vssd1 vssd1 vccd1 vccd1 _08681_ sky130_fd_sc_hd__a22o_1
XFILLER_0_84_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11315__X _06288_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19132__CLK clknet_leaf_141_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11732_ net565 _06693_ net470 vssd1 vssd1 vccd1 vccd1 _06704_ sky130_fd_sc_hd__a21o_1
XFILLER_0_138_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14451_ _08604_ _08605_ _08607_ _08609_ vssd1 vssd1 vccd1 vccd1 _08612_ sky130_fd_sc_hd__a211o_1
X_11663_ net1118 net1095 vssd1 vssd1 vccd1 vccd1 _06635_ sky130_fd_sc_hd__or2_1
XANTENNA__16591__A1 net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_94_3201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13402_ net238 net312 _07553_ _07873_ net1664 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[486\]
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_68_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10614_ _05559_ _05572_ _05573_ _05586_ vssd1 vssd1 vccd1 vccd1 _05587_ sky130_fd_sc_hd__o22a_1
X_17170_ _02839_ _02840_ _02842_ _02843_ _02848_ vssd1 vssd1 vccd1 vccd1 _02849_ sky130_fd_sc_hd__a221o_1
X_14382_ net992 ag2.body\[297\] vssd1 vssd1 vccd1 vccd1 _08543_ sky130_fd_sc_hd__xor2_1
X_11594_ obsg2.obstacleArray\[10\] net633 net509 obsg2.obstacleArray\[14\] net759
+ vssd1 vssd1 vccd1 vccd1 _06567_ sky130_fd_sc_hd__o221a_1
X_16121_ obsg2.obstacleArray\[78\] obsg2.obstacleArray\[79\] net423 vssd1 vssd1 vccd1
+ vccd1 _01800_ sky130_fd_sc_hd__mux2_1
XFILLER_0_106_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13333_ net664 _07846_ vssd1 vssd1 vccd1 vccd1 _07847_ sky130_fd_sc_hd__nor2_1
XANTENNA__19834__RESET_B net1414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10545_ ag2.body\[228\] net1136 vssd1 vssd1 vccd1 vccd1 _05518_ sky130_fd_sc_hd__nand2_1
XANTENNA__12146__X _07118_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_130_clk clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_130_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_64_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17540__B1 net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16052_ _01720_ _01730_ vssd1 vssd1 vccd1 vccd1 _01731_ sky130_fd_sc_hd__and2b_1
XFILLER_0_49_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13264_ net672 _07819_ vssd1 vssd1 vccd1 vccd1 _07820_ sky130_fd_sc_hd__nor2_1
X_10476_ _04614_ _05448_ _05435_ vssd1 vssd1 vccd1 vccd1 _05449_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_51_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_1480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15003_ net2569 net152 _01552_ control.body\[984\] vssd1 vssd1 vccd1 vccd1 _00338_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12904__A1 net245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11707__A2 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12215_ img_gen.control.current\[0\] _07182_ _07179_ net677 vssd1 vssd1 vccd1 vccd1
+ _07186_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_32_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10107__A net1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13195_ net289 _07785_ _07786_ net2014 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[365\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_104_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19811_ clknet_leaf_125_clk _00755_ net1410 vssd1 vssd1 vccd1 vccd1 ag2.body\[577\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_88_3005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12146_ _07115_ _07116_ _07117_ _07114_ vssd1 vssd1 vccd1 vccd1 _07118_ sky130_fd_sc_hd__a31o_1
XFILLER_0_138_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_88_3016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14657__A1 net1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_1407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10391__A1 net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14657__B2 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19742_ clknet_leaf_128_clk _00686_ net1325 vssd1 vssd1 vccd1 vccd1 control.body\[652\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_1529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16954_ ag2.body\[292\] net964 vssd1 vssd1 vccd1 vccd1 _02633_ sky130_fd_sc_hd__xor2_4
X_12077_ img_gen.tracker.frame\[132\] net629 net594 img_gen.tracker.frame\[141\] _07048_
+ vssd1 vssd1 vccd1 vccd1 _07049_ sky130_fd_sc_hd__a221o_1
XANTENNA__20312__Q ag2.randCord\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12132__A2 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15905_ ag2.body\[195\] net129 _01651_ ag2.body\[187\] vssd1 vssd1 vccd1 vccd1 _01141_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_75_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11028_ net1061 control.body\[1047\] vssd1 vssd1 vccd1 vccd1 _06001_ sky130_fd_sc_hd__or2_1
X_19673_ clknet_leaf_119_clk _00617_ net1386 vssd1 vssd1 vccd1 vccd1 control.body\[727\]
+ sky130_fd_sc_hd__dfrtp_1
X_16885_ ag2.body\[23\] net688 net722 ag2.body\[18\] vssd1 vssd1 vccd1 vccd1 _02564_
+ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__11340__B1 _06312_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18624_ clknet_leaf_0_clk img_gen.tracker.next_frame\[62\] net1248 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[62\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__10694__A2 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15836_ ag2.body\[262\] net201 net49 ag2.body\[254\] vssd1 vssd1 vccd1 vccd1 _01080_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_99_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12976__B net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18555_ clknet_leaf_43_clk _00081_ net1378 vssd1 vssd1 vccd1 vccd1 control.fsm.temp\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_15767_ _04897_ _01631_ vssd1 vssd1 vccd1 vccd1 _01637_ sky130_fd_sc_hd__and2b_2
X_12979_ net225 _07684_ _07685_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[251\]
+ sky130_fd_sc_hd__o21bai_1
X_17506_ ag2.body\[234\] net726 net933 _04074_ _03184_ vssd1 vssd1 vccd1 vccd1 _03185_
+ sky130_fd_sc_hd__a221o_1
X_14718_ net1033 ag2.body\[341\] vssd1 vssd1 vccd1 vccd1 _08879_ sky130_fd_sc_hd__nand2_1
XFILLER_0_86_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18486_ net1516 net1510 vssd1 vssd1 vccd1 vccd1 _00017_ sky130_fd_sc_hd__or2_1
X_15698_ ag2.body\[379\] net137 _01628_ ag2.body\[371\] vssd1 vssd1 vccd1 vccd1 _00957_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_34_1468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10496__B net1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17437_ ag2.body\[148\] net713 net693 ag2.body\[151\] _03115_ vssd1 vssd1 vccd1 vccd1
+ _03116_ sky130_fd_sc_hd__o221a_1
XFILLER_0_129_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14649_ _08805_ _08806_ _08807_ _08809_ vssd1 vssd1 vccd1 vccd1 _08810_ sky130_fd_sc_hd__or4_1
XFILLER_0_69_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_120_Right_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_16 _03446_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_27 _03442_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13396__A1 net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_38 _08924_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17368_ _03967_ _03046_ vssd1 vssd1 vccd1 vccd1 _03047_ sky130_fd_sc_hd__nor2_1
XFILLER_0_15_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19107_ clknet_leaf_1_clk img_gen.tracker.next_frame\[545\] net1244 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[545\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_15_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16319_ obsg2.obstacleArray\[68\] net409 vssd1 vssd1 vccd1 vccd1 _01998_ sky130_fd_sc_hd__or2_1
XFILLER_0_12_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_121_clk clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_121_clk
+ sky130_fd_sc_hd__clkbuf_8
X_17299_ ag2.body\[347\] net855 vssd1 vssd1 vccd1 vccd1 _02978_ sky130_fd_sc_hd__or2_1
XFILLER_0_82_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19038_ clknet_leaf_6_clk img_gen.tracker.next_frame\[476\] net1264 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[476\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14712__A net1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16403__S net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20409__RESET_B net1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14648__A1 net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15845__B1 _01644_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14648__B2 net1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17924__A_N net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13328__A net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12123__A2 net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13320__A1 net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1351 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout374_A net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09624_ _04589_ _04590_ _04594_ _04596_ vssd1 vssd1 vccd1 vccd1 _04597_ sky130_fd_sc_hd__or4b_2
XANTENNA__19155__CLK clknet_leaf_52_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16496__S1 net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12886__B _07639_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09541__A net1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11790__B net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09555_ net1193 control.body\[721\] vssd1 vssd1 vccd1 vccd1 _04528_ sky130_fd_sc_hd__xor2_1
XANTENNA__15262__B net58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_1622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_1562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout541_A net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout162_X net162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout639_A net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14820__B2 net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09486_ ag2.body\[368\] net1234 vssd1 vssd1 vccd1 vccd1 _04459_ sky130_fd_sc_hd__xor2_1
XFILLER_0_93_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16573__A1 net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1450_A net1451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout427_X net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout806_A net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1169_X net1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11398__B1 _05133_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11937__A2 net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16325__A1 net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20577_ clknet_leaf_107_clk sound_gen.osc1.at_max_nxt _00041_ vssd1 vssd1 vccd1 vccd1
+ sound_gen.at_max sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_112_clk clknet_4_10__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_112_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__19245__RESET_B net1482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10330_ control.body_update.curr_length\[1\] net923 _04554_ _05302_ vssd1 vssd1 vccd1
+ vccd1 _05303_ sky130_fd_sc_hd__a31o_1
XFILLER_0_61_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1388 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout796_X net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10261_ _05224_ _05225_ _05229_ _05233_ vssd1 vssd1 vccd1 vccd1 _05234_ sky130_fd_sc_hd__and4_1
XANTENNA_fanout1503_X net1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12000_ img_gen.tracker.frame\[445\] net614 net578 img_gen.tracker.frame\[454\] _06971_
+ vssd1 vssd1 vccd1 vccd1 _06972_ sky130_fd_sc_hd__o221a_1
XFILLER_0_121_1220 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10192_ ag2.body\[114\] net1186 vssd1 vssd1 vccd1 vccd1 _05165_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout963_X net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19193__Q ag2.body\[56\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14639__A1 net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1304 net1306 vssd1 vssd1 vccd1 vccd1 net1304 sky130_fd_sc_hd__clkbuf_4
XANTENNA__14639__B2 net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1315 net1324 vssd1 vssd1 vccd1 vccd1 net1315 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_100_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13238__A net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1326 net1327 vssd1 vssd1 vccd1 vccd1 net1326 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09435__B net1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1337 net1338 vssd1 vssd1 vccd1 vccd1 net1337 sky130_fd_sc_hd__clkbuf_2
Xfanout1348 net1351 vssd1 vssd1 vccd1 vccd1 net1348 sky130_fd_sc_hd__clkbuf_4
Xfanout350 net351 vssd1 vssd1 vccd1 vccd1 net350 sky130_fd_sc_hd__buf_2
Xfanout361 _02222_ vssd1 vssd1 vccd1 vccd1 net361 sky130_fd_sc_hd__clkbuf_4
Xfanout1359 net1362 vssd1 vssd1 vccd1 vccd1 net1359 sky130_fd_sc_hd__clkbuf_4
Xfanout372 _01907_ vssd1 vssd1 vccd1 vccd1 net372 sky130_fd_sc_hd__buf_2
X_13951_ ag2.body\[92\] net191 _08155_ ag2.body\[84\] vssd1 vssd1 vccd1 vccd1 _00173_
+ sky130_fd_sc_hd__a22o_1
Xfanout383 _06822_ vssd1 vssd1 vccd1 vccd1 net383 sky130_fd_sc_hd__buf_2
Xfanout394 net395 vssd1 vssd1 vccd1 vccd1 net394 sky130_fd_sc_hd__clkbuf_4
XANTENNA__17589__B1 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16549__A net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17053__A2 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12902_ _07453_ net339 net386 vssd1 vssd1 vccd1 vccd1 _07650_ sky130_fd_sc_hd__and3b_1
X_16670_ _02346_ _02347_ _02348_ _02216_ net362 vssd1 vssd1 vccd1 vccd1 _02349_ sky130_fd_sc_hd__a221o_1
X_13882_ ag2.body\[31\] net115 _08147_ ag2.body\[23\] vssd1 vssd1 vccd1 vccd1 _00112_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_9_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09451__A net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15621_ ag2.body\[454\] net123 _01613_ ag2.body\[446\] vssd1 vssd1 vccd1 vccd1 _00888_
+ sky130_fd_sc_hd__a22o_1
X_12833_ net286 _07616_ _07617_ net1849 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[173\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_35_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14069__A net1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18340_ _03828_ _03833_ _03835_ vssd1 vssd1 vccd1 vccd1 _03836_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_68_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15552_ ag2.body\[505\] net191 _01612_ ag2.body\[497\] vssd1 vssd1 vccd1 vccd1 _00827_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_56_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12764_ net237 _07585_ _07586_ net1754 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[135\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_57_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14503_ net1028 ag2.body\[181\] vssd1 vssd1 vccd1 vccd1 _08664_ sky130_fd_sc_hd__xor2_1
X_11715_ net566 _06683_ _06685_ _06686_ net469 vssd1 vssd1 vccd1 vccd1 _06687_ sky130_fd_sc_hd__a221o_1
X_18271_ net534 _03774_ vssd1 vssd1 vccd1 vccd1 _01383_ sky130_fd_sc_hd__and2_1
X_15483_ ag2.body\[571\] net109 _01605_ ag2.body\[563\] vssd1 vssd1 vccd1 vccd1 _00765_
+ sky130_fd_sc_hd__a22o_1
X_12695_ net259 net310 _07551_ _07552_ net1608 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[100\]
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_84_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17222_ _04103_ net887 net944 _04107_ vssd1 vssd1 vccd1 vccd1 _02901_ sky130_fd_sc_hd__a22o_1
XFILLER_0_83_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14434_ net1015 ag2.body\[22\] vssd1 vssd1 vccd1 vccd1 _08595_ sky130_fd_sc_hd__xnor2_1
X_11646_ net1124 _06618_ _06615_ _06485_ vssd1 vssd1 vccd1 vccd1 _06619_ sky130_fd_sc_hd__o211a_1
XANTENNA__11699__Y _06671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19798__CLK clknet_leaf_127_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16316__A1 net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14365_ net996 ag2.body\[600\] vssd1 vssd1 vccd1 vccd1 _08526_ sky130_fd_sc_hd__xor2_1
X_17153_ ag2.body\[611\] net715 net698 ag2.body\[614\] vssd1 vssd1 vccd1 vccd1 _02832_
+ sky130_fd_sc_hd__a22o_1
X_11577_ obsg2.obstacleArray\[81\] obsg2.obstacleArray\[85\] net514 vssd1 vssd1 vccd1
+ vccd1 _06550_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_103_clk clknet_4_10__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_103_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__17513__B1 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16104_ obsg2.obstacleArray\[66\] obsg2.obstacleArray\[67\] net426 vssd1 vssd1 vccd1
+ vccd1 _01783_ sky130_fd_sc_hd__mux2_1
XANTENNA__10061__B1 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13316_ net251 _07839_ _07840_ net1703 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[433\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11221__A net1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17084_ ag2.body\[192\] net737 net723 ag2.body\[194\] vssd1 vssd1 vccd1 vccd1 _02763_
+ sky130_fd_sc_hd__a22o_1
X_10528_ _05497_ _05498_ _05499_ _05500_ vssd1 vssd1 vccd1 vccd1 _05501_ sky130_fd_sc_hd__or4_1
XFILLER_0_68_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14296_ _08448_ _08451_ _08452_ _08456_ vssd1 vssd1 vccd1 vccd1 _08457_ sky130_fd_sc_hd__or4_1
Xhold809 control.body\[1010\] vssd1 vssd1 vccd1 vccd1 net2371 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16035_ net500 net462 net499 vssd1 vssd1 vccd1 vccd1 _01714_ sky130_fd_sc_hd__and3_1
X_13247_ net2068 net648 _07811_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[393\]
+ sky130_fd_sc_hd__and3_1
X_10459_ ag2.body\[448\] net1224 vssd1 vssd1 vccd1 vccd1 _05432_ sky130_fd_sc_hd__xor2_1
XFILLER_0_126_1186 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18004__A net46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_3698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16619__A2 net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13178_ _07780_ net253 _07778_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[355\]
+ sky130_fd_sc_hd__mux2_1
XANTENNA__10364__A1 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15827__B1 _01643_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10364__B2 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1304 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12129_ img_gen.tracker.frame\[570\] net549 net575 vssd1 vssd1 vccd1 vccd1 _07101_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_97_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19178__CLK clknet_leaf_53_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17986_ net46 _03604_ vssd1 vssd1 vccd1 vccd1 _03605_ sky130_fd_sc_hd__nor2_1
XFILLER_0_104_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15066__C net65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09506__B1 net1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13302__A1 net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11539__S1 net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19725_ clknet_leaf_133_clk _00669_ net1305 vssd1 vssd1 vccd1 vccd1 control.body\[667\]
+ sky130_fd_sc_hd__dfrtp_1
X_16937_ ag2.body\[526\] net943 vssd1 vssd1 vccd1 vccd1 _02616_ sky130_fd_sc_hd__xnor2_1
XANTENNA__17562__B net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16459__A _02057_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19656_ clknet_leaf_133_clk _00600_ net1309 vssd1 vssd1 vccd1 vccd1 control.body\[742\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09632__Y _04605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16868_ ag2.body\[467\] net850 vssd1 vssd1 vccd1 vccd1 _02547_ sky130_fd_sc_hd__or2_1
XANTENNA__10778__Y _05751_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18607_ clknet_leaf_17_clk img_gen.tracker.next_frame\[45\] net1318 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[45\] sky130_fd_sc_hd__dfrtp_1
X_15819_ ag2.body\[278\] net206 _01642_ ag2.body\[270\] vssd1 vssd1 vccd1 vccd1 _01064_
+ sky130_fd_sc_hd__a22o_1
X_19587_ clknet_leaf_118_clk _00531_ net1386 vssd1 vssd1 vccd1 vccd1 control.body\[801\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09809__A1 _04740_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16799_ _02476_ _02477_ net402 vssd1 vssd1 vccd1 vccd1 _02478_ sky130_fd_sc_hd__mux2_1
XANTENNA__14802__A1 net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14802__B2 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09340_ sound_gen.osc1.stayCount\[4\] _04343_ vssd1 vssd1 vccd1 vccd1 _04344_ sky130_fd_sc_hd__and2_1
X_18538_ clknet_leaf_135_clk _00064_ net1301 vssd1 vssd1 vccd1 vccd1 img_gen.updater.commands.count\[7\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_75_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10300__A net1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09271_ sound_gen.osc1.stayCount\[16\] sound_gen.osc1.stayCount\[14\] _04288_ vssd1
+ vssd1 vccd1 vccd1 _04294_ sky130_fd_sc_hd__a21o_1
XFILLER_0_30_1107 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18469_ net883 net871 net861 net851 vssd1 vssd1 vccd1 vccd1 _03955_ sky130_fd_sc_hd__a31o_1
XFILLER_0_75_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14707__A net975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20500_ clknet_leaf_22_clk _01387_ net1359 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[136\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_8_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20431_ clknet_leaf_23_clk _01318_ net1358 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[67\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__12041__A1 net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16307__A1 net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout122_A net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17504__B1 net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11131__A net1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12592__A2 net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20362_ clknet_leaf_21_clk _00002_ net1361 vssd1 vssd1 vccd1 vccd1 obsg2.obsNeeded\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_130_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17244__A2_N net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20293_ clknet_leaf_37_clk control.divider.next_count\[14\] net1349 vssd1 vssd1 vccd1
+ vccd1 control.divider.count\[14\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout1031_A ag2.randCord\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10970__A net1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14442__A net1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1129_A ag2.x\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout491_A net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout589_A net592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08986_ ag2.body\[80\] vssd1 vssd1 vccd1 vccd1 _04011_ sky130_fd_sc_hd__inv_2
XFILLER_0_23_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12897__A net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout377_X net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13844__A2 net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout756_A net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1498_A net1499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15273__A _04605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_1079 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09607_ net1146 control.body\[635\] vssd1 vssd1 vccd1 vccd1 _04580_ sky130_fd_sc_hd__xor2_1
XANTENNA__13505__B _07515_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout544_X net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09538_ net786 control.body\[1024\] _04505_ _04506_ _04508_ vssd1 vssd1 vccd1 vccd1
+ _04511_ sky130_fd_sc_hd__a2111o_1
XANTENNA__10210__A net1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout35_A net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16816__B net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_432 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09469_ _04135_ net1156 net1104 _04137_ _04441_ vssd1 vssd1 vccd1 vccd1 _04442_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout711_X net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1453_X net1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout809_X net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11500_ net1215 net1191 vssd1 vssd1 vccd1 vccd1 _06473_ sky130_fd_sc_hd__nor2_2
XFILLER_0_47_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12480_ net290 _07425_ _07430_ _07432_ net1617 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[5\]
+ sky130_fd_sc_hd__a32o_1
XANTENNA__10544__A_N net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_93_clk_X clknet_leaf_93_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11431_ _06400_ _06401_ _06402_ _06403_ vssd1 vssd1 vccd1 vccd1 _06404_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_134_4399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20629_ sound_gen.dac1.dacCount\[7\] vssd1 vssd1 vccd1 vccd1 net16 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_116_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14150_ net1006 ag2.body\[599\] vssd1 vssd1 vccd1 vccd1 _08311_ sky130_fd_sc_hd__xor2_1
X_11362_ net1148 control.body\[811\] vssd1 vssd1 vccd1 vccd1 _06335_ sky130_fd_sc_hd__xor2_1
XFILLER_0_22_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17647__B net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11791__B1 net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13101_ net243 _07742_ _07743_ net1965 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[315\]
+ sky130_fd_sc_hd__a22o_1
X_10313_ _05279_ _05284_ _05285_ vssd1 vssd1 vccd1 vccd1 _05286_ sky130_fd_sc_hd__or3_1
XFILLER_0_0_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14081_ net841 ag2.body\[560\] _04207_ net980 _08241_ vssd1 vssd1 vccd1 vccd1 _08242_
+ sky130_fd_sc_hd__a221o_1
X_11293_ _06260_ _06263_ _06264_ _06265_ vssd1 vssd1 vccd1 vccd1 _06266_ sky130_fd_sc_hd__or4_1
XANTENNA__14352__A net1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_957 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09736__B1 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13032_ net673 _07710_ vssd1 vssd1 vccd1 vccd1 _07711_ sky130_fd_sc_hd__nor2_1
X_10244_ _05213_ _05214_ _05215_ _05216_ _05207_ vssd1 vssd1 vccd1 vccd1 _05217_ sky130_fd_sc_hd__a221o_1
XANTENNA__09446__A net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11543__B1 net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1602 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15809__B1 _01641_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1101 net1106 vssd1 vssd1 vccd1 vccd1 net1101 sky130_fd_sc_hd__buf_4
XFILLER_0_24_1478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1112 ag2.x\[1\] vssd1 vssd1 vccd1 vccd1 net1112 sky130_fd_sc_hd__clkbuf_4
X_17840_ net790 net224 vssd1 vssd1 vccd1 vccd1 _03497_ sky130_fd_sc_hd__nor2_1
X_10175_ ag2.body\[417\] net1209 vssd1 vssd1 vccd1 vccd1 _05148_ sky130_fd_sc_hd__xor2_1
XANTENNA__20178__CLK clknet_leaf_88_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1123 net1129 vssd1 vssd1 vccd1 vccd1 net1123 sky130_fd_sc_hd__clkbuf_8
Xfanout1134 net1135 vssd1 vssd1 vccd1 vccd1 net1134 sky130_fd_sc_hd__clkbuf_4
Xfanout1145 net1156 vssd1 vssd1 vccd1 vccd1 net1145 sky130_fd_sc_hd__buf_2
Xfanout1156 ag2.y\[3\] vssd1 vssd1 vccd1 vccd1 net1156 sky130_fd_sc_hd__buf_4
XANTENNA__17382__B net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17771_ _03360_ _03365_ _03175_ vssd1 vssd1 vccd1 vccd1 _03450_ sky130_fd_sc_hd__o21a_1
Xfanout1167 net1173 vssd1 vssd1 vccd1 vccd1 net1167 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_101_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14983_ control.body\[1022\] net158 _01550_ control.body\[1014\] vssd1 vssd1 vccd1
+ vccd1 _00320_ sky130_fd_sc_hd__a22o_1
Xfanout180 net182 vssd1 vssd1 vccd1 vccd1 net180 sky130_fd_sc_hd__clkbuf_2
Xfanout1178 net1189 vssd1 vssd1 vccd1 vccd1 net1178 sky130_fd_sc_hd__buf_4
XFILLER_0_136_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout191 net192 vssd1 vssd1 vccd1 vccd1 net191 sky130_fd_sc_hd__clkbuf_2
X_19510_ clknet_leaf_113_clk _00454_ net1402 vssd1 vssd1 vccd1 vccd1 control.body\[884\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1189 ag2.y\[2\] vssd1 vssd1 vccd1 vccd1 net1189 sky130_fd_sc_hd__buf_4
X_16722_ obsg2.obstacleArray\[111\] net500 net481 obsg2.obstacleArray\[109\] _02400_
+ vssd1 vssd1 vccd1 vccd1 _02401_ sky130_fd_sc_hd__a221o_1
XANTENNA__09452__Y _04425_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13934_ ag2.body\[77\] net193 _08153_ ag2.body\[69\] vssd1 vssd1 vccd1 vccd1 _00158_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_92_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12600__A net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19441_ clknet_leaf_108_clk _00385_ net1421 vssd1 vssd1 vccd1 vccd1 control.body\[959\]
+ sky130_fd_sc_hd__dfrtp_1
X_16653_ net396 _02331_ _02330_ net360 vssd1 vssd1 vccd1 vccd1 _02332_ sky130_fd_sc_hd__a211o_1
X_13865_ _08030_ _08036_ vssd1 vssd1 vccd1 vccd1 _08139_ sky130_fd_sc_hd__nor2_1
XFILLER_0_53_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_104_3480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_104_3491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15604_ ag2.body\[470\] net121 _01619_ ag2.body\[462\] vssd1 vssd1 vccd1 vccd1 _00872_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11216__A net1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12816_ net286 _07608_ _07609_ net1635 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[164\]
+ sky130_fd_sc_hd__a22o_1
X_19372_ clknet_leaf_102_clk _00316_ net1426 vssd1 vssd1 vccd1 vccd1 control.body\[1018\]
+ sky130_fd_sc_hd__dfrtp_1
X_16584_ obsg2.obstacleArray\[66\] obsg2.obstacleArray\[67\] net446 vssd1 vssd1 vccd1
+ vccd1 _02263_ sky130_fd_sc_hd__mux2_1
XANTENNA__17322__A1_N net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13796_ img_gen.updater.commands.count\[15\] _08099_ vssd1 vssd1 vccd1 vccd1 _08102_
+ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_100_3366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18323_ _04947_ _08033_ vssd1 vssd1 vccd1 vccd1 _03819_ sky130_fd_sc_hd__nor2_1
XANTENNA__11074__A2 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_100_3377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15535_ ag2.body\[521\] net160 _01611_ ag2.body\[513\] vssd1 vssd1 vccd1 vccd1 _00811_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_100_3388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12747_ net258 _07576_ _07577_ net1779 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[127\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_57_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_1476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17734__B1 _02917_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10282__B1 _05253_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13431__A net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18254_ net353 _03633_ net37 obsg2.obstacleArray\[124\] vssd1 vssd1 vccd1 vccd1 _03766_
+ sky130_fd_sc_hd__a31o_1
X_12678_ net264 _07543_ _07544_ net1669 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[91\]
+ sky130_fd_sc_hd__a22o_1
X_15466_ ag2.body\[588\] net111 _01603_ ag2.body\[580\] vssd1 vssd1 vccd1 vccd1 _00750_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__10774__B net1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17205_ ag2.body\[176\] net738 _02878_ _02883_ vssd1 vssd1 vccd1 vccd1 _02884_ sky130_fd_sc_hd__a211o_1
XFILLER_0_53_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11629_ obsg2.obstacleArray\[32\] obsg2.obstacleArray\[36\] net510 vssd1 vssd1 vccd1
+ vccd1 _06602_ sky130_fd_sc_hd__mux2_1
X_14417_ net794 ag2.body\[535\] ag2.body\[528\] net844 vssd1 vssd1 vccd1 vccd1 _08578_
+ sky130_fd_sc_hd__a2bb2o_1
X_18185_ obsg2.obstacleArray\[89\] _03731_ net531 vssd1 vssd1 vccd1 vccd1 _01340_
+ sky130_fd_sc_hd__o21a_1
XANTENNA__17838__A net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_117_3885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15397_ control.body\[654\] net80 _01596_ net2356 vssd1 vssd1 vccd1 vccd1 _00688_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_117_3896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10034__B1 net1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17136_ _02811_ _02812_ _02813_ _02814_ vssd1 vssd1 vccd1 vccd1 _02815_ sky130_fd_sc_hd__a22o_1
XFILLER_0_128_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17557__B net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14348_ _08506_ _08507_ _08508_ vssd1 vssd1 vccd1 vccd1 _08509_ sky130_fd_sc_hd__or3_4
Xhold606 _00279_ vssd1 vssd1 vccd1 vccd1 net2168 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_1394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_1502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold617 control.body\[1055\] vssd1 vssd1 vccd1 vccd1 net2179 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10585__B2 _05557_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold628 control.divider.count\[10\] vssd1 vssd1 vccd1 vccd1 net2190 sky130_fd_sc_hd__dlygate4sd3_1
X_14279_ net994 ag2.body\[137\] vssd1 vssd1 vccd1 vccd1 _08440_ sky130_fd_sc_hd__xor2_1
XANTENNA__16170__C1 net347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17067_ ag2.body\[24\] net880 vssd1 vssd1 vccd1 vccd1 _02746_ sky130_fd_sc_hd__or2_1
Xhold639 control.body\[862\] vssd1 vssd1 vccd1 vccd1 net2201 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12334__X _07301_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xmax_cap358 _02227_ vssd1 vssd1 vccd1 vccd1 net358 sky130_fd_sc_hd__buf_4
XANTENNA__14262__A net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09727__B1 net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16018_ net860 _01696_ _01690_ vssd1 vssd1 vccd1 vccd1 _01697_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18568__CLK clknet_leaf_15_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19813__CLK clknet_leaf_124_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_1067 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17969_ _03590_ net45 vssd1 vssd1 vccd1 vccd1 _03593_ sky130_fd_sc_hd__nor2_1
XFILLER_0_58_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10014__B net1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15093__A _04553_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19708_ clknet_leaf_134_clk _00652_ net1307 vssd1 vssd1 vccd1 vccd1 control.body\[682\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_79_1490 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10949__B _05921_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19639_ clknet_leaf_123_clk _00583_ net1406 vssd1 vssd1 vccd1 vccd1 control.body\[757\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_0_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15821__A _04986_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19590__RESET_B net1386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09323_ sound_gen.dac1.dacCount\[2\] _04334_ vssd1 vssd1 vccd1 vccd1 _04335_ sky130_fd_sc_hd__and2_1
XANTENNA__14437__A net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10965__A net1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09254_ img_gen.updater.commands.rR1.rainbowRNG\[4\] vssd1 vssd1 vccd1 vccd1 _04279_
+ sky130_fd_sc_hd__inv_2
XANTENNA_fanout1079_A net1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_1274 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13060__B _07723_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09185_ ag2.body\[578\] vssd1 vssd1 vccd1 vccd1 _04210_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout504_A net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20424__RESET_B net1355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1246_A net1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20414_ clknet_leaf_32_clk _01301_ net1352 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[50\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__09818__X _04791_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17467__B net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11773__B1 net550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20345_ clknet_leaf_140_clk _01236_ net1293 vssd1 vssd1 vccd1 vccd1 img_gen.updater.commands.rR1.rainbowRNG\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15503__A2 net113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1034_X net1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1413_A net1414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20320__CLK clknet_leaf_43_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20276_ clknet_leaf_36_clk net1566 net1347 vssd1 vssd1 vccd1 vccd1 control.button2.Q\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10328__A1 _05283_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout494_X net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout873_A net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10328__B2 _05300_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19493__CLK clknet_leaf_113_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1201_X net1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_127_4192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08969_ ag2.body\[55\] vssd1 vssd1 vccd1 vccd1 _03994_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout759_X net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17008__A2 net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_123_4067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11980_ img_gen.tracker.frame\[547\] net541 net568 vssd1 vssd1 vccd1 vccd1 _06952_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_58_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_123_4089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_535 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19678__RESET_B net1386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10931_ net756 control.body\[1037\] _04252_ net1061 _05903_ vssd1 vssd1 vccd1 vccd1
+ _05904_ sky130_fd_sc_hd__o221a_1
XANTENNA__17930__B net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13235__B net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout926_X net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15731__A _05657_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13650_ control.divider.count\[16\] control.divider.count\[17\] _08004_ vssd1 vssd1
+ vccd1 vccd1 _08008_ sky130_fd_sc_hd__and3_1
X_10862_ _05826_ _05832_ _05833_ _05834_ vssd1 vssd1 vccd1 vccd1 _05835_ sky130_fd_sc_hd__or4_1
XFILLER_0_67_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout38_X net38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12601_ net328 _07501_ vssd1 vssd1 vccd1 vccd1 _07502_ sky130_fd_sc_hd__or2_1
XFILLER_0_67_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13581_ _03960_ control.divider.count\[7\] _07955_ vssd1 vssd1 vccd1 vccd1 _07956_
+ sky130_fd_sc_hd__a21o_1
X_10793_ ag2.body\[36\] net1128 vssd1 vssd1 vccd1 vccd1 _05766_ sky130_fd_sc_hd__nand2_1
XFILLER_0_112_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13251__A net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15320_ control.body\[712\] net73 _01589_ net2136 vssd1 vssd1 vccd1 vccd1 _00618_
+ sky130_fd_sc_hd__a22o_1
X_12532_ net606 net439 net469 net576 vssd1 vssd1 vccd1 vccd1 _07463_ sky130_fd_sc_hd__or4_1
XANTENNA__10264__B1 _04419_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_45_1689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_1502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15251_ control.body\[781\] net99 _01579_ net2171 vssd1 vssd1 vccd1 vccd1 _00559_
+ sky130_fd_sc_hd__a22o_1
X_12463_ net1621 _07420_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[0\] sky130_fd_sc_hd__and2_1
XFILLER_0_48_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_10_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20165__RESET_B net1484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14202_ _08361_ _08362_ vssd1 vssd1 vccd1 vccd1 _08363_ sky130_fd_sc_hd__nand2b_1
X_11414_ net1100 control.body\[853\] vssd1 vssd1 vccd1 vccd1 _06387_ sky130_fd_sc_hd__nand2_1
XFILLER_0_69_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15182_ _04494_ net53 vssd1 vssd1 vccd1 vccd1 _01572_ sky130_fd_sc_hd__nor2_2
XANTENNA__14950__B1 _01546_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12394_ img_gen.updater.commands.rR1.rainbowRNG\[10\] _07319_ _07338_ _07350_ _07358_
+ vssd1 vssd1 vccd1 vccd1 _07359_ sky130_fd_sc_hd__a221o_1
XANTENNA_clkbuf_leaf_73_clk_A clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14133_ net1009 ag2.body\[175\] vssd1 vssd1 vccd1 vccd1 _08294_ sky130_fd_sc_hd__or2_1
XFILLER_0_1_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_570 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11345_ ag2.body\[444\] net1127 vssd1 vssd1 vccd1 vccd1 _06318_ sky130_fd_sc_hd__xor2_1
XANTENNA__17945__X _03574_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09447__Y _04420_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19990_ clknet_leaf_64_clk _00934_ net1474 vssd1 vssd1 vccd1 vccd1 ag2.body\[404\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__16152__C1 net349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_3089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14064_ _08220_ _08223_ _08224_ vssd1 vssd1 vccd1 vccd1 _08225_ sky130_fd_sc_hd__or3_2
X_18941_ clknet_leaf_139_clk img_gen.tracker.next_frame\[379\] net1288 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[379\] sky130_fd_sc_hd__dfrtp_1
X_11276_ ag2.body\[120\] net1235 vssd1 vssd1 vccd1 vccd1 _06249_ sky130_fd_sc_hd__xor2_1
XANTENNA__11516__B1 _06485_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13015_ net668 _07702_ vssd1 vssd1 vccd1 vccd1 _07703_ sky130_fd_sc_hd__nor2_1
X_10227_ ag2.body\[561\] net1203 vssd1 vssd1 vccd1 vccd1 _05200_ sky130_fd_sc_hd__xor2_1
XANTENNA__17247__A2 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_88_clk_A clknet_4_12__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18872_ clknet_leaf_22_clk img_gen.tracker.next_frame\[310\] net1342 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[310\] sky130_fd_sc_hd__dfrtp_1
X_17823_ ag2.body\[7\] _03474_ _03476_ _03488_ vssd1 vssd1 vccd1 vccd1 _01222_ sky130_fd_sc_hd__a22o_1
X_10158_ ag2.body\[60\] net760 net744 ag2.body\[63\] _05123_ vssd1 vssd1 vccd1 vccd1
+ _05131_ sky130_fd_sc_hd__a221o_1
XANTENNA_clkbuf_leaf_131_clk_A clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold3 control.button3.Q\[1\] vssd1 vssd1 vccd1 vccd1 net1565 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11645__S net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_3542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17754_ _03428_ _03429_ _03430_ _03432_ vssd1 vssd1 vccd1 vccd1 _03433_ sky130_fd_sc_hd__and4_1
XFILLER_0_101_1498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14334__A1_N net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_3553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10089_ net758 control.body\[796\] control.body\[797\] net753 vssd1 vssd1 vccd1 vccd1
+ _05062_ sky130_fd_sc_hd__o22ai_1
X_14966_ control.body\[1024\] net157 net51 control.body\[1016\] vssd1 vssd1 vccd1
+ vccd1 _00306_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_106_3564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_11_clk_A clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20320__Q obsg2.randCord\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10769__B net1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16705_ _02378_ _02383_ net433 vssd1 vssd1 vccd1 vccd1 _02384_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_102_3428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13917_ ag2.body\[62\] net129 _08151_ ag2.body\[54\] vssd1 vssd1 vccd1 vccd1 _00143_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12687__D _07306_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17685_ _04168_ net869 net723 ag2.body\[474\] _03363_ vssd1 vssd1 vccd1 vccd1 _03364_
+ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_102_3439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14897_ control.body\[1090\] net178 _01540_ net2485 vssd1 vssd1 vccd1 vccd1 _00244_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_58_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19424_ clknet_leaf_111_clk _00368_ net1430 vssd1 vssd1 vccd1 vccd1 control.body\[974\]
+ sky130_fd_sc_hd__dfrtp_1
X_16636_ obsg2.obstacleArray\[56\] obsg2.obstacleArray\[57\] net445 vssd1 vssd1 vccd1
+ vccd1 _02315_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_146_clk_A clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13848_ ag2.body\[12\] net117 _08133_ net927 vssd1 vssd1 vccd1 vccd1 _00092_ sky130_fd_sc_hd__a22o_1
XFILLER_0_58_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19355_ clknet_leaf_101_clk _00299_ net1438 vssd1 vssd1 vccd1 vccd1 control.body\[1033\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_130_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16567_ obsg2.obstacleArray\[123\] net449 net390 _02245_ vssd1 vssd1 vccd1 vccd1
+ _02246_ sky130_fd_sc_hd__o211a_1
XANTENNA_clkbuf_leaf_26_clk_A clknet_4_4__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10785__A net1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_2760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13779_ _08088_ _08089_ vssd1 vssd1 vccd1 vccd1 _00067_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_80_2771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_119_3947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18306_ _03801_ vssd1 vssd1 vccd1 vccd1 _03802_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_119_3958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19366__CLK clknet_leaf_102_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15518_ ag2.body\[538\] net156 _01609_ ag2.body\[530\] vssd1 vssd1 vccd1 vccd1 _00796_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_61_2170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19286_ clknet_leaf_98_clk _00230_ net1447 vssd1 vssd1 vccd1 vccd1 control.body\[1108\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_61_2181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16498_ obsg2.obstacleArray\[16\] obsg2.obstacleArray\[17\] obsg2.obstacleArray\[18\]
+ obsg2.obstacleArray\[19\] net458 net399 vssd1 vssd1 vccd1 vccd1 _02177_ sky130_fd_sc_hd__mux4_1
XFILLER_0_84_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_1583 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_2192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18237_ net519 _03757_ vssd1 vssd1 vccd1 vccd1 _01366_ sky130_fd_sc_hd__nor2_1
XANTENNA__15194__B1 _01573_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15449_ ag2.body\[605\] net86 _01601_ ag2.body\[597\] vssd1 vssd1 vccd1 vccd1 _00735_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__15733__A2 net200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14544__X _08705_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18168_ _03604_ net36 vssd1 vssd1 vccd1 vccd1 _03723_ sky130_fd_sc_hd__nor2_1
XFILLER_0_128_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18278__A4 _03577_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09412__A2 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10009__B _04239_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold403 img_gen.tracker.frame\[315\] vssd1 vssd1 vccd1 vccd1 net1965 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_128_1078 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold414 img_gen.tracker.frame\[416\] vssd1 vssd1 vccd1 vccd1 net1976 sky130_fd_sc_hd__dlygate4sd3_1
X_17119_ ag2.body\[541\] net952 vssd1 vssd1 vccd1 vccd1 _02798_ sky130_fd_sc_hd__xor2_1
XANTENNA__17486__A2 net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold425 img_gen.tracker.frame\[337\] vssd1 vssd1 vccd1 vccd1 net1987 sky130_fd_sc_hd__dlygate4sd3_1
X_18099_ net44 _03681_ vssd1 vssd1 vccd1 vccd1 _03682_ sky130_fd_sc_hd__nor2_1
Xhold436 img_gen.tracker.frame\[111\] vssd1 vssd1 vccd1 vccd1 net1998 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12505__A net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold447 img_gen.tracker.frame\[438\] vssd1 vssd1 vccd1 vccd1 net2009 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold458 img_gen.tracker.frame\[462\] vssd1 vssd1 vccd1 vccd1 net2020 sky130_fd_sc_hd__dlygate4sd3_1
X_20130_ clknet_leaf_81_clk _01074_ net1449 vssd1 vssd1 vccd1 vccd1 ag2.body\[256\]
+ sky130_fd_sc_hd__dfrtp_4
X_09941_ _03984_ net1197 net754 ag2.body\[29\] _04913_ vssd1 vssd1 vccd1 vccd1 _04914_
+ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_74_2586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold469 img_gen.tracker.frame\[440\] vssd1 vssd1 vccd1 vccd1 net2031 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_96_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__20493__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout905 net908 vssd1 vssd1 vccd1 vccd1 net905 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_106_1387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout916 control.body_update.curr_length\[2\] vssd1 vssd1 vccd1 vccd1 net916 sky130_fd_sc_hd__buf_2
Xfanout927 ag2.body\[4\] vssd1 vssd1 vccd1 vccd1 net927 sky130_fd_sc_hd__clkbuf_4
X_20061_ clknet_leaf_72_clk _01005_ net1502 vssd1 vssd1 vccd1 vccd1 ag2.body\[331\]
+ sky130_fd_sc_hd__dfrtp_4
X_09872_ _04833_ _04834_ _04839_ _04844_ vssd1 vssd1 vccd1 vccd1 _04845_ sky130_fd_sc_hd__or4_2
XFILLER_0_110_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout938 net941 vssd1 vssd1 vccd1 vccd1 net938 sky130_fd_sc_hd__clkbuf_4
Xfanout949 net950 vssd1 vssd1 vccd1 vccd1 net949 sky130_fd_sc_hd__buf_4
XANTENNA__16446__B1 net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09814__A net1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout287_A net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09479__A2 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18199__B1 net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_2969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10679__B net1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20230__Q ag2.body\[164\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout454_A net459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_92_clk clknet_4_9__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_92_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_95_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1196_A net1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10494__B1 net1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_1494 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout621_A net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout242_X net242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout719_A net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09306_ _04325_ vssd1 vssd1 vccd1 vccd1 _04326_ sky130_fd_sc_hd__inv_2
XANTENNA__13071__A _07558_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14195__A2_N ag2.body\[167\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_135_4450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11994__B1 net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_4314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09237_ net883 vssd1 vssd1 vccd1 vccd1 _04262_ sky130_fd_sc_hd__inv_2
XFILLER_0_8_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_131_4325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16382__A net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1151_X net1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_1531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout507_X net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_1542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09939__B1 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09168_ ag2.body\[529\] vssd1 vssd1 vccd1 vccd1 _04193_ sky130_fd_sc_hd__inv_2
XANTENNA__17197__B net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout990_A net995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18123__B1 net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14614__B ag2.body\[58\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17477__A2 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17765__X _03444_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09099_ ag2.body\[350\] vssd1 vssd1 vccd1 vccd1 _04124_ sky130_fd_sc_hd__inv_2
X_11130_ net1099 control.body\[869\] vssd1 vssd1 vccd1 vccd1 _06103_ sky130_fd_sc_hd__nand2_1
X_20328_ clknet_leaf_105_clk sound_gen.osc1.timer_nxt\[14\] _00005_ vssd1 vssd1 vccd1
+ vccd1 sound_gen.osc1.timer\[2\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_129_4243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_129_4254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold970 _00509_ vssd1 vssd1 vccd1 vccd1 net2532 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_4265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout876_X net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold981 control.body\[792\] vssd1 vssd1 vccd1 vccd1 net2543 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14160__A1 net996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11061_ ag2.body\[439\] net1069 vssd1 vssd1 vccd1 vccd1 _06034_ sky130_fd_sc_hd__xnor2_1
Xhold992 control.body\[1030\] vssd1 vssd1 vccd1 vccd1 net2554 sky130_fd_sc_hd__dlygate4sd3_1
X_20259_ clknet_leaf_45_clk _01203_ net1379 vssd1 vssd1 vccd1 vccd1 ag2.body\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_38_1482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_1464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14160__B2 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_125_4129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18102__A net44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_1493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10012_ net903 _04979_ _04417_ vssd1 vssd1 vccd1 vccd1 _04985_ sky130_fd_sc_hd__a21o_2
XTAP_TAPCELL_ROW_34_1357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09724__A net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19239__CLK clknet_leaf_83_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14820_ net809 ag2.body\[157\] ag2.body\[152\] net845 vssd1 vssd1 vccd1 vccd1 _01491_
+ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__17941__A net48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13246__A net384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09443__B net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17660__B net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14751_ net837 ag2.body\[105\] ag2.body\[111\] net794 _08906_ vssd1 vssd1 vccd1 vccd1
+ _08912_ sky130_fd_sc_hd__a221o_1
XFILLER_0_25_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11963_ img_gen.tracker.frame\[493\] net617 net571 _06934_ vssd1 vssd1 vccd1 vccd1
+ _06935_ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_83_clk clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_83_clk
+ sky130_fd_sc_hd__clkbuf_8
X_13702_ track.highScore\[3\] _04642_ _08038_ _08041_ _08042_ vssd1 vssd1 vccd1 vccd1
+ _08043_ sky130_fd_sc_hd__o221ai_1
XANTENNA__10485__B1 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10914_ ag2.body\[459\] net1153 vssd1 vssd1 vccd1 vccd1 _05887_ sky130_fd_sc_hd__xnor2_1
X_17470_ _04194_ net863 net942 _04196_ vssd1 vssd1 vccd1 vccd1 _03149_ sky130_fd_sc_hd__o22a_1
XFILLER_0_131_1403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14682_ net1039 ag2.body\[92\] vssd1 vssd1 vccd1 vccd1 _08843_ sky130_fd_sc_hd__xnor2_1
X_11894_ _06864_ _06865_ net564 vssd1 vssd1 vccd1 vccd1 _06866_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16421_ _02096_ _02098_ _02099_ net364 vssd1 vssd1 vccd1 vccd1 _02100_ sky130_fd_sc_hd__a22o_1
XFILLER_0_67_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13633_ _07995_ _07996_ net222 vssd1 vssd1 vccd1 vccd1 control.divider.next_count\[11\]
+ sky130_fd_sc_hd__and3b_1
X_10845_ net758 ag2.body\[44\] _03988_ net1169 vssd1 vssd1 vccd1 vccd1 _05818_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_132_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__20346__RESET_B net1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14077__A net1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__20366__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19140_ clknet_leaf_139_clk net8 net1289 vssd1 vssd1 vccd1 vccd1 img_gen.control.button5.Q\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_16352_ obsg2.obstacleArray\[6\] net409 vssd1 vssd1 vccd1 vccd1 _02031_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_15_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12777__A2 net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13564_ _07931_ _07942_ ssdec1.in\[2\] vssd1 vssd1 vccd1 vccd1 _07943_ sky130_fd_sc_hd__mux2_1
X_10776_ ag2.body\[217\] net1210 vssd1 vssd1 vccd1 vccd1 _05749_ sky130_fd_sc_hd__xor2_1
XFILLER_0_32_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15303_ control.body\[730\] net77 _01586_ net2432 vssd1 vssd1 vccd1 vccd1 _00604_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_97_3276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19071_ clknet_leaf_29_clk img_gen.tracker.next_frame\[509\] net1336 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[509\] sky130_fd_sc_hd__dfrtp_1
X_12515_ net315 _07454_ vssd1 vssd1 vccd1 vccd1 _07455_ sky130_fd_sc_hd__or2_1
XFILLER_0_125_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16283_ _01960_ _01961_ net419 vssd1 vssd1 vccd1 vccd1 _01962_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_114_3800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_3287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13495_ net328 _07508_ _07813_ vssd1 vssd1 vccd1 vccd1 _07910_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_114_3811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18022_ net299 _03630_ vssd1 vssd1 vccd1 vccd1 _03631_ sky130_fd_sc_hd__nand2_1
XFILLER_0_129_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15234_ control.body\[798\] net96 _01577_ net2297 vssd1 vssd1 vccd1 vccd1 _00544_
+ sky130_fd_sc_hd__a22o_1
X_12446_ _07354_ _07388_ _07398_ _07406_ vssd1 vssd1 vccd1 vccd1 _07407_ sky130_fd_sc_hd__a31o_1
XANTENNA__14923__B1 _01543_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11737__B1 net553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11500__Y _06473_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17468__A2 net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15165_ control.body\[848\] net103 _01570_ net2495 vssd1 vssd1 vccd1 vccd1 _00482_
+ sky130_fd_sc_hd__a22o_1
X_12377_ img_gen.updater.commands.count\[7\] img_gen.updater.commands.count\[6\] img_gen.updater.commands.count\[5\]
+ vssd1 vssd1 vccd1 vccd1 _07342_ sky130_fd_sc_hd__and3_1
XFILLER_0_50_652 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16676__B1 net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11328_ net1168 control.body\[658\] vssd1 vssd1 vccd1 vccd1 _06301_ sky130_fd_sc_hd__xor2_1
XFILLER_0_65_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14116_ _08269_ _08270_ _08271_ _08272_ _08276_ vssd1 vssd1 vccd1 vccd1 _08277_ sky130_fd_sc_hd__a221o_1
X_19973_ clknet_leaf_63_clk _00917_ net1470 vssd1 vssd1 vccd1 vccd1 ag2.body\[419\]
+ sky130_fd_sc_hd__dfrtp_4
X_15096_ net2622 net145 _01563_ net2164 vssd1 vssd1 vccd1 vccd1 _00420_ sky130_fd_sc_hd__a22o_1
XFILLER_0_120_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18924_ clknet_leaf_140_clk img_gen.tracker.next_frame\[362\] net1291 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[362\] sky130_fd_sc_hd__dfrtp_1
X_14047_ net988 ag2.body\[185\] vssd1 vssd1 vccd1 vccd1 _08208_ sky130_fd_sc_hd__xnor2_1
X_11259_ _06227_ _06228_ _06231_ _04491_ vssd1 vssd1 vccd1 vccd1 _06232_ sky130_fd_sc_hd__a211o_1
XFILLER_0_43_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14151__B2 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14540__A net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_3604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_3615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12162__B1 net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_3626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18855_ clknet_leaf_18_clk img_gen.tracker.next_frame\[293\] net1323 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[293\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__10712__A1 net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17806_ _03474_ vssd1 vssd1 vccd1 vccd1 _03475_ sky130_fd_sc_hd__inv_2
XFILLER_0_94_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19529__RESET_B net1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18606__CLK clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18786_ clknet_leaf_13_clk img_gen.tracker.next_frame\[224\] net1284 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[224\] sky130_fd_sc_hd__dfrtp_1
X_15998_ net690 _01676_ vssd1 vssd1 vccd1 vccd1 _01677_ sky130_fd_sc_hd__nor2_1
XFILLER_0_89_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17737_ _03304_ _03309_ _03323_ vssd1 vssd1 vccd1 vccd1 _03416_ sky130_fd_sc_hd__o21a_1
XANTENNA__17570__B net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_1471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14949_ control.body\[1040\] net172 _01546_ net2260 vssd1 vssd1 vccd1 vccd1 _00290_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12465__A1 net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_74_clk clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_74_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_82_2811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_82_2822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10476__B1 _05435_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_2833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_527 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17668_ ag2.body\[450\] net861 vssd1 vssd1 vccd1 vccd1 _03347_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_63_2232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_2243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19407_ clknet_leaf_103_clk _00351_ net1431 vssd1 vssd1 vccd1 vccd1 control.body\[989\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_114_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16619_ obsg2.obstacleArray\[47\] net449 net390 vssd1 vssd1 vccd1 vccd1 _02298_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_63_2254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18756__CLK clknet_leaf_15_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17599_ ag2.body\[422\] net697 vssd1 vssd1 vccd1 vccd1 _03278_ sky130_fd_sc_hd__nor2_1
XANTENNA__20087__RESET_B net1492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19338_ clknet_leaf_100_clk net2407 net1443 vssd1 vssd1 vccd1 vccd1 control.body\[1048\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_46_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09633__A2 _04599_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11976__B1 net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10779__B2 _05739_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16914__B net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19269_ clknet_leaf_71_clk _00213_ net1503 vssd1 vssd1 vccd1 vccd1 ag2.body\[132\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_31_1098 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_323 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09022_ ag2.body\[156\] vssd1 vssd1 vccd1 vccd1 _04047_ sky130_fd_sc_hd__inv_2
XFILLER_0_66_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_76_2626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_76_2637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16852__A2_N net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_2648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14390__A1 net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold200 img_gen.tracker.frame\[451\] vssd1 vssd1 vccd1 vccd1 net1762 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_2047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17459__A2 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold211 img_gen.tracker.frame\[84\] vssd1 vssd1 vccd1 vccd1 net1773 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14390__B2 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_2058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_2069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold222 img_gen.tracker.frame\[333\] vssd1 vssd1 vccd1 vccd1 net1784 sky130_fd_sc_hd__dlygate4sd3_1
Xhold233 img_gen.tracker.frame\[163\] vssd1 vssd1 vccd1 vccd1 net1795 sky130_fd_sc_hd__dlygate4sd3_1
Xhold244 img_gen.tracker.frame\[456\] vssd1 vssd1 vccd1 vccd1 net1806 sky130_fd_sc_hd__dlygate4sd3_1
Xhold255 img_gen.tracker.frame\[160\] vssd1 vssd1 vccd1 vccd1 net1817 sky130_fd_sc_hd__dlygate4sd3_1
Xhold266 img_gen.tracker.frame\[532\] vssd1 vssd1 vccd1 vccd1 net1828 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold277 img_gen.tracker.frame\[437\] vssd1 vssd1 vccd1 vccd1 net1839 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14142__A1 net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20113_ clknet_leaf_79_clk _01057_ net1488 vssd1 vssd1 vccd1 vccd1 ag2.body\[287\]
+ sky130_fd_sc_hd__dfrtp_4
Xhold288 img_gen.tracker.frame\[44\] vssd1 vssd1 vccd1 vccd1 net1850 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14142__B2 net1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout702 _04268_ vssd1 vssd1 vccd1 vccd1 net702 sky130_fd_sc_hd__clkbuf_4
X_09924_ _04433_ _04640_ vssd1 vssd1 vccd1 vccd1 _04897_ sky130_fd_sc_hd__nor2_2
Xhold299 img_gen.tracker.frame\[297\] vssd1 vssd1 vccd1 vccd1 net1861 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout713 net714 vssd1 vssd1 vccd1 vccd1 net713 sky130_fd_sc_hd__buf_4
XANTENNA__16141__S net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout724 net725 vssd1 vssd1 vccd1 vccd1 net724 sky130_fd_sc_hd__buf_4
XFILLER_0_0_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1111_A net1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16419__B1 net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1209_A net1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout735 _04263_ vssd1 vssd1 vccd1 vccd1 net735 sky130_fd_sc_hd__buf_4
XANTENNA__15890__A1 ag2.body\[214\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout746 net747 vssd1 vssd1 vccd1 vccd1 net746 sky130_fd_sc_hd__buf_4
X_20044_ clknet_leaf_68_clk _00988_ net1498 vssd1 vssd1 vccd1 vccd1 ag2.body\[346\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA_input7_A gpio_in[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout757 _04232_ vssd1 vssd1 vccd1 vccd1 net757 sky130_fd_sc_hd__clkbuf_8
X_09855_ net1110 _04250_ control.body\[975\] net745 _04827_ vssd1 vssd1 vccd1 vccd1
+ _04828_ sky130_fd_sc_hd__o221a_1
XANTENNA_fanout192_X net192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout571_A net573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout768 _04230_ vssd1 vssd1 vccd1 vccd1 net768 sky130_fd_sc_hd__clkbuf_8
Xfanout779 net781 vssd1 vssd1 vccd1 vccd1 net779 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11900__B1 net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout669_A net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13066__A net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09786_ net890 _04758_ vssd1 vssd1 vccd1 vccd1 _04759_ sky130_fd_sc_hd__nor2_2
XANTENNA__19531__CLK clknet_leaf_118_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_1545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_134_Right_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17480__B net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1480_A net1484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_65_clk clknet_4_13__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_65_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout836_A _03965_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1199_X net1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_4_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_137_4501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_137_4512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1100 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_46_1740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout624_X net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15945__A2 net195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10219__B1 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10630_ net1194 control.body\[665\] vssd1 vssd1 vccd1 vccd1 _05603_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_27_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16824__B net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14809__A1_N net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_23_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_23_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10561_ ag2.body\[512\] net1228 vssd1 vssd1 vccd1 vccd1 _05534_ sky130_fd_sc_hd__and2b_1
XANTENNA__16355__C1 net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18834__RESET_B net1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14625__A net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12300_ _07202_ _07210_ vssd1 vssd1 vccd1 vccd1 _07267_ sky130_fd_sc_hd__and2b_1
XFILLER_0_122_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13280_ net234 _07825_ _07826_ net1820 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[411\]
+ sky130_fd_sc_hd__a22o_1
X_10492_ ag2.body\[547\] net1158 vssd1 vssd1 vccd1 vccd1 _05465_ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout993_X net993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19196__Q ag2.body\[59\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10872__B net1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_92_3140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11719__B1 net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12231_ _07188_ _07200_ vssd1 vssd1 vccd1 vccd1 _07201_ sky130_fd_sc_hd__or2_1
XANTENNA__13184__A2 net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09438__B net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09927__A3 _04897_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16658__B1 net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12162_ img_gen.tracker.frame\[405\] net584 net568 vssd1 vssd1 vccd1 vccd1 _07134_
+ sky130_fd_sc_hd__o21a_1
XANTENNA__17655__B net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11680__A_N net1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_1419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11113_ net775 control.body\[1098\] control.body\[1102\] net751 vssd1 vssd1 vccd1
+ vccd1 _06086_ sky130_fd_sc_hd__o2bb2a_1
X_16970_ ag2.body\[411\] net718 net691 ag2.body\[415\] vssd1 vssd1 vccd1 vccd1 _02649_
+ sky130_fd_sc_hd__o22a_1
X_12093_ _06661_ _07058_ _07064_ _07052_ net436 vssd1 vssd1 vccd1 vccd1 _07065_ sky130_fd_sc_hd__o311a_1
XANTENNA__18629__CLK clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12144__B1 net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15921_ ag2.body\[176\] net136 _01654_ ag2.body\[168\] vssd1 vssd1 vccd1 vccd1 _01154_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__15881__B2 ag2.body\[214\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11044_ _05963_ _06016_ _05985_ _05973_ vssd1 vssd1 vccd1 vccd1 _06017_ sky130_fd_sc_hd__or4b_2
XANTENNA__12695__A1 net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18640_ clknet_leaf_15_clk img_gen.tracker.next_frame\[78\] net1312 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[78\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__17622__A2 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15852_ ag2.body\[244\] net176 _01645_ ag2.body\[236\] vssd1 vssd1 vccd1 vccd1 _01094_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_137_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14803_ net844 ag2.body\[288\] ag2.body\[295\] net795 vssd1 vssd1 vccd1 vccd1 _01474_
+ sky130_fd_sc_hd__a22oi_1
XANTENNA__16830__B1 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18571_ clknet_leaf_15_clk img_gen.tracker.next_frame\[9\] net1313 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[9\] sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_101_Right_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15783_ ag2.body\[310\] net208 _01638_ ag2.body\[302\] vssd1 vssd1 vccd1 vccd1 _01032_
+ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_56_clk clknet_4_12__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_56_clk
+ sky130_fd_sc_hd__clkbuf_8
X_12995_ _07693_ net254 _07691_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[259\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17522_ _03197_ _03198_ _03199_ _03200_ vssd1 vssd1 vccd1 vccd1 _03201_ sky130_fd_sc_hd__or4_1
X_14734_ _08892_ _08893_ _08894_ _08891_ vssd1 vssd1 vccd1 vccd1 _08895_ sky130_fd_sc_hd__a211o_1
XANTENNA__09901__B net1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11946_ img_gen.tracker.frame\[121\] net618 vssd1 vssd1 vccd1 vccd1 _06918_ sky130_fd_sc_hd__or2_1
XFILLER_0_52_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17453_ ag2.body\[438\] net940 vssd1 vssd1 vccd1 vccd1 _03132_ sky130_fd_sc_hd__xnor2_1
X_14665_ net1038 ag2.body\[524\] vssd1 vssd1 vccd1 vccd1 _08826_ sky130_fd_sc_hd__xor2_1
XANTENNA__15936__A2 net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_99_3338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11670__A2 net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11877_ _06846_ _06848_ net570 vssd1 vssd1 vccd1 vccd1 _06849_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_99_3349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16404_ _02079_ _02082_ net364 vssd1 vssd1 vccd1 vccd1 _02083_ sky130_fd_sc_hd__mux2_1
XANTENNA__11224__A net1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13616_ control.divider.count\[5\] _07959_ net220 vssd1 vssd1 vccd1 vccd1 _07986_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_39_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10828_ ag2.body\[311\] net1067 vssd1 vssd1 vccd1 vccd1 _05801_ sky130_fd_sc_hd__xor2_1
X_17384_ ag2.body\[494\] net942 vssd1 vssd1 vccd1 vccd1 _03063_ sky130_fd_sc_hd__or2_1
X_14596_ net978 ag2.body\[307\] vssd1 vssd1 vccd1 vccd1 _08757_ sky130_fd_sc_hd__xor2_1
XFILLER_0_116_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19123_ clknet_leaf_141_clk img_gen.tracker.next_frame\[561\] net1294 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[561\] sky130_fd_sc_hd__dfrtp_1
X_16335_ obsg2.obstacleArray\[87\] net414 _02013_ net416 vssd1 vssd1 vccd1 vccd1 _02014_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_109_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13547_ net226 _07929_ vssd1 vssd1 vccd1 vccd1 _07930_ sky130_fd_sc_hd__nor2_1
XFILLER_0_137_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10759_ _05728_ _05729_ _05730_ _05731_ vssd1 vssd1 vccd1 vccd1 _05732_ sky130_fd_sc_hd__a22o_1
XANTENNA__12607__X _07505_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16897__B1 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19054_ clknet_leaf_8_clk img_gen.tracker.next_frame\[492\] net1272 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[492\] sky130_fd_sc_hd__dfrtp_1
X_16266_ net417 _01942_ _01944_ net369 vssd1 vssd1 vccd1 vccd1 _01945_ sky130_fd_sc_hd__a211o_1
X_13478_ net250 _07902_ _07903_ net1828 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[532\]
+ sky130_fd_sc_hd__a22o_1
X_18005_ obsg2.obstacleArray\[22\] _03618_ net533 vssd1 vssd1 vccd1 vccd1 _01273_
+ sky130_fd_sc_hd__o21a_1
X_15217_ control.body\[815\] net92 _01575_ net2208 vssd1 vssd1 vccd1 vccd1 _00529_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__19404__CLK clknet_leaf_103_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12429_ _06629_ _07390_ _06627_ vssd1 vssd1 vccd1 vccd1 _07391_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_125_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16197_ obsg2.obstacleArray\[62\] obsg2.obstacleArray\[63\] net424 vssd1 vssd1 vccd1
+ vccd1 _01876_ sky130_fd_sc_hd__mux2_1
XFILLER_0_124_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_1615 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_71_2501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15148_ net2311 net105 _01568_ control.body\[857\] vssd1 vssd1 vccd1 vccd1 _00467_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_26_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10933__A1 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10933__B2 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1069 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19956_ clknet_leaf_44_clk _00900_ net1381 vssd1 vssd1 vccd1 vccd1 ag2.body\[434\]
+ sky130_fd_sc_hd__dfrtp_4
X_15079_ net2597 net151 _01561_ net2242 vssd1 vssd1 vccd1 vccd1 _00405_ sky130_fd_sc_hd__a22o_1
XANTENNA__12135__B1 net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18907_ clknet_leaf_144_clk img_gen.tracker.next_frame\[345\] net1251 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[345\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__12686__A1 net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19887_ clknet_leaf_86_clk _00831_ net1460 vssd1 vssd1 vccd1 vccd1 ag2.body\[509\]
+ sky130_fd_sc_hd__dfrtp_4
Xclkbuf_4_0__f_clk clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_0__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_09640_ _04608_ _04610_ _04611_ _04612_ vssd1 vssd1 vccd1 vccd1 _04613_ sky130_fd_sc_hd__or4b_1
XANTENNA__10922__A2_N net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10303__A net1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18838_ clknet_leaf_4_clk img_gen.tracker.next_frame\[276\] net1277 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[276\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_69_2430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_69_2441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09571_ ag2.body\[204\] net763 net757 ag2.body\[205\] vssd1 vssd1 vccd1 vccd1 _04544_
+ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_65_2305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18769_ clknet_leaf_18_clk img_gen.tracker.next_frame\[207\] net1321 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[207\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_116_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_65_2316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_47_clk clknet_4_7__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_47_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__11646__C1 _06485_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10957__B net1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout152_A net154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11134__A net1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17535__A2_N net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12205__A4 _07147_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11949__B1 net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_1651 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16337__C1 net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12610__A1 net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20593_ net1525 vssd1 vssd1 vccd1 vccd1 gpio_oeb[5] sky130_fd_sc_hd__buf_2
XANTENNA__10973__A net1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_2109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1061_A net1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14445__A net1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16888__B1 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1159_A net1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09005_ ag2.body\[122\] vssd1 vssd1 vccd1 vccd1 _04030_ sky130_fd_sc_hd__inv_2
XFILLER_0_5_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_1268 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17475__B net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout786_A net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14115__A1 net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14115__B2 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_1435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout510 net515 vssd1 vssd1 vccd1 vccd1 net510 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout1114_X net1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12126__B1 net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1508 net9 vssd1 vssd1 vccd1 vccd1 net1508 sky130_fd_sc_hd__buf_2
Xfanout521 net528 vssd1 vssd1 vccd1 vccd1 net521 sky130_fd_sc_hd__buf_2
Xfanout532 net533 vssd1 vssd1 vccd1 vccd1 net532 sky130_fd_sc_hd__clkbuf_2
X_09907_ ag2.body\[132\] net1141 vssd1 vssd1 vccd1 vccd1 _04880_ sky130_fd_sc_hd__nand2_1
Xfanout543 net553 vssd1 vssd1 vccd1 vccd1 net543 sky130_fd_sc_hd__clkbuf_2
XANTENNA__12677__A1 net241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout953_A net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout554 net555 vssd1 vssd1 vccd1 vccd1 net554 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout574_X net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout565 net566 vssd1 vssd1 vccd1 vccd1 net565 sky130_fd_sc_hd__buf_2
X_20027_ clknet_leaf_67_clk _00971_ net1473 vssd1 vssd1 vccd1 vccd1 ag2.body\[361\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_22_1587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout576 net577 vssd1 vssd1 vccd1 vccd1 net576 sky130_fd_sc_hd__buf_2
XANTENNA__17604__A2 net961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09838_ net1204 control.body\[921\] vssd1 vssd1 vccd1 vccd1 _04811_ sky130_fd_sc_hd__or2_1
Xfanout587 net589 vssd1 vssd1 vccd1 vccd1 net587 sky130_fd_sc_hd__clkbuf_4
Xfanout598 _06476_ vssd1 vssd1 vccd1 vccd1 net598 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10213__A net1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10152__A2 net1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout65_A net67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16378__Y _02057_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09561__X _04534_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout741_X net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09769_ ag2.body\[236\] net1136 vssd1 vssd1 vccd1 vccd1 _04742_ sky130_fd_sc_hd__xor2_1
XANTENNA_fanout839_X net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_38_clk clknet_4_5__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_38_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout1483_X net1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11800_ net468 _06746_ _06741_ _06661_ vssd1 vssd1 vccd1 vccd1 _06772_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_29_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_1459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12780_ net667 _07593_ vssd1 vssd1 vccd1 vccd1 _07594_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_29_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10867__B net1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15379__B1 _01594_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11731_ _06697_ _06699_ _06700_ _06702_ vssd1 vssd1 vccd1 vccd1 _06703_ sky130_fd_sc_hd__a22o_1
XFILLER_0_138_212 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16040__A1 net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14450_ net846 ag2.body\[224\] ag2.body\[230\] net804 _08610_ vssd1 vssd1 vccd1 vccd1
+ _08611_ sky130_fd_sc_hd__o221a_1
XFILLER_0_22_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11662_ net317 _06634_ net480 vssd1 vssd1 vccd1 vccd1 coll.nextBadColl sky130_fd_sc_hd__a21boi_1
XFILLER_0_132_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13401_ net312 _07553_ net673 vssd1 vssd1 vccd1 vccd1 _07873_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_94_3202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10613_ _05574_ _05575_ _05580_ _05585_ vssd1 vssd1 vccd1 vccd1 _05586_ sky130_fd_sc_hd__or4_2
X_14381_ _08534_ _08539_ _08540_ _08541_ vssd1 vssd1 vccd1 vccd1 _08542_ sky130_fd_sc_hd__or4b_2
X_11593_ obsg2.obstacleArray\[8\] obsg2.obstacleArray\[9\] obsg2.obstacleArray\[12\]
+ obsg2.obstacleArray\[13\] net1123 net513 vssd1 vssd1 vccd1 vccd1 _06566_ sky130_fd_sc_hd__mux4_1
X_16120_ obsg2.obstacleArray\[76\] net423 net373 _01798_ vssd1 vssd1 vccd1 vccd1 _01799_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_64_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13332_ net332 _07505_ _07813_ vssd1 vssd1 vccd1 vccd1 _07846_ sky130_fd_sc_hd__and3_1
XANTENNA__09449__A net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10544_ net641 _04599_ vssd1 vssd1 vccd1 vccd1 _05517_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_91_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16051_ net433 _01719_ vssd1 vssd1 vccd1 vccd1 _01730_ sky130_fd_sc_hd__nand2_1
XFILLER_0_126_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10475_ _05436_ _05437_ _05442_ _05447_ vssd1 vssd1 vccd1 vccd1 _05448_ sky130_fd_sc_hd__or4_1
X_13263_ net384 _07454_ vssd1 vssd1 vccd1 vccd1 _07819_ sky130_fd_sc_hd__nor2_1
X_15002_ _05178_ net58 vssd1 vssd1 vccd1 vccd1 _01552_ sky130_fd_sc_hd__nor2_4
X_12214_ _07177_ _07181_ _04259_ img_gen.control.current\[0\] vssd1 vssd1 vccd1 vccd1
+ _07185_ sky130_fd_sc_hd__o211a_1
X_13194_ _07787_ net263 _07785_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[364\]
+ sky130_fd_sc_hd__mux2_1
XANTENNA__14106__A1 net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14106__B2 net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19810_ clknet_leaf_89_clk _00754_ net1410 vssd1 vssd1 vccd1 vccd1 ag2.body\[576\]
+ sky130_fd_sc_hd__dfrtp_4
X_12145_ img_gen.tracker.frame\[513\] net583 net560 vssd1 vssd1 vccd1 vccd1 _07117_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_124_1070 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_3006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14090__A net1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12603__A net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_3017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12117__B1 net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16953_ ag2.body\[290\] net864 vssd1 vssd1 vccd1 vccd1 _02632_ sky130_fd_sc_hd__xor2_4
X_19741_ clknet_leaf_129_clk _00685_ net1325 vssd1 vssd1 vccd1 vccd1 control.body\[651\]
+ sky130_fd_sc_hd__dfrtp_1
X_12076_ img_gen.tracker.frame\[135\] net611 net556 img_gen.tracker.frame\[138\] vssd1
+ vssd1 vccd1 vccd1 _07048_ sky130_fd_sc_hd__a22o_1
XFILLER_0_40_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17056__B1 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15904_ ag2.body\[194\] net132 _01651_ ag2.body\[186\] vssd1 vssd1 vccd1 vccd1 _01140_
+ sky130_fd_sc_hd__a22o_1
X_11027_ net1181 control.body\[1042\] vssd1 vssd1 vccd1 vccd1 _06000_ sky130_fd_sc_hd__xor2_1
X_19672_ clknet_leaf_134_clk _00616_ net1309 vssd1 vssd1 vccd1 vccd1 control.body\[726\]
+ sky130_fd_sc_hd__dfrtp_1
X_16884_ _03981_ net868 net858 _03982_ _02562_ vssd1 vssd1 vccd1 vccd1 _02563_ sky130_fd_sc_hd__a221o_1
XANTENNA__10123__A net1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11340__B2 _05856_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18623_ clknet_leaf_3_clk img_gen.tracker.next_frame\[61\] net1250 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[61\] sky130_fd_sc_hd__dfrtp_1
X_15835_ ag2.body\[261\] net204 net49 ag2.body\[253\] vssd1 vssd1 vccd1 vccd1 _01079_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_91_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_29_clk clknet_4_4__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_29_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_56_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18554_ clknet_leaf_37_clk _00080_ net1351 vssd1 vssd1 vccd1 vccd1 control.divider.fsm.current_mode\[0\]
+ sky130_fd_sc_hd__dfstp_1
X_15766_ ag2.body\[327\] net215 _01636_ ag2.body\[319\] vssd1 vssd1 vccd1 vccd1 _01017_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_99_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_1452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12978_ img_gen.tracker.frame\[251\] net646 _07684_ vssd1 vssd1 vccd1 vccd1 _07685_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_86_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17505_ ag2.body\[235\] net719 net692 ag2.body\[239\] vssd1 vssd1 vccd1 vccd1 _03184_
+ sky130_fd_sc_hd__a22o_1
X_14717_ net1032 ag2.body\[341\] vssd1 vssd1 vccd1 vccd1 _08878_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_16_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18485_ net1516 net1510 vssd1 vssd1 vccd1 vccd1 _00016_ sky130_fd_sc_hd__or2_1
X_11929_ _06894_ _06900_ net470 vssd1 vssd1 vccd1 vccd1 _06901_ sky130_fd_sc_hd__mux2_1
X_15697_ ag2.body\[378\] net130 _01628_ ag2.body\[370\] vssd1 vssd1 vccd1 vccd1 _00956_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_86_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17436_ _04042_ net966 net708 ag2.body\[149\] vssd1 vssd1 vccd1 vccd1 _03115_ sky130_fd_sc_hd__o22a_1
XFILLER_0_12_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14648_ net828 ag2.body\[514\] _04191_ net1039 _08808_ vssd1 vssd1 vccd1 vccd1 _08809_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_117_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_17 _08236_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_28 _03442_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17367_ net1044 net1043 vssd1 vssd1 vccd1 vccd1 _03046_ sky130_fd_sc_hd__nand2_1
XANTENNA_39 _08924_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14265__A net999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14579_ net833 ag2.body\[489\] ag2.body\[494\] net800 vssd1 vssd1 vccd1 vccd1 _08740_
+ sky130_fd_sc_hd__a22o_1
X_19106_ clknet_leaf_1_clk img_gen.tracker.next_frame\[544\] net1244 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[544\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16318_ obsg2.obstacleArray\[70\] obsg2.obstacleArray\[71\] net409 vssd1 vssd1 vccd1
+ vccd1 _01997_ sky130_fd_sc_hd__mux2_1
XANTENNA__11800__C1 _06661_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17298_ ag2.body\[347\] net855 vssd1 vssd1 vccd1 vccd1 _02977_ sky130_fd_sc_hd__nand2_1
XFILLER_0_15_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19037_ clknet_leaf_6_clk img_gen.tracker.next_frame\[475\] net1264 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[475\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__14345__A1 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17576__A ag2.body\[342\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16249_ net354 _01892_ vssd1 vssd1 vccd1 vccd1 _01928_ sky130_fd_sc_hd__or2_1
XANTENNA__14345__B2 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11401__B net1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_1566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_482 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17295__B net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_120_Left_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_1599 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10017__B net1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16098__A1 _01728_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12108__B1 net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12513__A _06638_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09094__A ag2.body\[337\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19939_ clknet_leaf_46_clk _00883_ net1376 vssd1 vssd1 vccd1 vccd1 ag2.body\[449\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__12659__A1 net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13856__B1 _08134_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17047__B1 net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13320__A2 net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09623_ net783 control.body\[800\] control.body\[804\] net758 _04595_ vssd1 vssd1
+ vccd1 vccd1 _04596_ sky130_fd_sc_hd__o221a_1
XANTENNA__10968__A net1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout367_A _02067_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09554_ net1050 control.body\[727\] vssd1 vssd1 vccd1 vccd1 _04527_ sky130_fd_sc_hd__or2_1
XANTENNA__10687__B net1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09485_ _04447_ _04457_ _04444_ vssd1 vssd1 vccd1 vccd1 _04458_ sky130_fd_sc_hd__o21ai_1
XANTENNA__11634__A2 net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12831__A1 net239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1276_A net1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17770__A1 _03193_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20427__CLK clknet_leaf_37_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14584__A1 net1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_237 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14584__B2 net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout701_A net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14175__A net1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1064_X net1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20576_ clknet_leaf_106_clk _01434_ _00040_ vssd1 vssd1 vccd1 vccd1 sound_gen.dac1.dacCount\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14336__A1 net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14336__B2 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11311__B net1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14462__X _08623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16730__C1 net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10208__A net1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1231_X net1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14903__A net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10260_ net1049 control.body\[791\] vssd1 vssd1 vccd1 vccd1 _05233_ sky130_fd_sc_hd__xnor2_1
XANTENNA__17412__A2_N net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout691_X net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12898__A1 net245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout789_X net789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10191_ ag2.body\[114\] net1186 vssd1 vssd1 vccd1 vccd1 _05164_ sky130_fd_sc_hd__or2_1
XANTENNA__12423__A net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1305 net1306 vssd1 vssd1 vccd1 vccd1 net1305 sky130_fd_sc_hd__clkbuf_2
Xfanout1316 net1324 vssd1 vssd1 vccd1 vccd1 net1316 sky130_fd_sc_hd__clkbuf_2
XANTENNA__10555__D_N _05517_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1327 net1330 vssd1 vssd1 vccd1 vccd1 net1327 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout956_X net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16389__X _02068_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1338 net1357 vssd1 vssd1 vccd1 vccd1 net1338 sky130_fd_sc_hd__clkbuf_4
Xfanout340 _07309_ vssd1 vssd1 vccd1 vccd1 net340 sky130_fd_sc_hd__clkbuf_2
Xfanout1349 net1350 vssd1 vssd1 vccd1 vccd1 net1349 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_121_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17038__B1 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout351 _01703_ vssd1 vssd1 vccd1 vccd1 net351 sky130_fd_sc_hd__clkbuf_4
Xfanout362 _02222_ vssd1 vssd1 vccd1 vccd1 net362 sky130_fd_sc_hd__clkbuf_4
X_13950_ ag2.body\[91\] net191 _08155_ ag2.body\[83\] vssd1 vssd1 vccd1 vccd1 _00172_
+ sky130_fd_sc_hd__a22o_1
Xfanout373 net375 vssd1 vssd1 vccd1 vccd1 net373 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_1384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17589__A1 ag2.body\[58\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout384 _06723_ vssd1 vssd1 vccd1 vccd1 net384 sky130_fd_sc_hd__clkbuf_4
XANTENNA__14672__A1_N net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout395 net396 vssd1 vssd1 vccd1 vccd1 net395 sky130_fd_sc_hd__clkbuf_4
XANTENNA__17589__B2 ag2.body\[61\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12901_ net293 _07647_ _07648_ net1912 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[209\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_96_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11981__B net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13881_ ag2.body\[30\] net115 _08147_ ag2.body\[22\] vssd1 vssd1 vccd1 vccd1 _00111_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11873__A2 net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15620_ ag2.body\[453\] net124 _01613_ ag2.body\[445\] vssd1 vssd1 vccd1 vccd1 _00887_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12796__C net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13254__A net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12832_ net261 _07616_ _07617_ net1826 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[172\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__09451__B net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13075__A1 net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09818__A2 net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14069__B ag2.body\[214\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11086__B1 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15551_ ag2.body\[504\] net188 _01612_ ag2.body\[496\] vssd1 vssd1 vccd1 vccd1 _00826_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_16_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11625__A2 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12763_ net684 _07585_ vssd1 vssd1 vccd1 vccd1 _07586_ sky130_fd_sc_hd__nor2_1
XFILLER_0_96_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14502_ _08655_ _08656_ _08661_ _08662_ vssd1 vssd1 vccd1 vccd1 _08663_ sky130_fd_sc_hd__or4_1
XFILLER_0_96_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18270_ _03549_ _03563_ _03564_ obsg2.obstacleArray\[132\] vssd1 vssd1 vccd1 vccd1
+ _03774_ sky130_fd_sc_hd__a31o_1
XFILLER_0_83_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11714_ img_gen.tracker.frame\[335\] net590 net576 vssd1 vssd1 vccd1 vccd1 _06686_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_84_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15482_ ag2.body\[570\] net112 _01605_ ag2.body\[562\] vssd1 vssd1 vccd1 vccd1 _00764_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_12_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10884__Y _05857_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12694_ net238 net310 _07551_ _07552_ net1609 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[99\]
+ sky130_fd_sc_hd__a32o_1
X_17221_ ag2.body\[314\] net866 vssd1 vssd1 vccd1 vccd1 _02900_ sky130_fd_sc_hd__xor2_1
X_14433_ net970 ag2.body\[19\] vssd1 vssd1 vccd1 vccd1 _08594_ sky130_fd_sc_hd__xor2_1
X_11645_ _06616_ _06617_ net507 vssd1 vssd1 vccd1 vccd1 _06618_ sky130_fd_sc_hd__mux2_1
XANTENNA__14610__A1_N net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17152_ _02825_ _02826_ _02830_ vssd1 vssd1 vccd1 vccd1 _02831_ sky130_fd_sc_hd__a21o_1
XFILLER_0_25_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14364_ net1026 ag2.body\[605\] vssd1 vssd1 vccd1 vccd1 _08525_ sky130_fd_sc_hd__xnor2_1
X_11576_ net505 _06547_ _06548_ _06546_ net1126 vssd1 vssd1 vccd1 vccd1 _06549_ sky130_fd_sc_hd__a221o_1
XANTENNA__12050__A2 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_5_clk_X clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_1554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16103_ obsg2.obstacleArray\[64\] net426 net374 _01781_ vssd1 vssd1 vccd1 vccd1 _01782_
+ sky130_fd_sc_hd__o211a_1
XANTENNA__14327__A1 net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13315_ net229 _07839_ _07840_ net1927 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[432\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__18967__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_1576 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14327__B2 net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17083_ _02758_ _02759_ _02760_ _02761_ vssd1 vssd1 vccd1 vccd1 _02762_ sky130_fd_sc_hd__a22o_1
X_10527_ net1204 control.body\[913\] vssd1 vssd1 vccd1 vccd1 _05500_ sky130_fd_sc_hd__xor2_1
XFILLER_0_122_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14295_ net1006 _04172_ _08454_ _08455_ vssd1 vssd1 vccd1 vccd1 _08456_ sky130_fd_sc_hd__a211o_1
XANTENNA__10118__A net1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10600__A3 _04238_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14813__A net1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16034_ net460 net495 vssd1 vssd1 vccd1 vccd1 _01713_ sky130_fd_sc_hd__nor2_1
X_10458_ ag2.body\[451\] net1153 vssd1 vssd1 vccd1 vccd1 _05431_ sky130_fd_sc_hd__xor2_1
X_13246_ net384 net338 _07439_ vssd1 vssd1 vccd1 vccd1 _07811_ sky130_fd_sc_hd__or3_1
XFILLER_0_126_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_111_3699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_1284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13177_ img_gen.tracker.frame\[355\] net646 vssd1 vssd1 vccd1 vccd1 _07780_ sky130_fd_sc_hd__and2_1
X_10389_ net1060 control.body\[1063\] vssd1 vssd1 vccd1 vccd1 _05362_ sky130_fd_sc_hd__nand2_1
XANTENNA__13148__B net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12128_ img_gen.tracker.frame\[573\] net588 vssd1 vssd1 vccd1 vccd1 _07100_ sky130_fd_sc_hd__or2_1
X_17985_ net354 _03603_ vssd1 vssd1 vccd1 vccd1 _03604_ sky130_fd_sc_hd__or2_1
XFILLER_0_104_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17029__B1 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12059_ img_gen.tracker.frame\[48\] net627 net609 img_gen.tracker.frame\[51\] vssd1
+ vssd1 vccd1 vccd1 _07031_ sky130_fd_sc_hd__a22o_1
X_19724_ clknet_leaf_133_clk net2256 net1305 vssd1 vssd1 vccd1 vccd1 control.body\[666\]
+ sky130_fd_sc_hd__dfrtp_1
X_16936_ ag2.body\[523\] net854 vssd1 vssd1 vccd1 vccd1 _02615_ sky130_fd_sc_hd__xor2_1
XFILLER_0_79_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09642__A net1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16867_ ag2.body\[467\] net848 vssd1 vssd1 vccd1 vccd1 _02546_ sky130_fd_sc_hd__nand2_1
X_19655_ clknet_leaf_133_clk _00599_ net1308 vssd1 vssd1 vccd1 vccd1 control.body\[741\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__15363__B net53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16788__C1 net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11864__A2 net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10788__A net1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17885__B1_N obsg2.obstacleCount\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13164__A net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15818_ ag2.body\[277\] net206 _01642_ ag2.body\[269\] vssd1 vssd1 vccd1 vccd1 _01063_
+ sky130_fd_sc_hd__a22o_1
X_18606_ clknet_leaf_16_clk img_gen.tracker.next_frame\[44\] net1318 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[44\] sky130_fd_sc_hd__dfrtp_1
X_19586_ clknet_leaf_118_clk _00530_ net1388 vssd1 vssd1 vccd1 vccd1 control.body\[800\]
+ sky130_fd_sc_hd__dfrtp_1
X_16798_ obsg2.obstacleArray\[132\] obsg2.obstacleArray\[133\] net457 vssd1 vssd1
+ vccd1 vccd1 _02477_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_430 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18537_ clknet_leaf_136_clk _00063_ net1300 vssd1 vssd1 vccd1 vccd1 img_gen.updater.commands.count\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_15749_ _05255_ net60 vssd1 vssd1 vccd1 vccd1 _01635_ sky130_fd_sc_hd__nor2_2
XANTENNA__17201__B1 net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09270_ sound_gen.osc1.stayCount\[12\] _04287_ _04288_ sound_gen.osc1.stayCount\[14\]
+ sound_gen.osc1.stayCount\[13\] vssd1 vssd1 vccd1 vccd1 _04293_ sky130_fd_sc_hd__a221o_1
X_18468_ _04261_ _03951_ _03953_ _03954_ vssd1 vssd1 vccd1 vccd1 _01424_ sky130_fd_sc_hd__o211a_1
XANTENNA__16555__A2 net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1119 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14566__A1 net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17419_ _03092_ _03093_ _03096_ _03097_ vssd1 vssd1 vccd1 vccd1 _03098_ sky130_fd_sc_hd__or4_4
XFILLER_0_1_1518 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14566__B2 net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18399_ net326 _03785_ _03888_ net464 vssd1 vssd1 vccd1 vccd1 _03889_ sky130_fd_sc_hd__a211o_1
X_20430_ clknet_leaf_23_clk _01317_ net1359 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[66\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__11412__A net1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20361_ clknet_leaf_21_clk _00001_ net1361 vssd1 vssd1 vccd1 vccd1 obsg2.obsNeeded\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09993__A1 net1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16414__S net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09993__B2 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_9_clk clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_9_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_3_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_1086 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20292_ clknet_leaf_37_clk control.divider.next_count\[13\] net1350 vssd1 vssd1 vccd1
+ vccd1 control.divider.count\[13\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_45_1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17268__B1 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1024_A ag2.randCord\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19122__CLK clknet_leaf_141_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20233__Q ag2.body\[167\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08985_ ag2.body\[79\] vssd1 vssd1 vccd1 vccd1 _04010_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout484_A _02373_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09552__A net1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15273__B net54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11855__A2 net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10698__A _04471_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout749_A _04233_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09606_ net1097 control.body\[637\] vssd1 vssd1 vccd1 vccd1 _04579_ sky130_fd_sc_hd__xor2_1
XFILLER_0_97_238 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13057__A1 net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13505__C _07813_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09537_ net769 control.body\[1027\] vssd1 vssd1 vccd1 vccd1 _04510_ sky130_fd_sc_hd__and2_1
XANTENNA__11306__B net1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11607__A2 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12804__A1 net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1181_X net1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09468_ ag2.body\[378\] net774 net768 ag2.body\[379\] vssd1 vssd1 vccd1 vccd1 _04441_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_109_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09681__B1 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16546__A2 net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout704_X net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09399_ _04344_ _04383_ vssd1 vssd1 vccd1 vccd1 _01403_ sky130_fd_sc_hd__nor2_1
XFILLER_0_30_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11430_ ag2.body\[394\] net1185 vssd1 vssd1 vccd1 vccd1 _06403_ sky130_fd_sc_hd__or2_1
XFILLER_0_11_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20628_ sound_gen.dac1.dacCount\[6\] vssd1 vssd1 vccd1 vccd1 net15 sky130_fd_sc_hd__clkbuf_1
XANTENNA__12032__A2 net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12137__B net616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16832__B net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11361_ _06332_ _06333_ vssd1 vssd1 vccd1 vccd1 _06334_ sky130_fd_sc_hd__nand2_1
X_20559_ clknet_leaf_109_clk toggle1.nextBlinkToggle\[1\] net1416 vssd1 vssd1 vccd1
+ vccd1 net26 sky130_fd_sc_hd__dfrtp_1
XANTENNA__16324__S net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14633__A net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18105__A net38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10312_ _05277_ _05278_ _05280_ _05281_ _05274_ vssd1 vssd1 vccd1 vccd1 _05285_ sky130_fd_sc_hd__a221o_1
X_13100_ net683 _07742_ vssd1 vssd1 vccd1 vccd1 _07743_ sky130_fd_sc_hd__nor2_1
XFILLER_0_120_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11292_ _06254_ _06255_ _06256_ _06259_ vssd1 vssd1 vccd1 vccd1 _06265_ sky130_fd_sc_hd__or4_1
X_14080_ net1007 ag2.body\[567\] vssd1 vssd1 vccd1 vccd1 _08241_ sky130_fd_sc_hd__xor2_1
XFILLER_0_127_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10880__B net1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10243_ ag2.body\[324\] net1141 vssd1 vssd1 vccd1 vccd1 _05216_ sky130_fd_sc_hd__or2_1
X_13031_ net342 _07539_ vssd1 vssd1 vccd1 vccd1 _07710_ sky130_fd_sc_hd__nor2_1
XANTENNA__13249__A net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_1349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17944__A net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09446__B net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10174_ ag2.body\[416\] net1234 vssd1 vssd1 vccd1 vccd1 _05147_ sky130_fd_sc_hd__xor2_1
XFILLER_0_101_1614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1102 net1103 vssd1 vssd1 vccd1 vccd1 net1102 sky130_fd_sc_hd__clkbuf_4
Xfanout1113 net1117 vssd1 vssd1 vccd1 vccd1 net1113 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_101_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1124 net1129 vssd1 vssd1 vccd1 vccd1 net1124 sky130_fd_sc_hd__clkbuf_2
Xfanout1135 net1137 vssd1 vssd1 vccd1 vccd1 net1135 sky130_fd_sc_hd__buf_2
X_17770_ _03193_ _03196_ _02861_ vssd1 vssd1 vccd1 vccd1 _03449_ sky130_fd_sc_hd__o21a_1
Xfanout1146 net1147 vssd1 vssd1 vccd1 vccd1 net1146 sky130_fd_sc_hd__buf_2
Xfanout1157 net1158 vssd1 vssd1 vccd1 vccd1 net1157 sky130_fd_sc_hd__buf_4
X_14982_ net2223 net158 _01550_ net2237 vssd1 vssd1 vccd1 vccd1 _00319_ sky130_fd_sc_hd__a22o_1
XANTENNA__13296__A1 net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1168 net1173 vssd1 vssd1 vccd1 vccd1 net1168 sky130_fd_sc_hd__clkbuf_2
Xfanout170 net171 vssd1 vssd1 vccd1 vccd1 net170 sky130_fd_sc_hd__buf_2
Xfanout1179 net1180 vssd1 vssd1 vccd1 vccd1 net1179 sky130_fd_sc_hd__buf_4
Xfanout181 net182 vssd1 vssd1 vccd1 vccd1 net181 sky130_fd_sc_hd__buf_2
X_16721_ obsg2.obstacleArray\[108\] net490 net486 obsg2.obstacleArray\[110\] vssd1
+ vssd1 vccd1 vccd1 _02400_ sky130_fd_sc_hd__a22o_1
Xfanout192 net218 vssd1 vssd1 vccd1 vccd1 net192 sky130_fd_sc_hd__clkbuf_2
X_13933_ ag2.body\[76\] net186 _08153_ ag2.body\[68\] vssd1 vssd1 vccd1 vccd1 _00157_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__18548__Q ag2.y\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11846__A2 net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12600__B net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1244 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19440_ clknet_leaf_108_clk _00384_ net1421 vssd1 vssd1 vccd1 vccd1 control.body\[958\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_44_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16652_ obsg2.obstacleArray\[4\] obsg2.obstacleArray\[5\] net446 vssd1 vssd1 vccd1
+ vccd1 _02331_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13864_ track.nextHighScore\[2\] net322 track.nextHighScore\[6\] _08137_ vssd1 vssd1
+ vccd1 vccd1 _08138_ sky130_fd_sc_hd__a31o_1
XFILLER_0_9_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19765__CLK clknet_leaf_127_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_3481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15603_ ag2.body\[469\] net121 _01619_ ag2.body\[461\] vssd1 vssd1 vccd1 vccd1 _00871_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_104_3492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14796__A1 net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12815_ net261 _07608_ _07609_ net1795 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[163\]
+ sky130_fd_sc_hd__a22o_1
X_19371_ clknet_leaf_102_clk _00315_ net1426 vssd1 vssd1 vccd1 vccd1 control.body\[1017\]
+ sky130_fd_sc_hd__dfrtp_1
X_16583_ _02208_ _02261_ vssd1 vssd1 vccd1 vccd1 _02262_ sky130_fd_sc_hd__or2_1
XANTENNA__14796__B2 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13795_ img_gen.updater.commands.count\[15\] _08099_ vssd1 vssd1 vccd1 vccd1 _08101_
+ sky130_fd_sc_hd__or2_1
XANTENNA__14808__A net1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18322_ _03789_ _03817_ _03785_ vssd1 vssd1 vccd1 vccd1 _03818_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_29_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_100_3367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15534_ ag2.body\[520\] net160 _01611_ ag2.body\[512\] vssd1 vssd1 vccd1 vccd1 _00810_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_100_3378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12746_ net237 _07576_ _07577_ net1672 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[126\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_60_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18253_ obsg2.obstacleArray\[123\] _03765_ net525 vssd1 vssd1 vccd1 vccd1 _01374_
+ sky130_fd_sc_hd__o21a_1
XANTENNA__10282__A1 _04982_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11503__Y _06476_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15465_ ag2.body\[587\] net108 _01603_ ag2.body\[579\] vssd1 vssd1 vccd1 vccd1 _00749_
+ sky130_fd_sc_hd__a22o_1
X_12677_ net241 _07543_ _07544_ net2163 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[90\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_38_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17204_ _02879_ _02880_ _02882_ vssd1 vssd1 vccd1 vccd1 _02883_ sky130_fd_sc_hd__or3_1
XFILLER_0_25_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14416_ net828 ag2.body\[530\] ag2.body\[535\] net794 vssd1 vssd1 vccd1 vccd1 _08577_
+ sky130_fd_sc_hd__a22o_1
X_18184_ _03625_ net41 vssd1 vssd1 vccd1 vccd1 _03731_ sky130_fd_sc_hd__nor2_1
X_11628_ net506 _06597_ _06600_ vssd1 vssd1 vccd1 vccd1 _06601_ sky130_fd_sc_hd__o21a_1
XFILLER_0_128_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15396_ net2188 net80 _01596_ net2315 vssd1 vssd1 vccd1 vccd1 _00687_ sky130_fd_sc_hd__a22o_1
XANTENNA__12023__A2 net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_3886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_117_3897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09975__A1 _04421_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17135_ ag2.body\[519\] net932 vssd1 vssd1 vccd1 vccd1 _02814_ sky130_fd_sc_hd__or2_1
XANTENNA__10263__A1_N _05211_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14347_ _08502_ _08503_ _08504_ _08505_ vssd1 vssd1 vccd1 vccd1 _08508_ sky130_fd_sc_hd__or4_1
XFILLER_0_68_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11559_ net505 _06530_ _06531_ net1124 vssd1 vssd1 vccd1 vccd1 _06532_ sky130_fd_sc_hd__a211o_1
XFILLER_0_53_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18015__A net45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14543__A net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold607 control.body\[1115\] vssd1 vssd1 vccd1 vccd1 net2169 sky130_fd_sc_hd__dlygate4sd3_1
Xhold618 _00281_ vssd1 vssd1 vccd1 vccd1 net2180 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17066_ ag2.body\[24\] net880 vssd1 vssd1 vccd1 vccd1 _02745_ sky130_fd_sc_hd__nand2_1
Xhold629 control.body\[784\] vssd1 vssd1 vccd1 vccd1 net2191 sky130_fd_sc_hd__dlygate4sd3_1
X_14278_ net1040 ag2.body\[140\] vssd1 vssd1 vccd1 vccd1 _08439_ sky130_fd_sc_hd__xor2_1
XFILLER_0_100_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1551 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16017_ net860 _01684_ vssd1 vssd1 vccd1 vccd1 _01696_ sky130_fd_sc_hd__nor2_1
XANTENNA__14720__A1 net1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13229_ _07804_ net263 _07802_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[382\]
+ sky130_fd_sc_hd__mux2_1
XANTENNA__13523__A2 net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14720__B2 net1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14830__X _01501_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11534__A1 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20053__Q ag2.body\[339\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19295__CLK clknet_leaf_98_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13287__A1 net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17968_ net43 vssd1 vssd1 vccd1 vccd1 _03592_ sky130_fd_sc_hd__inv_2
XFILLER_0_97_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15093__B net58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19707_ clknet_leaf_134_clk _00651_ net1307 vssd1 vssd1 vccd1 vccd1 control.body\[681\]
+ sky130_fd_sc_hd__dfrtp_1
X_16919_ ag2.body\[563\] net716 net705 ag2.body\[565\] vssd1 vssd1 vccd1 vccd1 _02598_
+ sky130_fd_sc_hd__o22a_1
XANTENNA__11837__A2 net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17899_ net351 _03533_ vssd1 vssd1 vccd1 vccd1 _03535_ sky130_fd_sc_hd__and2_1
XFILLER_0_117_1610 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13039__A1 net233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19638_ clknet_leaf_123_clk _00582_ net1406 vssd1 vssd1 vccd1 vccd1 control.body\[756\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_0_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16776__A2 net494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16917__B net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11126__B net1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14787__A1 net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15821__B net59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19569_ clknet_leaf_116_clk _00513_ net1387 vssd1 vssd1 vccd1 vccd1 control.body\[831\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14787__B2 net974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14718__A net1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09322_ sound_gen.at_max sound_gen.dac1.dacCount\[1\] sound_gen.dac1.dacCount\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04334_ sky130_fd_sc_hd__and3_1
XANTENNA__19977__RESET_B net1470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09253_ img_gen.updater.commands.rR1.rainbowRNG\[5\] vssd1 vssd1 vccd1 vccd1 _04278_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_63_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout232_A net233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20228__Q ag2.body\[162\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09184_ ag2.body\[577\] vssd1 vssd1 vccd1 vccd1 _04209_ sky130_fd_sc_hd__inv_2
XANTENNA__13211__A1 net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20413_ clknet_leaf_33_clk _01300_ net1352 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[49\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__17489__B1 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10981__A net1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14453__A net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1141_A net1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1239_A net1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20344_ clknet_leaf_140_clk _01235_ net1293 vssd1 vssd1 vccd1 vccd1 img_gen.updater.commands.rR1.rainbowRNG\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_47_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16700__A2 net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout699_A net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09718__B2 net1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20275_ clknet_leaf_36_clk net3 net1347 vssd1 vssd1 vccd1 vccd1 control.button2.Q\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_41_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1027_X net1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10328__A2 _05286_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout866_A net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout487_X net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_127_4182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17661__B1 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_4193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08968_ ag2.body\[53\] vssd1 vssd1 vccd1 vccd1 _03993_ sky130_fd_sc_hd__inv_2
XANTENNA__19788__CLK clknet_leaf_127_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout654_X net654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17413__B1 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10930_ net755 control.body\[1037\] control.body\[1033\] net780 vssd1 vssd1 vccd1
+ vccd1 _05903_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__11637__A_N _06511_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09766__D_N _04539_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16827__B net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15731__B net60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11036__B net1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout821_X net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10861_ net1121 control.body\[692\] vssd1 vssd1 vccd1 vccd1 _05834_ sky130_fd_sc_hd__xor2_1
XANTENNA__14778__B2 net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout919_X net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12600_ net580 net471 net569 _07312_ vssd1 vssd1 vccd1 vccd1 _07501_ sky130_fd_sc_hd__or4_1
XFILLER_0_38_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13580_ control.divider.count\[6\] _07949_ _07950_ control.divider.count\[5\] vssd1
+ vssd1 vccd1 vccd1 _07955_ sky130_fd_sc_hd__o22a_1
XFILLER_0_6_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_967 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10792_ _05761_ _05763_ _05764_ _05685_ vssd1 vssd1 vccd1 vccd1 _05765_ sky130_fd_sc_hd__or4b_1
XFILLER_0_52_1163 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19199__Q ag2.body\[62\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10875__B net1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10264__A1 net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12531_ net283 net334 _07444_ _07460_ _07462_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[26\]
+ sky130_fd_sc_hd__a41o_1
XANTENNA__13251__B net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17939__A net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19168__CLK clknet_leaf_52_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15250_ control.body\[780\] net99 _01579_ net2103 vssd1 vssd1 vccd1 vccd1 _00558_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_30_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12462_ net678 _07419_ vssd1 vssd1 vccd1 vccd1 _07420_ sky130_fd_sc_hd__nor2_1
XFILLER_0_129_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17658__B net866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14201_ net833 ag2.body\[361\] ag2.body\[362\] net826 vssd1 vssd1 vccd1 vccd1 _08362_
+ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_10_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11413_ net1100 control.body\[853\] vssd1 vssd1 vccd1 vccd1 _06386_ sky130_fd_sc_hd__or2_1
XANTENNA__09957__A1 _04421_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15181_ control.body\[847\] net103 _01571_ net2401 vssd1 vssd1 vccd1 vccd1 _00497_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_129_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12393_ _07318_ _07332_ _07337_ _07357_ vssd1 vssd1 vccd1 vccd1 _07358_ sky130_fd_sc_hd__a31o_1
XANTENNA__10891__A net1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14363__A net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10077__A2_N net479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10567__A2 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14132_ net1009 ag2.body\[175\] vssd1 vssd1 vccd1 vccd1 _08293_ sky130_fd_sc_hd__nand2_1
XFILLER_0_65_1557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11344_ ag2.body\[447\] net1055 vssd1 vssd1 vccd1 vccd1 _06317_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_112_3750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_558 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_709 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18940_ clknet_leaf_139_clk img_gen.tracker.next_frame\[378\] net1288 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[378\] sky130_fd_sc_hd__dfrtp_1
X_14063_ _08215_ _08216_ _08218_ _08219_ vssd1 vssd1 vccd1 vccd1 _08224_ sky130_fd_sc_hd__or4_1
X_11275_ ag2.body\[123\] net1164 vssd1 vssd1 vccd1 vccd1 _06248_ sky130_fd_sc_hd__xor2_1
XANTENNA__11516__A1 net1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13014_ net342 _07527_ vssd1 vssd1 vccd1 vccd1 _07702_ sky130_fd_sc_hd__nor2_1
XFILLER_0_98_1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17393__B net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10226_ ag2.body\[566\] net1077 vssd1 vssd1 vccd1 vccd1 _05199_ sky130_fd_sc_hd__xor2_1
X_18871_ clknet_leaf_22_clk img_gen.tracker.next_frame\[309\] net1358 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[309\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__18444__A2 _04791_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17961__X _03586_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17822_ _03486_ _03487_ vssd1 vssd1 vccd1 vccd1 _03488_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_100_490 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10157_ _03996_ net1128 _04232_ ag2.body\[61\] _05125_ vssd1 vssd1 vccd1 vccd1 _05130_
+ sky130_fd_sc_hd__a221o_1
XANTENNA__17652__B1 net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09904__B net1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold4 control.button2.Q\[0\] vssd1 vssd1 vccd1 vccd1 net1566 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_1620 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_106_3543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10088_ net1172 _04242_ control.body\[797\] net753 _05060_ vssd1 vssd1 vccd1 vccd1
+ _05061_ sky130_fd_sc_hd__a221o_1
X_14965_ control.body\[1039\] net172 _01547_ net2525 vssd1 vssd1 vccd1 vccd1 _00305_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11819__A2 net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17753_ _02868_ _02873_ _02897_ _02961_ _03431_ vssd1 vssd1 vccd1 vccd1 _03432_ sky130_fd_sc_hd__o2111a_1
XTAP_TAPCELL_ROW_106_3554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10402__Y _05375_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_3565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1604 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16704_ _02380_ _02382_ net497 vssd1 vssd1 vccd1 vccd1 _02383_ sky130_fd_sc_hd__mux2_1
X_13916_ ag2.body\[61\] net129 _08151_ ag2.body\[53\] vssd1 vssd1 vccd1 vccd1 _00142_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_57_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17684_ ag2.body\[473\] net730 net710 ag2.body\[476\] vssd1 vssd1 vccd1 vccd1 _03363_
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_18_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10131__A net1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_3429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14896_ net2178 net178 _01540_ control.body\[1081\] vssd1 vssd1 vccd1 vccd1 _00243_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_57_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16758__A2 net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16635_ obsg2.obstacleArray\[59\] net450 net391 _02313_ vssd1 vssd1 vccd1 vccd1 _02314_
+ sky130_fd_sc_hd__o211a_1
X_19423_ clknet_leaf_107_clk _00367_ net1434 vssd1 vssd1 vccd1 vccd1 control.body\[973\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__15641__B net64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13847_ ag2.body\[11\] net127 _08133_ ag2.body\[3\] vssd1 vssd1 vccd1 vccd1 _00091_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_134_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16566_ obsg2.obstacleArray\[122\] net444 vssd1 vssd1 vccd1 vccd1 _02245_ sky130_fd_sc_hd__or2_1
X_19354_ clknet_leaf_101_clk _00298_ net1438 vssd1 vssd1 vccd1 vccd1 control.body\[1032\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_80_2750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13778_ img_gen.updater.commands.count\[10\] _08086_ _08070_ vssd1 vssd1 vccd1 vccd1
+ _08089_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_80_2761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_904 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_80_2772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18305_ track.nextHighScore\[1\] net326 net325 vssd1 vssd1 vccd1 vccd1 _03801_ sky130_fd_sc_hd__o21a_1
X_15517_ ag2.body\[537\] net155 _01609_ ag2.body\[529\] vssd1 vssd1 vccd1 vccd1 _00795_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_119_3948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12729_ net237 _07568_ _07569_ net1606 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[117\]
+ sky130_fd_sc_hd__a22o_1
X_19285_ clknet_leaf_98_clk _00229_ net1446 vssd1 vssd1 vccd1 vccd1 control.body\[1107\]
+ sky130_fd_sc_hd__dfrtp_1
X_16497_ net365 _02175_ _02174_ _02076_ vssd1 vssd1 vccd1 vccd1 _02176_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_119_3959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_61_2171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_2182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_2193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18236_ _03677_ net37 obsg2.obstacleArray\[115\] vssd1 vssd1 vccd1 vccd1 _03757_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_44_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15448_ ag2.body\[604\] net86 _01601_ ag2.body\[596\] vssd1 vssd1 vccd1 vccd1 _00734_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_5_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16930__A2 net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18167_ net532 _03722_ vssd1 vssd1 vccd1 vccd1 _01331_ sky130_fd_sc_hd__and2_1
XFILLER_0_83_1613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15379_ net2241 net69 _01594_ net2493 vssd1 vssd1 vccd1 vccd1 _00672_ sky130_fd_sc_hd__a22o_1
XFILLER_0_41_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold404 img_gen.tracker.frame\[57\] vssd1 vssd1 vccd1 vccd1 net1966 sky130_fd_sc_hd__dlygate4sd3_1
X_17118_ ag2.body\[540\] net963 vssd1 vssd1 vccd1 vccd1 _02797_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_78_2690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18098_ _03545_ _03613_ vssd1 vssd1 vccd1 vccd1 _03681_ sky130_fd_sc_hd__nand2_1
XANTENNA__16143__B1 net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold415 img_gen.tracker.frame\[212\] vssd1 vssd1 vccd1 vccd1 net1977 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12064__Y _07036_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold426 img_gen.tracker.frame\[477\] vssd1 vssd1 vccd1 vccd1 net1988 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold437 img_gen.tracker.frame\[282\] vssd1 vssd1 vccd1 vccd1 net1999 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12505__B _06638_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_2565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold448 img_gen.tracker.frame\[41\] vssd1 vssd1 vccd1 vccd1 net2010 sky130_fd_sc_hd__dlygate4sd3_1
X_17049_ ag2.body\[260\] net711 net740 ag2.body\[256\] vssd1 vssd1 vccd1 vccd1 _02728_
+ sky130_fd_sc_hd__a2bb2o_1
X_09940_ ag2.body\[28\] net1128 vssd1 vssd1 vccd1 vccd1 _04913_ sky130_fd_sc_hd__xor2_1
Xhold459 img_gen.tracker.frame\[508\] vssd1 vssd1 vccd1 vccd1 net2021 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_74_2587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10306__A net1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_115_Right_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20060_ clknet_leaf_72_clk _01004_ net1500 vssd1 vssd1 vccd1 vccd1 ag2.body\[330\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_96_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout906 net908 vssd1 vssd1 vccd1 vccd1 net906 sky130_fd_sc_hd__buf_2
X_09871_ _04840_ _04841_ _04842_ _04843_ vssd1 vssd1 vccd1 vccd1 _04844_ sky130_fd_sc_hd__or4_1
XANTENNA__19930__CLK clknet_leaf_51_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout917 net918 vssd1 vssd1 vccd1 vccd1 net917 sky130_fd_sc_hd__buf_4
Xfanout928 net929 vssd1 vssd1 vccd1 vccd1 net928 sky130_fd_sc_hd__buf_4
Xfanout939 net940 vssd1 vssd1 vccd1 vccd1 net939 sky130_fd_sc_hd__buf_4
XANTENNA__10025__B net1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12521__A net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10730__A2 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout182_A net183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11137__A net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10041__A net1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16749__A2 net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09884__B1 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09830__A net1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11691__B1 net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1091_A net1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout447_A net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13352__A _07519_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13432__A1 net236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09305_ sound_gen.osc1.count\[5\] sound_gen.osc1.count\[4\] _04323_ vssd1 vssd1 vccd1
+ vccd1 _04325_ sky130_fd_sc_hd__and3_1
XFILLER_0_130_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15709__B1 _01629_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13071__B _07639_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_135_4440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17759__A net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_135_4451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout614_A net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout235_X net235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1356_A net1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18371__A1 net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_4304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17111__X _02790_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09236_ net969 vssd1 vssd1 vccd1 vccd1 _04261_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_131_4315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_131_4326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17478__B net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_20_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_17_Right_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_40_1532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_255 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout402_X net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09167_ ag2.body\[527\] vssd1 vssd1 vccd1 vccd1 _04192_ sky130_fd_sc_hd__inv_2
XFILLER_0_126_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1144_X net1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11746__A1 net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_3_0_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09098_ ag2.body\[349\] vssd1 vssd1 vccd1 vccd1 _04123_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout983_A net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20327_ clknet_leaf_105_clk sound_gen.osc1.timer_nxt\[12\] _00004_ vssd1 vssd1 vccd1
+ vccd1 sound_gen.osc1.timer\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_102_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16602__S net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13499__A1 net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1311_X net1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10216__A net1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_4244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold960 _00663_ vssd1 vssd1 vccd1 vccd1 net2522 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_4255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold971 control.body\[910\] vssd1 vssd1 vccd1 vccd1 net2533 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout95_A net100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1552 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_129_4266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11060_ _06029_ _06030_ _06031_ _06032_ vssd1 vssd1 vccd1 vccd1 _06033_ sky130_fd_sc_hd__and4_1
Xhold982 control.body\[891\] vssd1 vssd1 vccd1 vccd1 net2544 sky130_fd_sc_hd__dlygate4sd3_1
X_20258_ clknet_leaf_43_clk _01202_ net1379 vssd1 vssd1 vccd1 vccd1 ag2.body\[0\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_101_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_99_1620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_38_1472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold993 _00312_ vssd1 vssd1 vccd1 vccd1 net2555 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_53_1926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout771_X net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_1494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18102__B _03683_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout869_X net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12171__A1 net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10011_ _04433_ _04791_ vssd1 vssd1 vccd1 vccd1 _04984_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_34_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_1506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_34_1358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09724__B net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20189_ clknet_leaf_88_clk _01133_ net1459 vssd1 vssd1 vccd1 vccd1 ag2.body\[203\]
+ sky130_fd_sc_hd__dfrtp_4
XPHY_EDGE_ROW_26_Right_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_34_1369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10721__A2 net1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13246__B net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_4_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15660__A2 net144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_103_clk_X clknet_leaf_103_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14750_ _08908_ _08909_ _08910_ vssd1 vssd1 vccd1 vccd1 _08911_ sky130_fd_sc_hd__or3b_1
XANTENNA__19899__RESET_B net1464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout50_X net50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11962_ img_gen.tracker.frame\[496\] net599 net583 img_gen.tracker.frame\[502\] _06933_
+ vssd1 vssd1 vccd1 vccd1 _06934_ sky130_fd_sc_hd__o221a_1
XANTENNA__17937__A1 net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_1214 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13701_ track.highScore\[2\] _04424_ _04637_ vssd1 vssd1 vccd1 vccd1 _08042_ sky130_fd_sc_hd__or3b_1
X_10913_ ag2.body\[458\] net1175 vssd1 vssd1 vccd1 vccd1 _05886_ sky130_fd_sc_hd__xnor2_1
XANTENNA__15461__B net63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14681_ _08837_ _08838_ _08839_ _08841_ vssd1 vssd1 vccd1 vccd1 _08842_ sky130_fd_sc_hd__a211o_1
XANTENNA__11682__B1 net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11893_ img_gen.tracker.frame\[73\] img_gen.tracker.frame\[76\] img_gen.tracker.frame\[79\]
+ img_gen.tracker.frame\[82\] net1216 net1190 vssd1 vssd1 vccd1 vccd1 _06865_ sky130_fd_sc_hd__mux4_1
XANTENNA__10886__A net1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16420_ obsg2.obstacleArray\[116\] obsg2.obstacleArray\[117\] obsg2.obstacleArray\[118\]
+ obsg2.obstacleArray\[119\] net455 net398 vssd1 vssd1 vccd1 vccd1 _02099_ sky130_fd_sc_hd__mux4_1
X_13632_ control.divider.count\[10\] control.divider.count\[9\] _07990_ control.divider.count\[11\]
+ vssd1 vssd1 vccd1 vccd1 _07996_ sky130_fd_sc_hd__a31o_1
X_10844_ ag2.body\[41\] net777 net767 ag2.body\[43\] vssd1 vssd1 vccd1 vccd1 _05817_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__13423__A1 net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14620__B1 ag2.body\[63\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_118_clk_X clknet_leaf_118_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16351_ _01930_ _01979_ _01996_ _02029_ vssd1 vssd1 vccd1 vccd1 _02030_ sky130_fd_sc_hd__a31o_1
XANTENNA__18558__CLK clknet_leaf_132_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13563_ _07933_ _07938_ vssd1 vssd1 vccd1 vccd1 _07942_ sky130_fd_sc_hd__and2_1
XFILLER_0_41_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10775_ ag2.body\[220\] net1140 vssd1 vssd1 vccd1 vccd1 _05748_ sky130_fd_sc_hd__xor2_1
XFILLER_0_137_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_35_Right_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19803__CLK clknet_leaf_124_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17165__A2 net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15302_ net2644 net78 _01586_ control.body\[721\] vssd1 vssd1 vccd1 vccd1 _00603_
+ sky130_fd_sc_hd__a22o_1
X_19070_ clknet_leaf_29_clk img_gen.tracker.next_frame\[508\] net1338 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[508\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__11985__B2 net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12514_ net387 net339 _07453_ vssd1 vssd1 vccd1 vccd1 _07454_ sky130_fd_sc_hd__or3_1
X_16282_ obsg2.obstacleArray\[20\] obsg2.obstacleArray\[21\] net412 vssd1 vssd1 vccd1
+ vccd1 _01961_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_114_3801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_3277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13494_ net276 _07908_ _07909_ net2051 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[542\]
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_97_3288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16912__A2 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18021_ _03541_ _03585_ vssd1 vssd1 vccd1 vccd1 _03630_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_114_3812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15233_ control.body\[797\] net96 _01577_ net2216 vssd1 vssd1 vccd1 vccd1 _00543_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_81_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12445_ _07355_ _07405_ _07403_ _07400_ vssd1 vssd1 vccd1 vccd1 _07406_ sky130_fd_sc_hd__o211ai_1
XANTENNA__16125__B1 net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15164_ _06182_ net63 vssd1 vssd1 vccd1 vccd1 _01570_ sky130_fd_sc_hd__and2_2
XFILLER_0_129_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12376_ img_gen.updater.commands.count\[14\] img_gen.updater.commands.count\[15\]
+ img_gen.updater.commands.count\[13\] _07340_ vssd1 vssd1 vccd1 vccd1 _07341_ sky130_fd_sc_hd__or4_1
XFILLER_0_50_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14115_ net832 ag2.body\[569\] ag2.body\[575\] net791 _08275_ vssd1 vssd1 vccd1 vccd1
+ _08276_ sky130_fd_sc_hd__a221o_1
XFILLER_0_132_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11327_ _06292_ _06294_ _06299_ vssd1 vssd1 vccd1 vccd1 _06300_ sky130_fd_sc_hd__or3_1
X_19972_ clknet_leaf_62_clk _00916_ net1470 vssd1 vssd1 vccd1 vccd1 ag2.body\[418\]
+ sky130_fd_sc_hd__dfrtp_4
X_15095_ control.body\[913\] net147 _01563_ net2093 vssd1 vssd1 vccd1 vccd1 _00419_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__10126__A net1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14821__A net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14046_ net1014 ag2.body\[191\] vssd1 vssd1 vccd1 vccd1 _08207_ sky130_fd_sc_hd__xnor2_1
X_18923_ clknet_leaf_140_clk img_gen.tracker.next_frame\[361\] net1290 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[361\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11258_ net1228 control.body\[768\] vssd1 vssd1 vccd1 vccd1 _06231_ sky130_fd_sc_hd__xor2_1
XPHY_EDGE_ROW_44_Right_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_108_3605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_3616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09563__C1 _04484_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10209_ net1230 control.body\[992\] vssd1 vssd1 vccd1 vccd1 _05182_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_108_3627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09634__B net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18854_ clknet_leaf_18_clk img_gen.tracker.next_frame\[292\] net1319 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[292\] sky130_fd_sc_hd__dfrtp_1
X_11189_ _04055_ net1209 net749 ag2.body\[182\] _06157_ vssd1 vssd1 vccd1 vccd1 _06162_
+ sky130_fd_sc_hd__a221o_1
X_17805_ net223 _08110_ net663 vssd1 vssd1 vccd1 vccd1 _03474_ sky130_fd_sc_hd__o21a_1
X_15997_ net870 net861 vssd1 vssd1 vccd1 vccd1 _01676_ sky130_fd_sc_hd__xnor2_2
X_18785_ clknet_leaf_12_clk img_gen.tracker.next_frame\[223\] net1285 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[223\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_136_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15651__A2 net139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17736_ _03340_ _03344_ _02703_ _03206_ vssd1 vssd1 vccd1 vccd1 _03415_ sky130_fd_sc_hd__o211a_2
X_14948_ net893 _04634_ net65 vssd1 vssd1 vccd1 vccd1 _01546_ sky130_fd_sc_hd__and3_2
XANTENNA__13662__A1 net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_2812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_82_2823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09650__A net1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17667_ ag2.body\[451\] net851 vssd1 vssd1 vccd1 vccd1 _03346_ sky130_fd_sc_hd__nand2_1
XFILLER_0_106_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_2834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14879_ net2374 net178 _01538_ control.body\[1098\] vssd1 vssd1 vccd1 vccd1 _00228_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_67_2380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14268__A net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_63_2233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19406_ clknet_leaf_103_clk net2385 net1427 vssd1 vssd1 vccd1 vccd1 control.body\[988\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_63_2244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16618_ obsg2.obstacleArray\[46\] net441 vssd1 vssd1 vccd1 vccd1 _02297_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_63_2255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17598_ ag2.body\[423\] net931 vssd1 vssd1 vccd1 vccd1 _03277_ sky130_fd_sc_hd__xor2_1
XFILLER_0_106_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13414__A1 net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_53_Right_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16549_ net463 _02220_ vssd1 vssd1 vccd1 vccd1 _02228_ sky130_fd_sc_hd__xnor2_4
X_19337_ clknet_leaf_103_clk net2180 net1431 vssd1 vssd1 vccd1 vccd1 control.body\[1063\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11404__B net1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19268_ clknet_leaf_71_clk _00212_ net1503 vssd1 vssd1 vccd1 vccd1 ag2.body\[131\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__17298__B net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14715__B ag2.body\[339\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09021_ ag2.body\[155\] vssd1 vssd1 vccd1 vccd1 _04046_ sky130_fd_sc_hd__inv_2
XFILLER_0_115_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18219_ obsg2.obstacleArray\[106\] _03748_ net524 vssd1 vssd1 vccd1 vccd1 _01357_
+ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_76_2627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19199_ clknet_leaf_89_clk _00143_ net1455 vssd1 vssd1 vccd1 vccd1 ag2.body\[62\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_14_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_2638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20056__RESET_B net1504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_2649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11420__A net1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold201 img_gen.tracker.frame\[253\] vssd1 vssd1 vccd1 vccd1 net1763 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_2048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold212 img_gen.tracker.frame\[254\] vssd1 vssd1 vccd1 vccd1 net1774 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_2059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold223 img_gen.tracker.frame\[85\] vssd1 vssd1 vccd1 vccd1 net1785 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold234 img_gen.tracker.frame\[92\] vssd1 vssd1 vccd1 vccd1 net1796 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold245 img_gen.tracker.frame\[409\] vssd1 vssd1 vccd1 vccd1 net1807 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14731__A net993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold256 img_gen.tracker.frame\[148\] vssd1 vssd1 vccd1 vccd1 net1818 sky130_fd_sc_hd__dlygate4sd3_1
Xhold267 img_gen.tracker.frame\[546\] vssd1 vssd1 vccd1 vccd1 net1829 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_62_Right_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold278 img_gen.tracker.frame\[293\] vssd1 vssd1 vccd1 vccd1 net1840 sky130_fd_sc_hd__dlygate4sd3_1
X_20112_ clknet_leaf_80_clk _01056_ net1487 vssd1 vssd1 vccd1 vccd1 ag2.body\[286\]
+ sky130_fd_sc_hd__dfrtp_4
X_09923_ _04891_ _04893_ _04895_ vssd1 vssd1 vccd1 vccd1 _04896_ sky130_fd_sc_hd__or3_1
XANTENNA__09825__A net1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout703 net704 vssd1 vssd1 vccd1 vccd1 net703 sky130_fd_sc_hd__clkbuf_4
Xhold289 img_gen.tracker.frame\[272\] vssd1 vssd1 vccd1 vccd1 net1851 sky130_fd_sc_hd__dlygate4sd3_1
Xfanout714 _04266_ vssd1 vssd1 vccd1 vccd1 net714 sky130_fd_sc_hd__clkbuf_8
XANTENNA__12153__A1 net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16419__A1 net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout725 _04264_ vssd1 vssd1 vccd1 vccd1 net725 sky130_fd_sc_hd__buf_4
XANTENNA_fanout397_A net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20043_ clknet_leaf_68_clk _00987_ net1495 vssd1 vssd1 vccd1 vccd1 ag2.body\[345\]
+ sky130_fd_sc_hd__dfrtp_4
Xfanout736 _04263_ vssd1 vssd1 vccd1 vccd1 net736 sky130_fd_sc_hd__buf_2
XANTENNA__13347__A net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09854_ net1230 control.body\[968\] vssd1 vssd1 vccd1 vccd1 _04827_ sky130_fd_sc_hd__xnor2_1
Xfanout747 _04234_ vssd1 vssd1 vccd1 vccd1 net747 sky130_fd_sc_hd__buf_4
Xfanout758 net766 vssd1 vssd1 vccd1 vccd1 net758 sky130_fd_sc_hd__buf_4
XANTENNA_fanout1104_A net1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout769 net770 vssd1 vssd1 vccd1 vccd1 net769 sky130_fd_sc_hd__clkbuf_4
XANTENNA__17711__S0 net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17761__B _02790_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13066__B _07726_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09785_ net917 net913 net909 vssd1 vssd1 vccd1 vccd1 _04758_ sky130_fd_sc_hd__a21o_4
XANTENNA_fanout564_A net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_72_clk_A clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout731_A _04263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout352_X net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_137_4502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout829_A net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1473_A net1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17395__A2 net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_71_Right_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1094_X net1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19826__CLK clknet_leaf_124_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_137_4513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13082__A net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19239__RESET_B net1480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_90 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_1741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_42_1605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout617_X net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_87_clk_A clknet_4_12__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18850__CLK clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10560_ net1228 ag2.body\[512\] vssd1 vssd1 vccd1 vccd1 _05533_ sky130_fd_sc_hd__and2b_1
XFILLER_0_107_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_23_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_130_clk_A clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09219_ control.body\[858\] vssd1 vssd1 vccd1 vccd1 _04244_ sky130_fd_sc_hd__inv_2
X_10491_ ag2.body\[550\] net1084 vssd1 vssd1 vccd1 vccd1 _05464_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_134_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_92_3130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_1630 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_3141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11330__A net1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12230_ _07198_ _07199_ vssd1 vssd1 vccd1 vccd1 _07200_ sky130_fd_sc_hd__nand2_1
XANTENNA_clkbuf_leaf_10_clk_A clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout986_X net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_15_Left_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16658__A1 net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_80_Right_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12392__A1 net1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12161_ img_gen.tracker.frame\[387\] net601 net585 img_gen.tracker.frame\[393\] _07132_
+ vssd1 vssd1 vccd1 vccd1 _07133_ sky130_fd_sc_hd__o221a_1
XANTENNA__16332__S net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14641__A net1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18113__A net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_145_clk_A clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_1409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11112_ net765 control.body\[1100\] control.body\[1101\] net756 vssd1 vssd1 vccd1
+ vccd1 _06085_ sky130_fd_sc_hd__o22a_1
X_12092_ net566 _07060_ _07063_ net470 vssd1 vssd1 vccd1 vccd1 _07064_ sky130_fd_sc_hd__o211a_1
Xhold790 _00270_ vssd1 vssd1 vccd1 vccd1 net2352 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_25_clk_A clknet_4_4__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15920_ _05921_ net57 vssd1 vssd1 vccd1 vccd1 _01654_ sky130_fd_sc_hd__nor2_2
XANTENNA__17952__A net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15881__A2 net192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11043_ _05452_ net477 _06015_ _04634_ vssd1 vssd1 vccd1 vccd1 _06016_ sky130_fd_sc_hd__a22o_1
XFILLER_0_99_1461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19356__CLK clknet_leaf_102_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15851_ ag2.body\[243\] net175 _01645_ ag2.body\[235\] vssd1 vssd1 vccd1 vccd1 _01093_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__17671__B net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14802_ net838 ag2.body\[289\] ag2.body\[295\] net795 vssd1 vssd1 vccd1 vccd1 _01473_
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_99_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15782_ ag2.body\[309\] net209 _01638_ ag2.body\[301\] vssd1 vssd1 vccd1 vccd1 _01031_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_73_1601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18570_ clknet_leaf_14_clk img_gen.tracker.next_frame\[8\] net1278 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[8\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__20333__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12994_ img_gen.tracker.frame\[259\] net645 vssd1 vssd1 vccd1 vccd1 _07693_ sky130_fd_sc_hd__and2_1
XFILLER_0_98_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_24_Left_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14733_ net1003 _04026_ ag2.body\[115\] net821 vssd1 vssd1 vccd1 vccd1 _08894_ sky130_fd_sc_hd__a22o_1
X_17521_ ag2.body\[487\] net929 vssd1 vssd1 vccd1 vccd1 _03200_ sky130_fd_sc_hd__xor2_1
XANTENNA__15191__B net58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11945_ img_gen.tracker.frame\[133\] net618 net572 _06916_ vssd1 vssd1 vccd1 vccd1
+ _06917_ sky130_fd_sc_hd__o211a_1
XFILLER_0_118_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14088__A net1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17452_ _04154_ net861 net703 ag2.body\[437\] vssd1 vssd1 vccd1 vccd1 _03131_ sky130_fd_sc_hd__o22a_1
XFILLER_0_129_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11505__A net1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14664_ net984 ag2.body\[522\] vssd1 vssd1 vccd1 vccd1 _08825_ sky130_fd_sc_hd__xor2_1
X_11876_ img_gen.tracker.frame\[253\] net615 net543 img_gen.tracker.frame\[259\] _06847_
+ vssd1 vssd1 vccd1 vccd1 _06848_ sky130_fd_sc_hd__o221a_1
XFILLER_0_52_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_99_3328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16403_ _02080_ _02081_ net403 vssd1 vssd1 vccd1 vccd1 _02082_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_99_3339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13615_ control.divider.count\[5\] control.divider.count\[4\] _07958_ vssd1 vssd1
+ vccd1 vccd1 _07985_ sky130_fd_sc_hd__and3_1
X_10827_ ag2.body\[310\] net1090 vssd1 vssd1 vccd1 vccd1 _05800_ sky130_fd_sc_hd__xor2_1
X_17383_ ag2.body\[494\] net942 vssd1 vssd1 vccd1 vccd1 _03062_ sky130_fd_sc_hd__nand2_1
X_14595_ net993 ag2.body\[305\] vssd1 vssd1 vccd1 vccd1 _08756_ sky130_fd_sc_hd__xor2_1
XFILLER_0_131_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11958__A1 net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16334_ obsg2.obstacleArray\[86\] net411 vssd1 vssd1 vccd1 vccd1 _02013_ sky130_fd_sc_hd__or2_1
XFILLER_0_82_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19122_ clknet_leaf_141_clk img_gen.tracker.next_frame\[560\] net1262 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[560\] sky130_fd_sc_hd__dfrtp_1
X_13546_ net2132 net659 _07929_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[574\]
+ sky130_fd_sc_hd__and3_1
X_10758_ net1179 control.body\[890\] vssd1 vssd1 vccd1 vccd1 _05731_ sky130_fd_sc_hd__or2_1
X_19053_ clknet_leaf_10_clk img_gen.tracker.next_frame\[491\] net1273 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[491\] sky130_fd_sc_hd__dfrtp_1
X_16265_ obsg2.obstacleArray\[49\] net413 _01943_ net418 vssd1 vssd1 vccd1 vccd1 _01944_
+ sky130_fd_sc_hd__o211a_1
X_13477_ net230 _07902_ _07903_ net1848 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[531\]
+ sky130_fd_sc_hd__a22o_1
X_10689_ ag2.body\[148\] net1141 vssd1 vssd1 vccd1 vccd1 _05662_ sky130_fd_sc_hd__xor2_1
XPHY_EDGE_ROW_33_Left_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18004_ net46 _03617_ vssd1 vssd1 vccd1 vccd1 _03618_ sky130_fd_sc_hd__nor2_1
X_15216_ net2646 net92 _01575_ net2341 vssd1 vssd1 vccd1 vccd1 _00528_ sky130_fd_sc_hd__a22o_1
XFILLER_0_125_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12428_ net1094 net1045 vssd1 vssd1 vccd1 vccd1 _07390_ sky130_fd_sc_hd__or2_1
X_16196_ obsg2.obstacleArray\[60\] obsg2.obstacleArray\[61\] net424 vssd1 vssd1 vccd1
+ vccd1 _01875_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_1185 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11186__A2 net1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_1627 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_2502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15147_ control.body\[864\] net105 _01568_ net2276 vssd1 vssd1 vccd1 vccd1 _00466_
+ sky130_fd_sc_hd__a22o_1
X_12359_ _06631_ _06635_ _07251_ _07292_ _07253_ vssd1 vssd1 vccd1 vccd1 _07326_ sky130_fd_sc_hd__a41o_1
XANTENNA__18023__A net45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1168 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19955_ clknet_leaf_62_clk _00899_ net1381 vssd1 vssd1 vccd1 vccd1 ag2.body\[433\]
+ sky130_fd_sc_hd__dfrtp_4
X_15078_ net2623 net147 _01561_ net2269 vssd1 vssd1 vccd1 vccd1 _00404_ sky130_fd_sc_hd__a22o_1
XFILLER_0_10_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11569__S0 net1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14029_ net811 ag2.body\[28\] _03985_ net1007 _08185_ vssd1 vssd1 vccd1 vccd1 _08190_
+ sky130_fd_sc_hd__o221a_1
X_18906_ clknet_leaf_144_clk img_gen.tracker.next_frame\[344\] net1251 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[344\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_103_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12071__A net1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19886_ clknet_leaf_85_clk _00830_ net1462 vssd1 vssd1 vccd1 vccd1 ag2.body\[508\]
+ sky130_fd_sc_hd__dfrtp_4
X_18837_ clknet_leaf_142_clk img_gen.tracker.next_frame\[275\] net1260 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[275\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_69_2420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_2431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18723__CLK clknet_leaf_142_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_42_Left_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19849__CLK clknet_leaf_93_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_2442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09570_ _04063_ net1208 net1184 _04064_ _04542_ vssd1 vssd1 vccd1 vccd1 _04543_ sky130_fd_sc_hd__a221o_1
X_18768_ clknet_leaf_16_clk img_gen.tracker.next_frame\[206\] net1321 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[206\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_65_2306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14832__B1 _08623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_65_2317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17719_ obsg2.obstacleArray\[130\] obsg2.obstacleArray\[131\] net427 vssd1 vssd1
+ vccd1 vccd1 _03398_ sky130_fd_sc_hd__mux2_1
XFILLER_0_136_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18699_ clknet_leaf_10_clk img_gen.tracker.next_frame\[137\] net1274 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[137\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_114_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11415__A net1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_19_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18873__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19999__CLK clknet_leaf_66_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16925__B net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14726__A net1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14060__A1 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18326__A1 _04944_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17129__A2 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14060__B2 net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_520 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20592_ net1524 vssd1 vssd1 vccd1 vccd1 gpio_oeb[4] sky130_fd_sc_hd__buf_2
XFILLER_0_73_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_1663 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_51_Left_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout312_A net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1054_A net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09004_ ag2.body\[121\] vssd1 vssd1 vccd1 vccd1 _04029_ sky130_fd_sc_hd__inv_2
XFILLER_0_103_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17756__B _03434_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout100_X net100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1221_A ag2.y\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17301__A2 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09555__A net1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout500 net501 vssd1 vssd1 vccd1 vccd1 net500 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout681_A _04393_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout511 net515 vssd1 vssd1 vccd1 vccd1 net511 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout779_A net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1509 net1511 vssd1 vssd1 vccd1 vccd1 net1509 sky130_fd_sc_hd__clkbuf_2
X_09906_ ag2.body\[130\] net1188 vssd1 vssd1 vccd1 vccd1 _04879_ sky130_fd_sc_hd__nand2_1
XANTENNA__11149__X _06122_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout522 net523 vssd1 vssd1 vccd1 vccd1 net522 sky130_fd_sc_hd__buf_2
XFILLER_0_22_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13077__A net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout533 net534 vssd1 vssd1 vccd1 vccd1 net533 sky130_fd_sc_hd__buf_2
XFILLER_0_96_1601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1107_X net1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout544 net545 vssd1 vssd1 vccd1 vccd1 net544 sky130_fd_sc_hd__clkbuf_4
Xfanout555 _06651_ vssd1 vssd1 vccd1 vccd1 net555 sky130_fd_sc_hd__buf_4
XANTENNA__16499__S0 net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20026_ clknet_leaf_67_clk _00970_ net1473 vssd1 vssd1 vccd1 vccd1 ag2.body\[360\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_77_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout566 net567 vssd1 vssd1 vccd1 vccd1 net566 sky130_fd_sc_hd__clkbuf_4
X_09837_ _04806_ _04807_ _04808_ _04809_ vssd1 vssd1 vccd1 vccd1 _04810_ sky130_fd_sc_hd__a22o_1
Xfanout577 _06649_ vssd1 vssd1 vccd1 vccd1 net577 sky130_fd_sc_hd__clkbuf_4
Xfanout588 net589 vssd1 vssd1 vccd1 vccd1 net588 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_119_1310 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout946_A net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout599 net602 vssd1 vssd1 vccd1 vccd1 net599 sky130_fd_sc_hd__buf_2
XANTENNA_fanout567_X net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16273__C1 net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09768_ ag2.body\[238\] net1085 vssd1 vssd1 vccd1 vccd1 _04741_ sky130_fd_sc_hd__xor2_1
XFILLER_0_119_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout58_A net59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13524__B _07807_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout734_X net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09699_ ag2.body\[67\] net1162 vssd1 vssd1 vccd1 vccd1 _04672_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_29_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_1364 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11730_ img_gen.tracker.frame\[215\] net591 _06649_ _06701_ vssd1 vssd1 vccd1 vccd1
+ _06702_ sky130_fd_sc_hd__o211a_1
XFILLER_0_90_1277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16040__A2 net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16835__B net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11661_ _06612_ _06633_ _06623_ _06559_ vssd1 vssd1 vccd1 vccd1 _06634_ sky130_fd_sc_hd__and4bb_2
XFILLER_0_37_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout901_X net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14051__A1 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12708__X _07558_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18108__A net44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14051__B2 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13400_ net283 net312 _07551_ _07872_ net1646 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[485\]
+ sky130_fd_sc_hd__a32o_1
X_10612_ _05581_ _05582_ _05583_ _05584_ vssd1 vssd1 vccd1 vccd1 _05585_ sky130_fd_sc_hd__or4_1
X_14380_ net834 ag2.body\[417\] ag2.body\[423\] net792 _08538_ vssd1 vssd1 vccd1 vccd1
+ _08541_ sky130_fd_sc_hd__o221a_1
XANTENNA__12062__B1 net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_94_3203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11592_ _06563_ _06564_ net507 vssd1 vssd1 vccd1 vccd1 _06565_ sky130_fd_sc_hd__mux2_1
XFILLER_0_92_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13331_ net275 _07844_ _07845_ net1758 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[443\]
+ sky130_fd_sc_hd__a22o_1
X_10543_ ag2.body\[230\] net1085 vssd1 vssd1 vccd1 vccd1 _05516_ sky130_fd_sc_hd__or2_1
XFILLER_0_52_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09449__B net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17540__A2 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16050_ net463 _01727_ vssd1 vssd1 vccd1 vccd1 _01729_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_106_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13262_ net282 _07817_ _07818_ net1856 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[401\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__17666__B net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10474_ _05443_ _05444_ _05445_ _05446_ vssd1 vssd1 vccd1 vccd1 _05447_ sky130_fd_sc_hd__or4_1
XFILLER_0_121_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15001_ control.body\[1007\] net153 _01551_ control.body\[999\] vssd1 vssd1 vccd1
+ vccd1 _00337_ sky130_fd_sc_hd__a22o_1
XANTENNA__17828__A0 net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12213_ img_gen.control.current\[1\] img_gen.control.current\[0\] _07182_ _07184_
+ _07178_ vssd1 vssd1 vccd1 vccd1 img_gen.control.next\[0\] sky130_fd_sc_hd__o32a_1
XFILLER_0_62_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14371__A net1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13193_ img_gen.tracker.frame\[364\] net658 vssd1 vssd1 vccd1 vccd1 _07787_ sky130_fd_sc_hd__and2_1
XFILLER_0_102_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12144_ img_gen.tracker.frame\[507\] net599 net544 img_gen.tracker.frame\[510\] vssd1
+ vssd1 vccd1 vccd1 _07116_ sky130_fd_sc_hd__o22a_1
XFILLER_0_62_1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16500__B1 _02075_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_88_3007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_88_3018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17682__A ag2.body\[478\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19740_ clknet_leaf_129_clk _00684_ net1304 vssd1 vssd1 vccd1 vccd1 control.body\[650\]
+ sky130_fd_sc_hd__dfrtp_1
X_16952_ _02623_ _02624_ _02627_ _02630_ vssd1 vssd1 vccd1 vccd1 _02631_ sky130_fd_sc_hd__or4_1
X_12075_ img_gen.tracker.frame\[123\] net611 net594 img_gen.tracker.frame\[129\] _07046_
+ vssd1 vssd1 vccd1 vccd1 _07047_ sky130_fd_sc_hd__a221o_1
XFILLER_0_104_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10404__A net1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15903_ ag2.body\[193\] net129 _01651_ ag2.body\[185\] vssd1 vssd1 vccd1 vccd1 _01139_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_40_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11026_ _05992_ _05993_ _05998_ _05991_ _05990_ vssd1 vssd1 vccd1 vccd1 _05999_ sky130_fd_sc_hd__a2111oi_2
X_19671_ clknet_leaf_135_clk _00615_ net1302 vssd1 vssd1 vccd1 vccd1 control.body\[725\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11876__B1 net543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16883_ ag2.body\[17\] net730 net688 ag2.body\[23\] vssd1 vssd1 vccd1 vccd1 _02562_
+ sky130_fd_sc_hd__a22o_1
X_18622_ clknet_leaf_3_clk img_gen.tracker.next_frame\[60\] net1248 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[60\] sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_4_2__f_clk_A clknet_3_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09912__B net1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15834_ ag2.body\[260\] net204 net49 ag2.body\[252\] vssd1 vssd1 vccd1 vccd1 _01078_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_63_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18005__B1 net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18553_ clknet_leaf_37_clk _00079_ net1349 vssd1 vssd1 vccd1 vccd1 control.divider.fsm.current_mode\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_15765_ ag2.body\[326\] net216 _01636_ ag2.body\[318\] vssd1 vssd1 vccd1 vccd1 _01016_
+ sky130_fd_sc_hd__a22o_1
X_12977_ net2035 net645 _07684_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[250\]
+ sky130_fd_sc_hd__and3_1
XANTENNA__14290__A1 net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14225__A1_N net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14290__B2 net806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17504_ ag2.body\[233\] net735 net854 _04072_ _03182_ vssd1 vssd1 vccd1 vccd1 _03183_
+ sky130_fd_sc_hd__a221o_1
X_14716_ net978 ag2.body\[339\] vssd1 vssd1 vccd1 vccd1 _08877_ sky130_fd_sc_hd__or2_1
XFILLER_0_87_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_16_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11928_ _06895_ _06896_ _06897_ _06899_ vssd1 vssd1 vccd1 vccd1 _06900_ sky130_fd_sc_hd__o31a_1
XANTENNA__16567__B1 net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15696_ ag2.body\[377\] net137 _01628_ ag2.body\[369\] vssd1 vssd1 vccd1 vccd1 _00955_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_16_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18484_ net1515 net1509 vssd1 vssd1 vccd1 vccd1 _00015_ sky130_fd_sc_hd__or2_1
XFILLER_0_118_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17435_ ag2.body\[146\] net865 vssd1 vssd1 vccd1 vccd1 _03114_ sky130_fd_sc_hd__xor2_1
X_14647_ net991 ag2.body\[513\] vssd1 vssd1 vccd1 vccd1 _08808_ sky130_fd_sc_hd__xor2_1
XANTENNA__14042__A1 net1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11859_ net567 _06827_ _06828_ _06830_ vssd1 vssd1 vccd1 vccd1 _06831_ sky130_fd_sc_hd__a22o_1
XFILLER_0_28_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14546__A net975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14042__B2 net1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13450__A _07581_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_18 _08509_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17366_ _03020_ _03023_ _03042_ _03044_ vssd1 vssd1 vccd1 vccd1 _03045_ sky130_fd_sc_hd__a211o_1
XANTENNA_29 _03442_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14578_ net802 ag2.body\[494\] _04179_ net1009 vssd1 vssd1 vccd1 vccd1 _08739_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__10793__B net1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20229__CLK clknet_leaf_66_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19105_ clknet_leaf_1_clk img_gen.tracker.next_frame\[543\] net1244 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[543\] sky130_fd_sc_hd__dfrtp_1
X_16317_ _01912_ _01990_ _01994_ _01995_ _01919_ vssd1 vssd1 vccd1 vccd1 _01996_ sky130_fd_sc_hd__a311o_1
XFILLER_0_6_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13529_ _07624_ _07807_ vssd1 vssd1 vccd1 vccd1 _07923_ sky130_fd_sc_hd__or2_1
XANTENNA__11800__B1 _06741_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17297_ ag2.body\[349\] net708 net694 ag2.body\[351\] _02975_ vssd1 vssd1 vccd1 vccd1
+ _02976_ sky130_fd_sc_hd__a221o_1
XFILLER_0_12_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14833__X _01504_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20056__Q ag2.body\[342\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16248_ _01912_ _01926_ _01919_ vssd1 vssd1 vccd1 vccd1 _01927_ sky130_fd_sc_hd__a21o_1
XANTENNA__09927__X _04900_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19036_ clknet_leaf_6_clk img_gen.tracker.next_frame\[474\] net1264 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[474\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__17576__B net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16179_ net373 _01857_ _01856_ net348 vssd1 vssd1 vccd1 vccd1 _01858_ sky130_fd_sc_hd__a211o_1
XFILLER_0_23_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11564__C1 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12513__B net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19938_ clknet_leaf_46_clk _00882_ net1375 vssd1 vssd1 vccd1 vccd1 ag2.body\[448\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_103_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19869_ clknet_leaf_95_clk _00813_ net1440 vssd1 vssd1 vccd1 vccd1 ag2.body\[523\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__10033__B net1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18200__B net40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09622_ net1148 control.body\[803\] vssd1 vssd1 vccd1 vccd1 _04595_ sky130_fd_sc_hd__xnor2_1
XANTENNA__19513__RESET_B net1403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1217 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16001__A net871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14805__B1 ag2.body\[290\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09553_ net1049 control.body\[727\] vssd1 vssd1 vccd1 vccd1 _04526_ sky130_fd_sc_hd__nand2_1
XANTENNA__14281__A1 net1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout262_A net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14281__B2 net809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_1549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09484_ _04449_ _04456_ _04451_ _04453_ vssd1 vssd1 vccd1 vccd1 _04457_ sky130_fd_sc_hd__or4b_1
XFILLER_0_17_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12796__A_N _07423_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16147__S net429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10984__A net1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout527_A net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1171_A net1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1269_A net1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18619__CLK clknet_leaf_144_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12044__B1 net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_1460 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1283 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11398__A2 _04425_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14743__X _08904_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10048__X _05021_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20575_ clknet_leaf_106_clk _01433_ _00039_ vssd1 vssd1 vccd1 vccd1 sound_gen.dac1.dacCount\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout315_X net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_13__f_clk_A clknet_3_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1057_X net1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1436_A net1442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14191__A net974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1224_X net1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10190_ ag2.body\[113\] net1212 vssd1 vssd1 vccd1 vccd1 _05163_ sky130_fd_sc_hd__xor2_1
XANTENNA__13519__B net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout684_X net684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1306 net1310 vssd1 vssd1 vccd1 vccd1 net1306 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__16610__S net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1317 net1324 vssd1 vssd1 vccd1 vccd1 net1317 sky130_fd_sc_hd__clkbuf_4
Xfanout1328 net1330 vssd1 vssd1 vccd1 vccd1 net1328 sky130_fd_sc_hd__clkbuf_4
Xfanout330 net331 vssd1 vssd1 vccd1 vccd1 net330 sky130_fd_sc_hd__buf_1
Xfanout1339 net1341 vssd1 vssd1 vccd1 vccd1 net1339 sky130_fd_sc_hd__clkbuf_4
Xfanout341 net342 vssd1 vssd1 vccd1 vccd1 net341 sky130_fd_sc_hd__clkbuf_4
Xfanout352 net354 vssd1 vssd1 vccd1 vccd1 net352 sky130_fd_sc_hd__buf_4
XFILLER_0_100_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18235__B1 net527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout851_X net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11858__B1 net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout374 net375 vssd1 vssd1 vccd1 vccd1 net374 sky130_fd_sc_hd__buf_4
XFILLER_0_96_1442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout949_X net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17589__A2 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout385 _06676_ vssd1 vssd1 vccd1 vccd1 net385 sky130_fd_sc_hd__buf_2
Xfanout396 _02216_ vssd1 vssd1 vccd1 vccd1 net396 sky130_fd_sc_hd__buf_4
X_12900_ _07649_ net267 _07647_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[208\]
+ sky130_fd_sc_hd__mux2_1
X_20009_ clknet_leaf_61_clk _00953_ net1468 vssd1 vssd1 vccd1 vccd1 ag2.body\[391\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__19254__RESET_B net1492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09732__B net1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13880_ ag2.body\[29\] net115 _08147_ ag2.body\[21\] vssd1 vssd1 vccd1 vccd1 _00110_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_92_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_hold739_A coll.badColl vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10878__B net1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12831_ net239 _07616_ _07617_ net1776 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[171\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12796__D net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09451__C net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15550_ _04416_ _04944_ net61 vssd1 vssd1 vccd1 vccd1 _01612_ sky130_fd_sc_hd__a21oi_4
X_12762_ net305 _07584_ vssd1 vssd1 vccd1 vccd1 _07585_ sky130_fd_sc_hd__nor2_1
XFILLER_0_9_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14501_ net983 _04087_ ag2.body\[263\] net795 _08659_ vssd1 vssd1 vccd1 vccd1 _08662_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_55_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11713_ img_gen.tracker.frame\[329\] net606 net551 img_gen.tracker.frame\[332\] _06684_
+ vssd1 vssd1 vccd1 vccd1 _06685_ sky130_fd_sc_hd__o221a_1
XFILLER_0_68_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15481_ ag2.body\[569\] net111 _01605_ ag2.body\[561\] vssd1 vssd1 vccd1 vccd1 _00763_
+ sky130_fd_sc_hd__a22o_1
X_12693_ net310 _07551_ net673 vssd1 vssd1 vccd1 vccd1 _07552_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_83_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14366__A net1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17220_ _04106_ net967 net707 ag2.body\[317\] vssd1 vssd1 vccd1 vccd1 _02899_ sky130_fd_sc_hd__o22a_1
X_14432_ _08586_ _08589_ _08591_ _08592_ vssd1 vssd1 vccd1 vccd1 _08593_ sky130_fd_sc_hd__or4_1
XFILLER_0_108_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11644_ obsg2.obstacleArray\[130\] obsg2.obstacleArray\[134\] net513 vssd1 vssd1
+ vccd1 vccd1 _06617_ sky130_fd_sc_hd__mux2_1
XANTENNA__12035__B1 net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19544__CLK clknet_leaf_118_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17151_ ag2.body\[612\] net958 vssd1 vssd1 vccd1 vccd1 _02830_ sky130_fd_sc_hd__xor2_1
X_14363_ net979 ag2.body\[602\] vssd1 vssd1 vccd1 vccd1 _08524_ sky130_fd_sc_hd__xnor2_1
XANTENNA__11502__B net1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11575_ obsg2.obstacleArray\[82\] net514 net507 vssd1 vssd1 vccd1 vccd1 _06548_ sky130_fd_sc_hd__o21a_1
X_16102_ obsg2.obstacleArray\[65\] net431 vssd1 vssd1 vccd1 vccd1 _01781_ sky130_fd_sc_hd__or2_1
XANTENNA__17513__A2 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13314_ net664 _07839_ vssd1 vssd1 vccd1 vccd1 _07840_ sky130_fd_sc_hd__nor2_1
XANTENNA__10061__A2 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17082_ ag2.body\[197\] net947 vssd1 vssd1 vccd1 vccd1 _02761_ sky130_fd_sc_hd__or2_1
X_10526_ net1229 control.body\[912\] vssd1 vssd1 vccd1 vccd1 _05499_ sky130_fd_sc_hd__xor2_1
XANTENNA__20521__CLK clknet_leaf_93_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16721__B1 net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14294_ net817 ag2.body\[475\] _04170_ net1025 _08450_ vssd1 vssd1 vccd1 vccd1 _08455_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_68_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16033_ _01680_ _01681_ vssd1 vssd1 vccd1 vccd1 _01712_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_106_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13245_ net283 net314 _07435_ _07810_ net1668 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[392\]
+ sky130_fd_sc_hd__a32o_1
XANTENNA__09907__B net1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10457_ ag2.body\[449\] net1198 vssd1 vssd1 vccd1 vccd1 _05430_ sky130_fd_sc_hd__xor2_1
XFILLER_0_27_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10349__B1 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12614__A net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11010__A1 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13176_ net231 _07778_ _07779_ net1918 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[354\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11010__B2 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10388_ net1205 control.body\[1057\] vssd1 vssd1 vccd1 vccd1 _05361_ sky130_fd_sc_hd__xor2_1
XANTENNA__16485__C1 net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11561__A2 net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12127_ _07095_ _07096_ _07098_ net558 vssd1 vssd1 vccd1 vccd1 _07099_ sky130_fd_sc_hd__a22o_1
X_17984_ net381 _01890_ net485 vssd1 vssd1 vccd1 vccd1 _03603_ sky130_fd_sc_hd__or3b_1
XFILLER_0_104_1475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16520__S _02057_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10134__A net1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13838__B2 net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09506__A2 net1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19723_ clknet_leaf_132_clk _00667_ net1303 vssd1 vssd1 vccd1 vccd1 control.body\[665\]
+ sky130_fd_sc_hd__dfrtp_1
X_12058_ img_gen.tracker.frame\[87\] net610 net555 img_gen.tracker.frame\[90\] _07029_
+ vssd1 vssd1 vccd1 vccd1 _07030_ sky130_fd_sc_hd__a221oi_2
X_16935_ ag2.body\[522\] net864 vssd1 vssd1 vccd1 vccd1 _02614_ sky130_fd_sc_hd__xor2_1
XFILLER_0_79_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13445__A _07578_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11009_ net750 control.body\[1086\] net895 vssd1 vssd1 vccd1 vccd1 _05982_ sky130_fd_sc_hd__o21a_1
X_19654_ clknet_leaf_133_clk _00598_ net1309 vssd1 vssd1 vccd1 vccd1 control.body\[740\]
+ sky130_fd_sc_hd__dfrtp_1
X_16866_ _02538_ _02544_ vssd1 vssd1 vccd1 vccd1 _02545_ sky130_fd_sc_hd__or2_1
XFILLER_0_88_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18605_ clknet_leaf_17_clk img_gen.tracker.next_frame\[43\] net1318 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[43\] sky130_fd_sc_hd__dfrtp_1
X_15817_ ag2.body\[276\] net205 _01642_ ag2.body\[268\] vssd1 vssd1 vccd1 vccd1 _01062_
+ sky130_fd_sc_hd__a22o_1
X_19585_ clknet_leaf_116_clk _00529_ net1385 vssd1 vssd1 vccd1 vccd1 control.body\[815\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14828__X _01499_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16797_ obsg2.obstacleArray\[134\] obsg2.obstacleArray\[135\] net457 vssd1 vssd1
+ vccd1 vccd1 _02476_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20511__RESET_B net1403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15460__B1 _01602_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18536_ clknet_leaf_136_clk _00062_ net1300 vssd1 vssd1 vccd1 vccd1 img_gen.updater.commands.count\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_15748_ ag2.body\[343\] net216 _01634_ ag2.body\[335\] vssd1 vssd1 vccd1 vccd1 _01001_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_5_1622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18467_ net969 net883 net871 vssd1 vssd1 vccd1 vccd1 _03954_ sky130_fd_sc_hd__a21o_1
XANTENNA__14015__A1 net999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15679_ ag2.body\[393\] net141 _01627_ ag2.body\[385\] vssd1 vssd1 vccd1 vccd1 _00939_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_114_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14015__B2 net1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12348__X _07315_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13180__A net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17418_ ag2.body\[285\] net707 net692 ag2.body\[287\] _03091_ vssd1 vssd1 vccd1 vccd1
+ _03097_ sky130_fd_sc_hd__a221o_1
XANTENNA__12026__B1 net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18398_ _03886_ _03887_ _03785_ vssd1 vssd1 vccd1 vccd1 _03888_ sky130_fd_sc_hd__o21ba_1
XANTENNA__12577__A1 net247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17349_ _03021_ _03022_ _03025_ _03027_ vssd1 vssd1 vccd1 vccd1 _03028_ sky130_fd_sc_hd__or4b_1
XANTENNA__18911__CLK clknet_leaf_142_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10309__A net1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17504__A2 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20360_ clknet_leaf_21_clk _00000_ net1361 vssd1 vssd1 vccd1 vccd1 obsg2.obsNeeded\[0\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_130_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19019_ clknet_leaf_6_clk img_gen.tracker.next_frame\[457\] net1264 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[457\] sky130_fd_sc_hd__dfrtp_1
X_20291_ clknet_leaf_37_clk control.divider.next_count\[12\] net1350 vssd1 vssd1 vccd1
+ vccd1 control.divider.count\[12\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_686 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11001__A1 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11001__B2 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08984_ ag2.body\[78\] vssd1 vssd1 vccd1 vccd1 _04009_ sky130_fd_sc_hd__inv_2
XANTENNA__16430__S net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10044__A net1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1017_A net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18217__B1 net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09833__A net1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19417__CLK clknet_leaf_105_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10979__A net1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11574__S net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10698__B net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09605_ net1195 control.body\[633\] vssd1 vssd1 vccd1 vccd1 _04578_ sky130_fd_sc_hd__xor2_1
XFILLER_0_39_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15451__B1 _01601_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout265_X net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1386_A net1404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09536_ net779 control.body\[1025\] control.body\[1027\] net769 _04504_ vssd1 vssd1
+ vccd1 vccd1 _04509_ sky130_fd_sc_hd__o221a_1
XFILLER_0_52_1323 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09467_ ag2.body\[377\] net778 net763 ag2.body\[380\] _04439_ vssd1 vssd1 vccd1 vccd1
+ _04440_ sky130_fd_sc_hd__a221o_1
XFILLER_0_94_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14186__A net1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout432_X net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16953__X _02632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout811_A net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15203__B1 _01574_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11162__X _06135_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12017__B1 net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20544__CLK clknet_leaf_105_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09398_ net2172 _04343_ net270 vssd1 vssd1 vccd1 vccd1 _04383_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_65_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11322__B net1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20627_ sound_gen.dac1.dacCount\[5\] vssd1 vssd1 vccd1 vccd1 net14 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_80_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_129_Right_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11360_ net774 control.body\[810\] control.body\[808\] net783 vssd1 vssd1 vccd1 vccd1
+ _06333_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__16703__B1 net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20558_ clknet_leaf_109_clk toggle1.nextBlinkToggle\[0\] net1416 vssd1 vssd1 vccd1
+ vccd1 net25 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_46_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout899_X net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11791__A2 net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10311_ _05273_ _05275_ _05276_ _05282_ vssd1 vssd1 vccd1 vccd1 _05284_ sky130_fd_sc_hd__or4_1
XFILLER_0_127_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11291_ net1062 control.body\[1111\] vssd1 vssd1 vccd1 vccd1 _06264_ sky130_fd_sc_hd__xor2_1
X_20489_ clknet_leaf_37_clk _01376_ net1353 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[125\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_104_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13030_ net283 _07708_ _07709_ net1653 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[278\]
+ sky130_fd_sc_hd__a22o_1
X_10242_ ag2.body\[324\] net1141 vssd1 vssd1 vccd1 vccd1 _05215_ sky130_fd_sc_hd__nand2_1
XANTENNA__09736__A2 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17944__B net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09446__C net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11543__A2 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12740__A1 net237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16340__S net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10173_ _05050_ _05088_ _05119_ _05145_ vssd1 vssd1 vccd1 vccd1 _05146_ sky130_fd_sc_hd__and4_1
Xfanout1103 net1106 vssd1 vssd1 vccd1 vccd1 net1103 sky130_fd_sc_hd__clkbuf_4
XANTENNA__18121__A net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1114 net1117 vssd1 vssd1 vccd1 vccd1 net1114 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10897__A4 _05075_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1125 net1126 vssd1 vssd1 vccd1 vccd1 net1125 sky130_fd_sc_hd__clkbuf_4
Xfanout1136 net1137 vssd1 vssd1 vccd1 vccd1 net1136 sky130_fd_sc_hd__clkbuf_4
Xfanout1147 net1156 vssd1 vssd1 vccd1 vccd1 net1147 sky130_fd_sc_hd__clkbuf_4
Xfanout1158 net1166 vssd1 vssd1 vccd1 vccd1 net1158 sky130_fd_sc_hd__buf_4
X_14981_ control.body\[1020\] net153 _01550_ net2537 vssd1 vssd1 vccd1 vccd1 _00318_
+ sky130_fd_sc_hd__a22o_1
Xfanout160 net161 vssd1 vssd1 vccd1 vccd1 net160 sky130_fd_sc_hd__buf_2
Xfanout171 net183 vssd1 vssd1 vccd1 vccd1 net171 sky130_fd_sc_hd__clkbuf_2
Xfanout1169 net1173 vssd1 vssd1 vccd1 vccd1 net1169 sky130_fd_sc_hd__buf_4
XANTENNA__11926__S0 net1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16720_ obsg2.obstacleArray\[104\] net491 net482 obsg2.obstacleArray\[105\] _02398_
+ vssd1 vssd1 vccd1 vccd1 _02399_ sky130_fd_sc_hd__a221o_1
Xfanout182 net183 vssd1 vssd1 vccd1 vccd1 net182 sky130_fd_sc_hd__clkbuf_2
Xfanout193 net194 vssd1 vssd1 vccd1 vccd1 net193 sky130_fd_sc_hd__buf_2
XANTENNA__09462__B net1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13932_ ag2.body\[75\] net193 _08153_ ag2.body\[67\] vssd1 vssd1 vccd1 vccd1 _00156_
+ sky130_fd_sc_hd__a22o_1
X_16651_ obsg2.obstacleArray\[7\] _02213_ net392 _02329_ vssd1 vssd1 vccd1 vccd1 _02330_
+ sky130_fd_sc_hd__o211a_1
X_13863_ net322 track.nextHighScore\[6\] _08136_ track.nextHighScore\[7\] vssd1 vssd1
+ vccd1 vccd1 _08137_ sky130_fd_sc_hd__a31o_1
XFILLER_0_57_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17024__X _02703_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15602_ ag2.body\[468\] net121 _01619_ net2511 vssd1 vssd1 vccd1 vccd1 _00870_ sky130_fd_sc_hd__a22o_1
XFILLER_0_97_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12814_ net239 _07608_ _07609_ net1831 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[162\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_9_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_3482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_762 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19370_ clknet_leaf_102_clk _00314_ net1436 vssd1 vssd1 vccd1 vccd1 control.body\[1016\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_104_3493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16582_ _01700_ _02207_ vssd1 vssd1 vccd1 vccd1 _02261_ sky130_fd_sc_hd__and2_1
X_13794_ _08095_ _08098_ _08100_ vssd1 vssd1 vccd1 vccd1 _00071_ sky130_fd_sc_hd__and3_1
XFILLER_0_9_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16295__B net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18321_ _03809_ _03812_ _03815_ _03791_ vssd1 vssd1 vccd1 vccd1 _03817_ sky130_fd_sc_hd__a31o_1
XFILLER_0_56_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12745_ net682 _07576_ vssd1 vssd1 vccd1 vccd1 _07577_ sky130_fd_sc_hd__nor2_1
XFILLER_0_35_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15533_ _05305_ net62 vssd1 vssd1 vccd1 vccd1 _01611_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_100_3368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1576 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_3379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18252_ _03693_ net35 vssd1 vssd1 vccd1 vccd1 _03765_ sky130_fd_sc_hd__nor2_1
XANTENNA__10282__A2 _05254_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15464_ ag2.body\[586\] net111 _01603_ ag2.body\[578\] vssd1 vssd1 vccd1 vccd1 _00748_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__15745__A1 ag2.body\[340\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12676_ net680 _07543_ vssd1 vssd1 vccd1 vccd1 _07544_ sky130_fd_sc_hd__nor2_1
XFILLER_0_38_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12559__A1 net226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17203_ ag2.body\[181\] net703 _02876_ _02877_ _02881_ vssd1 vssd1 vccd1 vccd1 _02882_
+ sky130_fd_sc_hd__a221o_1
X_14415_ net844 ag2.body\[528\] ag2.body\[529\] net837 vssd1 vssd1 vccd1 vccd1 _08576_
+ sky130_fd_sc_hd__a2bb2o_1
X_11627_ net504 _06598_ _06599_ net475 vssd1 vssd1 vccd1 vccd1 _06600_ sky130_fd_sc_hd__o31a_1
X_18183_ obsg2.obstacleArray\[88\] _03730_ net531 vssd1 vssd1 vccd1 vccd1 _01339_
+ sky130_fd_sc_hd__o21a_1
X_15395_ net2647 net82 _01596_ control.body\[644\] vssd1 vssd1 vccd1 vccd1 _00686_
+ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_7_Left_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10129__A net1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_117_3887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10034__A2 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11231__A1 net1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14346_ net970 _04220_ _04221_ net1006 _08500_ vssd1 vssd1 vccd1 vccd1 _08507_ sky130_fd_sc_hd__a221o_1
X_17134_ ag2.body\[519\] net932 vssd1 vssd1 vccd1 vccd1 _02813_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_117_3898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11558_ obsg2.obstacleArray\[66\] net633 _06465_ obsg2.obstacleArray\[70\] net507
+ vssd1 vssd1 vccd1 vccd1 _06531_ sky130_fd_sc_hd__o221a_1
XANTENNA__11231__B2 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1205 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold608 control.divider.count\[20\] vssd1 vssd1 vccd1 vccd1 net2170 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17065_ ag2.body\[25\] net868 vssd1 vssd1 vccd1 vccd1 _02744_ sky130_fd_sc_hd__nand2_1
X_10509_ _05474_ _05479_ _05480_ _05481_ vssd1 vssd1 vccd1 vccd1 _05482_ sky130_fd_sc_hd__and4_1
X_14277_ net986 ag2.body\[138\] vssd1 vssd1 vccd1 vccd1 _08438_ sky130_fd_sc_hd__xor2_1
XANTENNA__16170__A1 net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold619 control.body\[1088\] vssd1 vssd1 vccd1 vccd1 net2181 sky130_fd_sc_hd__dlygate4sd3_1
X_11489_ net1198 net1079 vssd1 vssd1 vccd1 vccd1 _06462_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10990__B1 net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16016_ _01689_ _01694_ vssd1 vssd1 vccd1 vccd1 _01695_ sky130_fd_sc_hd__nor2_2
XANTENNA__09727__A2 net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13228_ img_gen.tracker.frame\[382\] net658 vssd1 vssd1 vccd1 vccd1 _07804_ sky130_fd_sc_hd__and2_1
XFILLER_0_0_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_1563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16458__C1 net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12731__A1 net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09924__Y _04897_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13159_ net231 _07770_ _07771_ net1696 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[345\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_97_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09653__A net1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17967_ net319 _03531_ net296 vssd1 vssd1 vccd1 vccd1 _03591_ sky130_fd_sc_hd__or3b_1
XANTENNA__13287__A2 _07827_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15681__B1 _01627_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13175__A net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19706_ clknet_leaf_134_clk _00650_ net1307 vssd1 vssd1 vccd1 vccd1 control.body\[680\]
+ sky130_fd_sc_hd__dfrtp_1
X_16918_ ag2.body\[566\] net698 net689 ag2.body\[567\] _02596_ vssd1 vssd1 vccd1 vccd1
+ _02597_ sky130_fd_sc_hd__o221a_1
X_17898_ net354 _03531_ vssd1 vssd1 vccd1 vccd1 _03534_ sky130_fd_sc_hd__nor2_1
XANTENNA__16225__A2 net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19637_ clknet_leaf_124_clk _00581_ net1405 vssd1 vssd1 vccd1 vccd1 control.body\[755\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11407__B net1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16849_ net704 ag2.body\[173\] _04052_ net884 vssd1 vssd1 vccd1 vccd1 _02528_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_117_1622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_0_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15390__A _05857_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20567__CLK clknet_leaf_43_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19568_ clknet_leaf_116_clk _00512_ net1389 vssd1 vssd1 vccd1 vccd1 control.body\[830\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_76_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14718__B ag2.body\[341\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12798__A1 net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09321_ _04319_ net272 sound_gen.osc1.count\[0\] vssd1 vssd1 vccd1 vccd1 _01435_
+ sky130_fd_sc_hd__mux2_1
X_18519_ net1514 net1508 vssd1 vssd1 vccd1 vccd1 _00050_ sky130_fd_sc_hd__or2_1
XFILLER_0_125_96 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19499_ clknet_leaf_113_clk _00443_ net1396 vssd1 vssd1 vccd1 vccd1 control.body\[889\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_1430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11423__A net1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09252_ img_gen.updater.commands.rR1.rainbowRNG\[6\] vssd1 vssd1 vccd1 vccd1 _04277_
+ sky130_fd_sc_hd__inv_2
XANTENNA__15736__B2 ag2.body\[340\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16933__B net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11142__B net1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15200__A3 _04758_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09183_ ag2.body\[564\] vssd1 vssd1 vccd1 vccd1 _04208_ sky130_fd_sc_hd__inv_2
XANTENNA__10039__A net1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17426__A2_N net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11758__C1 net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout225_A net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20412_ clknet_leaf_32_clk _01299_ net1352 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[48\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_133_4390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09828__A net1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18150__A2 _03577_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11773__A2 net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20343_ clknet_leaf_140_clk _01234_ net1292 vssd1 vssd1 vccd1 vccd1 img_gen.updater.commands.rR1.rainbowRNG\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1134_A net1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20274_ clknet_leaf_42_clk net1586 net1373 vssd1 vssd1 vccd1 vccd1 control.button3.Q\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__17764__B _03299_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout594_A net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16160__S net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_1990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_4183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08967_ ag2.body\[50\] vssd1 vssd1 vccd1 vccd1 _03992_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_127_4194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout761_A net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout859_A net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_123_4069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10502__A net1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_4_clk_X clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18957__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10221__B net1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16621__C1 net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10500__A3 _05462_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10860_ net1072 control.body\[694\] vssd1 vssd1 vccd1 vccd1 _05833_ sky130_fd_sc_hd__xor2_1
XFILLER_0_6_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout40_A _03702_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12789__A1 net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09519_ net896 net900 net890 vssd1 vssd1 vccd1 vccd1 _04492_ sky130_fd_sc_hd__a21o_1
XANTENNA__17779__X _03458_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10791_ _05756_ _05757_ _05760_ _05762_ vssd1 vssd1 vccd1 vccd1 _05764_ sky130_fd_sc_hd__or4_1
XANTENNA_fanout814_X net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11997__C1 net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_979 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11333__A net1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12530_ img_gen.tracker.frame\[26\] net651 _07461_ vssd1 vssd1 vccd1 vccd1 _07462_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_52_1175 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10264__A2 _04471_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17939__B net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16843__B net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12461_ _06644_ _07307_ vssd1 vssd1 vccd1 vccd1 _07419_ sky130_fd_sc_hd__and2b_1
XANTENNA__18116__A net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14200_ net833 ag2.body\[361\] ag2.body\[362\] net826 vssd1 vssd1 vccd1 vccd1 _08361_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_10_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11412_ net1149 control.body\[851\] vssd1 vssd1 vccd1 vccd1 _06385_ sky130_fd_sc_hd__xor2_1
XFILLER_0_69_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15180_ control.body\[846\] net101 _01571_ net2355 vssd1 vssd1 vccd1 vccd1 _00496_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_34_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12392_ net1217 _07354_ _07356_ _07295_ _07353_ vssd1 vssd1 vccd1 vccd1 _07357_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_50_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16688__C1 _02228_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14131_ net807 ag2.body\[373\] _08288_ _08291_ vssd1 vssd1 vccd1 vccd1 _08292_ sky130_fd_sc_hd__a211o_1
XANTENNA__12961__A1 net254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11343_ ag2.body\[440\] net1224 vssd1 vssd1 vccd1 vccd1 _06316_ sky130_fd_sc_hd__xor2_1
XANTENNA__17955__A net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16152__A1 net379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_3740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_3751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14062_ _08221_ _08222_ vssd1 vssd1 vccd1 vccd1 _08223_ sky130_fd_sc_hd__nand2_1
X_11274_ ag2.body\[122\] net1186 vssd1 vssd1 vccd1 vccd1 _06247_ sky130_fd_sc_hd__xor2_1
XFILLER_0_39_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12713__A1 net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13013_ net288 _07699_ _07700_ net1902 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[269\]
+ sky130_fd_sc_hd__a22o_1
X_10225_ ag2.body\[564\] net1132 vssd1 vssd1 vccd1 vccd1 _05198_ sky130_fd_sc_hd__xor2_1
XANTENNA__16070__S net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18870_ clknet_leaf_26_clk img_gen.tracker.next_frame\[308\] net1344 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[308\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__10724__B1 net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17821_ _03974_ _08124_ vssd1 vssd1 vccd1 vccd1 _03487_ sky130_fd_sc_hd__xnor2_1
X_10156_ ag2.body\[62\] net1080 vssd1 vssd1 vccd1 vccd1 _05129_ sky130_fd_sc_hd__xor2_1
XANTENNA__18559__Q ag2.x\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14466__B2 net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20174__RESET_B net1480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold5 control.divider.detect.signal vssd1 vssd1 vccd1 vccd1 net1567 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12477__B1 net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17752_ _02722_ _02928_ _02938_ _02994_ vssd1 vssd1 vccd1 vccd1 _03431_ sky130_fd_sc_hd__and4_1
X_10087_ net1193 control.body\[793\] vssd1 vssd1 vccd1 vccd1 _05060_ sky130_fd_sc_hd__xor2_1
X_14964_ control.body\[1038\] net159 _01547_ net2339 vssd1 vssd1 vccd1 vccd1 _00304_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_106_3544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1632 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_106_3555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16703_ obsg2.obstacleArray\[86\] net488 net484 obsg2.obstacleArray\[85\] _02381_
+ vssd1 vssd1 vccd1 vccd1 _02382_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_106_3566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13915_ ag2.body\[60\] net120 _08151_ ag2.body\[52\] vssd1 vssd1 vccd1 vccd1 _00141_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_76_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14218__A1 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_3419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17683_ _04169_ net848 net710 ag2.body\[476\] vssd1 vssd1 vccd1 vccd1 _03362_ sky130_fd_sc_hd__a22o_1
XANTENNA__14218__B2 net813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14895_ net2181 net177 _01540_ control.body\[1080\] vssd1 vssd1 vccd1 vccd1 _00242_
+ sky130_fd_sc_hd__a22o_1
XANTENNA_clkload3_A clknet_4_7__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19882__CLK clknet_leaf_83_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11942__S net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_1529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13723__A net26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19422_ clknet_leaf_111_clk _00366_ net1427 vssd1 vssd1 vccd1 vccd1 control.body\[972\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16634_ obsg2.obstacleArray\[58\] net445 vssd1 vssd1 vccd1 vccd1 _02313_ sky130_fd_sc_hd__or2_1
XFILLER_0_18_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13846_ ag2.body\[10\] net116 _08133_ ag2.body\[2\] vssd1 vssd1 vccd1 vccd1 _00090_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_71_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19353_ clknet_leaf_101_clk _00297_ net1438 vssd1 vssd1 vccd1 vccd1 control.body\[1047\]
+ sky130_fd_sc_hd__dfrtp_1
X_16565_ _02207_ _02242_ vssd1 vssd1 vccd1 vccd1 _02244_ sky130_fd_sc_hd__nand2_1
X_13777_ img_gen.updater.commands.count\[10\] _07235_ _08081_ vssd1 vssd1 vccd1 vccd1
+ _08088_ sky130_fd_sc_hd__and3_1
XANTENNA__17168__B1 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10989_ _04605_ _05956_ _05960_ _05961_ vssd1 vssd1 vccd1 vccd1 _05962_ sky130_fd_sc_hd__nor4_1
XFILLER_0_70_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_80_2751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_2762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18304_ net323 _03787_ _03793_ net321 vssd1 vssd1 vccd1 vccd1 _03800_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_127_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_119_3938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_2773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19112__CLK clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15516_ ag2.body\[536\] net155 _01609_ ag2.body\[528\] vssd1 vssd1 vccd1 vccd1 _00794_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_119_3949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12728_ net683 _07568_ vssd1 vssd1 vccd1 vccd1 _07569_ sky130_fd_sc_hd__nor2_1
XFILLER_0_73_927 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19284_ clknet_leaf_98_clk _00228_ net1447 vssd1 vssd1 vccd1 vccd1 control.body\[1106\]
+ sky130_fd_sc_hd__dfrtp_1
X_16496_ obsg2.obstacleArray\[28\] obsg2.obstacleArray\[29\] obsg2.obstacleArray\[30\]
+ obsg2.obstacleArray\[31\] net458 net400 vssd1 vssd1 vccd1 vccd1 _02175_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_61_2172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_2183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18235_ obsg2.obstacleArray\[114\] _03756_ net527 vssd1 vssd1 vccd1 vccd1 _01365_
+ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_61_2194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12659_ net262 _07533_ _07534_ net1944 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[82\]
+ sky130_fd_sc_hd__a22o_1
X_15447_ ag2.body\[603\] net86 _01601_ ag2.body\[595\] vssd1 vssd1 vccd1 vccd1 _00733_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__14554__A net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12626__X _07515_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18026__A net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11530__X _06503_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09648__A net1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18166_ net351 _03539_ _03705_ obsg2.obstacleArray\[80\] vssd1 vssd1 vccd1 vccd1
+ _03722_ sky130_fd_sc_hd__a31o_1
XFILLER_0_128_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15378_ control.body\[669\] net68 _01594_ net2403 vssd1 vssd1 vccd1 vccd1 _00671_
+ sky130_fd_sc_hd__a22o_1
X_20599__1531 vssd1 vssd1 vccd1 vccd1 _20599__1531/HI net1531 sky130_fd_sc_hd__conb_1
XANTENNA__20325__SET_B net1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12345__Y _07312_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16679__C1 net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11755__A2 net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17117_ ag2.body\[536\] net739 net727 ag2.body\[538\] vssd1 vssd1 vccd1 vccd1 _02796_
+ sky130_fd_sc_hd__a22o_1
X_14329_ net835 ag2.body\[425\] _04152_ net1029 vssd1 vssd1 vccd1 vccd1 _08490_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_78_2691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10146__X _05119_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold405 img_gen.tracker.frame\[86\] vssd1 vssd1 vccd1 vccd1 net1967 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_561 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18097_ obsg2.obstacleArray\[52\] _03680_ net524 vssd1 vssd1 vccd1 vccd1 _01303_
+ sky130_fd_sc_hd__o21a_1
XANTENNA__14841__X _01512_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold416 img_gen.tracker.frame\[324\] vssd1 vssd1 vccd1 vccd1 net1978 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10963__B1 _05919_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold427 img_gen.tracker.frame\[428\] vssd1 vssd1 vccd1 vccd1 net1989 sky130_fd_sc_hd__dlygate4sd3_1
Xhold438 img_gen.tracker.frame\[65\] vssd1 vssd1 vccd1 vccd1 net2000 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12505__C net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17048_ ag2.body\[257\] net735 net711 ag2.body\[260\] vssd1 vssd1 vccd1 vccd1 _02727_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_74_2566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold449 img_gen.tracker.frame\[482\] vssd1 vssd1 vccd1 vccd1 net2011 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_2588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09870_ ag2.body\[156\] net1139 vssd1 vssd1 vccd1 vccd1 _04843_ sky130_fd_sc_hd__xor2_1
Xfanout907 net908 vssd1 vssd1 vccd1 vccd1 net907 sky130_fd_sc_hd__buf_4
Xfanout918 net919 vssd1 vssd1 vccd1 vccd1 net918 sky130_fd_sc_hd__clkbuf_2
XANTENNA__12802__A net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout929 obsg2.randCord\[7\] vssd1 vssd1 vccd1 vccd1 net929 sky130_fd_sc_hd__buf_4
XANTENNA__16446__A2 _02059_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14457__A1 net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18999_ clknet_leaf_2_clk img_gen.tracker.next_frame\[437\] net1248 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[437\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__14457__B2 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11418__A net1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11137__B _04420_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09884__A1 ag2.body\[161\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09884__B2 ag2.body\[164\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15406__B1 _01581_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16603__C1 net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10494__A2 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13352__B net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_743 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1084_A net1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09304_ sound_gen.osc1.count\[4\] _04323_ vssd1 vssd1 vccd1 vccd1 _04324_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_135_4430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_4441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16906__B1 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_135_4452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09235_ obsg2.arraySet vssd1 vssd1 vccd1 vccd1 _04260_ sky130_fd_sc_hd__inv_2
XANTENNA__11994__A2 net600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_4305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_131_4316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16155__S net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_4327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14464__A net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout607_A net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_1533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09939__A2 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09558__A net1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09166_ ag2.body\[516\] vssd1 vssd1 vccd1 vccd1 _04191_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_40_1555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15994__S net223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19098__RESET_B net1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09097_ ag2.body\[347\] vssd1 vssd1 vccd1 vccd1 _04122_ sky130_fd_sc_hd__inv_2
XFILLER_0_62_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1137_X net1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09845__X _04818_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20326_ clknet_leaf_46_clk _01222_ net1377 vssd1 vssd1 vccd1 vccd1 ag2.body\[7\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_43_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold950 control.body\[734\] vssd1 vssd1 vccd1 vccd1 net2512 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_4245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_3080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout976_A ag2.randCord\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold961 control.body\[895\] vssd1 vssd1 vccd1 vccd1 net2523 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout597_X net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1580 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_129_4256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_79_Left_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold972 _00432_ vssd1 vssd1 vccd1 vccd1 net2534 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20257_ clknet_leaf_70_clk _01201_ net1497 vssd1 vssd1 vccd1 vccd1 ag2.body\[143\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_129_4267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold983 control.body\[849\] vssd1 vssd1 vccd1 vccd1 net2545 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold994 control.body\[976\] vssd1 vssd1 vccd1 vccd1 net2556 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10010_ _04433_ net638 vssd1 vssd1 vccd1 vccd1 _04983_ sky130_fd_sc_hd__nor2_1
XANTENNA__09572__B1 net1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_1495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13527__B net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout764_X net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09999_ net1145 control.body\[731\] vssd1 vssd1 vccd1 vccd1 _04972_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_34_1359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14448__A1 net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09724__C net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20188_ clknet_leaf_89_clk _01132_ net1454 vssd1 vssd1 vccd1 vccd1 ag2.body\[202\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__15645__B1 _01623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14448__B2 net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17941__C _03570_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13246__C _07439_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16397__Y _02076_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11047__B net1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11961_ img_gen.tracker.frame\[499\] net544 vssd1 vssd1 vccd1 vccd1 _06933_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout931_X net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17398__B1 net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13700_ _04635_ _08039_ _08040_ vssd1 vssd1 vccd1 vccd1 _08041_ sky130_fd_sc_hd__o21a_1
X_10912_ _04538_ _04980_ _04447_ vssd1 vssd1 vccd1 vccd1 _05885_ sky130_fd_sc_hd__a21bo_1
X_14680_ net973 _04140_ _04141_ net1018 _08840_ vssd1 vssd1 vccd1 vccd1 _08841_ sky130_fd_sc_hd__a221o_1
XANTENNA__09740__B net1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19135__CLK clknet_leaf_132_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10485__A2 net1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11892_ img_gen.tracker.frame\[85\] img_gen.tracker.frame\[88\] img_gen.tracker.frame\[91\]
+ img_gen.tracker.frame\[94\] net1219 net1195 vssd1 vssd1 vccd1 vccd1 _06864_ sky130_fd_sc_hd__mux4_1
XANTENNA_fanout43_X net43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13631_ control.divider.count\[11\] control.divider.count\[10\] _07992_ vssd1 vssd1
+ vccd1 vccd1 _07995_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_88_Left_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10843_ ag2.body\[42\] net774 net766 ag2.body\[44\] vssd1 vssd1 vccd1 vccd1 _05816_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_131_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14620__A1 net1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14620__B2 net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16350_ _01919_ _02004_ _02012_ _02028_ _01929_ vssd1 vssd1 vccd1 vccd1 _02029_ sky130_fd_sc_hd__o311a_1
X_13562_ ssdec1.in\[1\] _04282_ _07941_ _07937_ vssd1 vssd1 vccd1 vccd1 net19 sky130_fd_sc_hd__a31oi_1
XFILLER_0_55_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17669__B net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10774_ ag2.body\[222\] net1091 vssd1 vssd1 vccd1 vccd1 _05747_ sky130_fd_sc_hd__xor2_1
XFILLER_0_67_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14578__A1_N net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15301_ control.body\[728\] net77 _01586_ control.body\[720\] vssd1 vssd1 vccd1 vccd1
+ _00602_ sky130_fd_sc_hd__a22o_1
XANTENNA__19285__CLK clknet_leaf_98_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12513_ _06638_ net439 net565 net551 vssd1 vssd1 vccd1 vccd1 _07453_ sky130_fd_sc_hd__or4_2
X_16281_ obsg2.obstacleArray\[22\] obsg2.obstacleArray\[23\] net412 vssd1 vssd1 vccd1
+ vccd1 _01960_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_97_3267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13493_ net250 _07908_ _07909_ net2067 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[541\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__14374__A net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_97_3278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_114_3802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18020_ obsg2.obstacleArray\[26\] _03629_ net531 vssd1 vssd1 vccd1 vccd1 _01277_
+ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_114_3813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_97_3289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13187__A1 net241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15232_ control.body\[796\] net98 _01577_ net2395 vssd1 vssd1 vccd1 vccd1 _00542_
+ sky130_fd_sc_hd__a22o_1
X_12444_ net1192 _07379_ _07404_ net589 vssd1 vssd1 vccd1 vccd1 _07405_ sky130_fd_sc_hd__a22o_1
XANTENNA__17956__Y _03582_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1300 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20262__CLK clknet_leaf_43_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12934__A1 net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11737__A2 net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15163_ control.body\[863\] net98 _01569_ net2405 vssd1 vssd1 vccd1 vccd1 _00481_
+ sky130_fd_sc_hd__a22o_1
X_12375_ img_gen.updater.commands.count\[10\] img_gen.updater.commands.count\[11\]
+ img_gen.updater.commands.count\[8\] img_gen.updater.commands.count\[9\] vssd1 vssd1
+ vccd1 vccd1 _07340_ sky130_fd_sc_hd__or4_1
XANTENNA__10407__A net1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_97_Left_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14114_ net971 ag2.body\[571\] vssd1 vssd1 vccd1 vccd1 _08275_ sky130_fd_sc_hd__xor2_1
XANTENNA__16676__A2 net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11326_ _06295_ _06296_ _06297_ _06298_ vssd1 vssd1 vccd1 vccd1 _06299_ sky130_fd_sc_hd__or4_1
X_19971_ clknet_leaf_62_clk _00915_ net1470 vssd1 vssd1 vccd1 vccd1 ag2.body\[417\]
+ sky130_fd_sc_hd__dfrtp_4
X_15094_ control.body\[912\] net148 _01563_ net2150 vssd1 vssd1 vccd1 vccd1 _00418_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__14687__A1 net986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14687__B2 net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1518 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14045_ net1025 ag2.body\[189\] vssd1 vssd1 vccd1 vccd1 _08206_ sky130_fd_sc_hd__xor2_1
X_18922_ clknet_leaf_140_clk img_gen.tracker.next_frame\[360\] net1291 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[360\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__09474__Y _04447_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11257_ net1075 control.body\[774\] vssd1 vssd1 vccd1 vccd1 _06230_ sky130_fd_sc_hd__xnor2_1
XANTENNA__12622__A net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12698__B1 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_108_3606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10208_ net1229 control.body\[992\] vssd1 vssd1 vccd1 vccd1 _05181_ sky130_fd_sc_hd__nand2_1
XANTENNA__12162__A2 net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_3617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1131 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10845__A1_N net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18853_ clknet_leaf_18_clk img_gen.tracker.next_frame\[291\] net1323 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[291\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_108_3628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11188_ ag2.body\[178\] net774 _06153_ _06155_ _06156_ vssd1 vssd1 vccd1 vccd1 _06161_
+ sky130_fd_sc_hd__a2111o_1
XANTENNA__14439__A1 net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14439__B2 net1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17804_ _03288_ _03469_ _03473_ vssd1 vssd1 vccd1 vccd1 _01218_ sky130_fd_sc_hd__and3b_1
X_10139_ net1201 control.body\[817\] vssd1 vssd1 vccd1 vccd1 _05112_ sky130_fd_sc_hd__xor2_1
XANTENNA__10142__A net1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18784_ clknet_leaf_12_clk img_gen.tracker.next_frame\[222\] net1284 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[222\] sky130_fd_sc_hd__dfrtp_1
X_15996_ control.fsm.temp\[2\] control.body_update.direction\[2\] net223 vssd1 vssd1
+ vccd1 vccd1 _01208_ sky130_fd_sc_hd__mux2_1
XANTENNA__14844__D1 _01499_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17735_ _03248_ _03251_ _03412_ _03413_ _02652_ vssd1 vssd1 vccd1 vccd1 _03414_ sky130_fd_sc_hd__o2111a_1
X_14947_ net2571 net168 _01545_ net2141 vssd1 vssd1 vccd1 vccd1 _00289_ sky130_fd_sc_hd__a22o_1
XANTENNA__17389__B1 net728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13662__A2 net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15939__A1 ag2.body\[161\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17666_ ag2.body\[451\] net851 vssd1 vssd1 vccd1 vccd1 _03345_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_82_2824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_2370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14878_ control.body\[1105\] net179 _01538_ control.body\[1097\] vssd1 vssd1 vccd1
+ vccd1 _00227_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_67_2381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10796__B net1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19405_ clknet_leaf_103_clk _00349_ net1432 vssd1 vssd1 vccd1 vccd1 control.body\[987\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_63_2234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16617_ net394 _02295_ _02294_ net361 vssd1 vssd1 vccd1 vccd1 _02296_ sky130_fd_sc_hd__a211o_1
XFILLER_0_15_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13829_ _08124_ _08125_ _08123_ vssd1 vssd1 vccd1 vccd1 _08126_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_9_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_63_2245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14611__A1 net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17597_ _03009_ _03021_ _03022_ _03275_ vssd1 vssd1 vccd1 vccd1 _03276_ sky130_fd_sc_hd__or4b_1
XTAP_TAPCELL_ROW_63_2256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14611__B2 net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1624 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19336_ clknet_leaf_100_clk net2299 net1443 vssd1 vssd1 vccd1 vccd1 control.body\[1062\]
+ sky130_fd_sc_hd__dfrtp_1
X_16548_ net461 _02220_ vssd1 vssd1 vccd1 vccd1 _02227_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_46_927 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17579__B net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16483__B net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11976__A2 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19267_ clknet_leaf_71_clk _00211_ net1503 vssd1 vssd1 vccd1 vccd1 ag2.body\[130\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_116_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_14_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16479_ obsg2.obstacleArray\[38\] net452 vssd1 vssd1 vccd1 vccd1 _02158_ sky130_fd_sc_hd__or2_1
XFILLER_0_5_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09020_ ag2.body\[154\] vssd1 vssd1 vccd1 vccd1 _04045_ sky130_fd_sc_hd__inv_2
X_18218_ _03660_ net40 vssd1 vssd1 vccd1 vccd1 _03748_ sky130_fd_sc_hd__nor2_1
XFILLER_0_72_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18652__CLK clknet_leaf_131_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19198_ clknet_leaf_53_clk _00142_ net1455 vssd1 vssd1 vccd1 vccd1 ag2.body\[61\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__11189__B1 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_2628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_2639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18149_ net529 _03713_ vssd1 vssd1 vccd1 vccd1 _01322_ sky130_fd_sc_hd__and2_1
XANTENNA__19191__RESET_B net1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold202 img_gen.tracker.frame\[58\] vssd1 vssd1 vccd1 vccd1 net1764 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10936__B1 _05798_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_2049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold213 img_gen.tracker.frame\[128\] vssd1 vssd1 vccd1 vccd1 net1775 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_339 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold224 img_gen.tracker.frame\[25\] vssd1 vssd1 vccd1 vccd1 net1786 sky130_fd_sc_hd__dlygate4sd3_1
Xhold235 img_gen.tracker.frame\[312\] vssd1 vssd1 vccd1 vccd1 net1797 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold246 img_gen.tracker.frame\[216\] vssd1 vssd1 vccd1 vccd1 net1808 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14678__A1 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19008__CLK clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14678__B2 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold257 img_gen.tracker.frame\[229\] vssd1 vssd1 vccd1 vccd1 net1819 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1607 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20111_ clknet_leaf_79_clk _01055_ net1487 vssd1 vssd1 vccd1 vccd1 ag2.body\[285\]
+ sky130_fd_sc_hd__dfrtp_4
Xhold268 img_gen.tracker.frame\[463\] vssd1 vssd1 vccd1 vccd1 net1830 sky130_fd_sc_hd__dlygate4sd3_1
X_09922_ ag2.body\[312\] net788 net772 ag2.body\[315\] _04894_ vssd1 vssd1 vccd1 vccd1
+ _04895_ sky130_fd_sc_hd__a221o_1
Xhold279 img_gen.tracker.frame\[203\] vssd1 vssd1 vccd1 vccd1 net1841 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1175 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12532__A net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout704 net705 vssd1 vssd1 vccd1 vccd1 net704 sky130_fd_sc_hd__buf_2
XFILLER_0_102_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout715 net716 vssd1 vssd1 vccd1 vccd1 net715 sky130_fd_sc_hd__clkbuf_4
XANTENNA__13350__A1 net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout726 net727 vssd1 vssd1 vccd1 vccd1 net726 sky130_fd_sc_hd__clkbuf_4
Xfanout737 _04262_ vssd1 vssd1 vccd1 vccd1 net737 sky130_fd_sc_hd__buf_4
X_20042_ clknet_leaf_68_clk _00986_ net1498 vssd1 vssd1 vccd1 vccd1 ag2.body\[344\]
+ sky130_fd_sc_hd__dfrtp_4
X_09853_ net1181 control.body\[970\] vssd1 vssd1 vccd1 vccd1 _04826_ sky130_fd_sc_hd__xor2_1
XANTENNA__13347__B _07515_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_4120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout748 _04233_ vssd1 vssd1 vccd1 vccd1 net748 sky130_fd_sc_hd__buf_4
XANTENNA__15627__B1 _01621_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout759 net760 vssd1 vssd1 vccd1 vccd1 net759 sky130_fd_sc_hd__buf_4
XANTENNA_fanout292_A net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17711__S1 net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11900__A2 net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09784_ net1110 control.body\[949\] vssd1 vssd1 vccd1 vccd1 _04757_ sky130_fd_sc_hd__xor2_1
XANTENNA__09841__A net1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13363__A net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout557_A _06651_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1299_A net1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_137_4503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_137_4514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13082__B _07564_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_1720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14602__A1 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout724_A net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14602__B2 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1087_X net1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10219__A2 _04758_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_27_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_27_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_42_1617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16355__A1 net420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_142_clk clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_142_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_23_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09218_ control.body\[815\] vssd1 vssd1 vccd1 vccd1 _04243_ sky130_fd_sc_hd__inv_2
XFILLER_0_17_673 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10490_ ag2.body\[546\] net1180 vssd1 vssd1 vccd1 vccd1 _05463_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_51_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_92_3120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_3131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11719__A2 _06644_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12916__A1 net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_3142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09149_ ag2.body\[482\] vssd1 vssd1 vccd1 vccd1 _04174_ sky130_fd_sc_hd__inv_2
XANTENNA__17709__S net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13184__A4 _07515_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17936__C _03566_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12160_ img_gen.tracker.frame\[384\] net618 net542 img_gen.tracker.frame\[390\] vssd1
+ vssd1 vccd1 vccd1 _07132_ sky130_fd_sc_hd__o22a_1
XFILLER_0_60_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout881_X net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11111_ net775 control.body\[1098\] _06081_ _06082_ _06083_ vssd1 vssd1 vccd1 vccd1
+ _06084_ sky130_fd_sc_hd__o2111a_1
XANTENNA_fanout979_X net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20309_ clknet_leaf_21_clk _01209_ net1361 vssd1 vssd1 vccd1 vccd1 obsg2.arraySet
+ sky130_fd_sc_hd__dfrtp_1
X_12091_ net577 _07062_ vssd1 vssd1 vccd1 vccd1 _07063_ sky130_fd_sc_hd__or2_1
Xhold780 control.body\[738\] vssd1 vssd1 vccd1 vccd1 net2342 sky130_fd_sc_hd__dlygate4sd3_1
Xhold791 control.body\[933\] vssd1 vssd1 vccd1 vccd1 net2353 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_6_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12144__A2 net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11042_ _06005_ _06007_ _06011_ _06014_ vssd1 vssd1 vccd1 vccd1 _06015_ sky130_fd_sc_hd__and4b_1
XANTENNA__17952__B net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18280__A1 net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15850_ ag2.body\[242\] net173 _01645_ ag2.body\[234\] vssd1 vssd1 vccd1 vccd1 _01092_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_36_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14801_ _01470_ _01471_ _01468_ _01469_ vssd1 vssd1 vccd1 vccd1 _01472_ sky130_fd_sc_hd__a211o_1
XANTENNA__16830__A2 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15781_ ag2.body\[308\] net209 _01638_ ag2.body\[300\] vssd1 vssd1 vccd1 vccd1 _01030_
+ sky130_fd_sc_hd__a22o_1
X_12993_ net233 _07691_ _07692_ net1956 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[258\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_118_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_1613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20598__1530 vssd1 vssd1 vccd1 vccd1 _20598__1530/HI net1530 sky130_fd_sc_hd__conb_1
X_17520_ ag2.body\[480\] net881 vssd1 vssd1 vccd1 vccd1 _03199_ sky130_fd_sc_hd__xor2_1
XFILLER_0_8_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13273__A net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14732_ net993 ag2.body\[113\] vssd1 vssd1 vccd1 vccd1 _08893_ sky130_fd_sc_hd__or2_1
XFILLER_0_98_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11944_ img_gen.tracker.frame\[142\] net585 net544 img_gen.tracker.frame\[139\] _06915_
+ vssd1 vssd1 vccd1 vccd1 _06916_ sky130_fd_sc_hd__o221a_1
XFILLER_0_118_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17451_ ag2.body\[434\] net724 net717 ag2.body\[435\] vssd1 vssd1 vccd1 vccd1 _03130_
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_73_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11875_ img_gen.tracker.frame\[256\] net598 net582 img_gen.tracker.frame\[262\] vssd1
+ vssd1 vccd1 vccd1 _06847_ sky130_fd_sc_hd__o22a_1
X_14663_ net1001 ag2.body\[520\] vssd1 vssd1 vccd1 vccd1 _08824_ sky130_fd_sc_hd__xor2_1
XFILLER_0_15_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_99_3329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16402_ obsg2.obstacleArray\[108\] obsg2.obstacleArray\[109\] net453 vssd1 vssd1
+ vccd1 vccd1 _02081_ sky130_fd_sc_hd__mux2_1
X_13614_ _07959_ _07984_ vssd1 vssd1 vccd1 vccd1 control.divider.next_count\[4\] sky130_fd_sc_hd__nor2_1
X_10826_ ag2.body\[308\] net1141 vssd1 vssd1 vccd1 vccd1 _05799_ sky130_fd_sc_hd__xor2_1
XFILLER_0_39_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17382_ ag2.body\[488\] net886 vssd1 vssd1 vccd1 vccd1 _03061_ sky130_fd_sc_hd__xor2_1
XFILLER_0_89_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14594_ net845 ag2.body\[304\] ag2.body\[308\] net815 vssd1 vssd1 vccd1 vccd1 _08755_
+ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__19920__CLK clknet_leaf_53_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19121_ clknet_leaf_141_clk img_gen.tracker.next_frame\[559\] net1294 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[559\] sky130_fd_sc_hd__dfrtp_1
X_16333_ net371 _02011_ _02008_ _01912_ vssd1 vssd1 vccd1 vccd1 _02012_ sky130_fd_sc_hd__o211a_1
XFILLER_0_6_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10757_ net1179 control.body\[890\] vssd1 vssd1 vccd1 vccd1 _05730_ sky130_fd_sc_hd__nand2_1
X_13545_ net2156 net659 _07929_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[573\]
+ sky130_fd_sc_hd__and3_1
XANTENNA__12080__A1 net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_995 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_472 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_133_clk clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_133_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__11521__A _06490_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19052_ clknet_leaf_8_clk img_gen.tracker.next_frame\[490\] net1273 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[490\] sky130_fd_sc_hd__dfrtp_1
X_16264_ obsg2.obstacleArray\[48\] net405 vssd1 vssd1 vccd1 vccd1 _01943_ sky130_fd_sc_hd__or2_1
XANTENNA__16897__A2 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13476_ net666 _07902_ vssd1 vssd1 vccd1 vccd1 _07903_ sky130_fd_sc_hd__nor2_1
X_10688_ ag2.body\[151\] net1065 vssd1 vssd1 vccd1 vccd1 _05661_ sky130_fd_sc_hd__xor2_1
XFILLER_0_109_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_1439 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18003_ net299 _03616_ vssd1 vssd1 vccd1 vccd1 _03617_ sky130_fd_sc_hd__nand2_1
XANTENNA__12907__A1 net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15215_ net2176 net92 _01575_ net2517 vssd1 vssd1 vccd1 vccd1 _00527_ sky130_fd_sc_hd__a22o_1
X_12427_ _07354_ _07387_ _07388_ vssd1 vssd1 vccd1 vccd1 _07389_ sky130_fd_sc_hd__and3_1
XANTENNA__11240__B net1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16195_ net373 _01871_ _01873_ net346 vssd1 vssd1 vccd1 vccd1 _01874_ sky130_fd_sc_hd__a211o_1
XANTENNA__10137__A net1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_1197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12358_ _06631_ _06635_ vssd1 vssd1 vccd1 vccd1 _07325_ sky130_fd_sc_hd__nand2_1
XFILLER_0_26_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15146_ _04421_ _05051_ net50 vssd1 vssd1 vccd1 vccd1 _01568_ sky130_fd_sc_hd__o21a_2
XTAP_TAPCELL_ROW_71_2503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_1639 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11309_ _06278_ _06279_ _06280_ _06281_ vssd1 vssd1 vccd1 vccd1 _06282_ sky130_fd_sc_hd__or4_1
X_19954_ clknet_leaf_44_clk _00898_ net1381 vssd1 vssd1 vccd1 vccd1 ag2.body\[432\]
+ sky130_fd_sc_hd__dfrtp_4
X_15077_ control.body\[929\] net147 _01561_ net2250 vssd1 vssd1 vccd1 vccd1 _00403_
+ sky130_fd_sc_hd__a22o_1
X_12289_ _04389_ _07257_ _04391_ vssd1 vssd1 vccd1 vccd1 _07259_ sky130_fd_sc_hd__o21a_1
XFILLER_0_77_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12135__A2 net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14028_ _08184_ _08186_ _08187_ _08188_ vssd1 vssd1 vccd1 vccd1 _08189_ sky130_fd_sc_hd__or4_1
X_18905_ clknet_leaf_144_clk img_gen.tracker.next_frame\[343\] net1251 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[343\] sky130_fd_sc_hd__dfrtp_1
X_19885_ clknet_leaf_86_clk _00829_ net1462 vssd1 vssd1 vccd1 vccd1 ag2.body\[507\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__10146__A1 _04520_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12071__B net1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15609__B1 _01620_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18836_ clknet_leaf_141_clk img_gen.tracker.next_frame\[274\] net1262 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[274\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_69_2421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_2432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09661__A net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18767_ clknet_leaf_16_clk img_gen.tracker.next_frame\[205\] net1315 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[205\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__14279__A net994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15979_ net1043 _08119_ vssd1 vssd1 vccd1 vccd1 _01664_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_65_2307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_65_2318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17718_ obsg2.obstacleArray\[128\] obsg2.obstacleArray\[129\] net427 vssd1 vssd1
+ vccd1 vccd1 _03397_ sky130_fd_sc_hd__mux2_1
X_18698_ clknet_leaf_29_clk img_gen.tracker.next_frame\[136\] net1274 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[136\] sky130_fd_sc_hd__dfrtp_1
X_17649_ ag2.body\[32\] net880 vssd1 vssd1 vccd1 vccd1 _03328_ sky130_fd_sc_hd__xor2_1
XFILLER_0_8_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13399__A1 net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_318 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_450 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_532 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19319_ clknet_leaf_104_clk _00263_ net1433 vssd1 vssd1 vccd1 vccd1 control.body\[1077\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_46_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11949__A2 net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16337__A1 net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17102__B net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20591_ net1523 vssd1 vssd1 vccd1 vccd1 gpio_oeb[3] sky130_fd_sc_hd__buf_2
Xclkbuf_leaf_124_clk clknet_4_9__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_124_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__12527__A net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout138_A net139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_1675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16888__A2 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09003_ ag2.body\[120\] vssd1 vssd1 vccd1 vccd1 _04028_ sky130_fd_sc_hd__inv_2
XFILLER_0_84_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11150__B net1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13820__A_N _08113_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_102_clk_X clknet_leaf_102_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout305_A _07445_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1047_A net1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09836__A net1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11577__S net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13358__A net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout501 _01708_ vssd1 vssd1 vccd1 vccd1 net501 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_6_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1214_A ag2.y\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12126__A2 net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout512 net515 vssd1 vssd1 vccd1 vccd1 net512 sky130_fd_sc_hd__clkbuf_2
X_09905_ ag2.body\[130\] net1188 vssd1 vssd1 vccd1 vccd1 _04878_ sky130_fd_sc_hd__or2_1
XFILLER_0_10_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_1459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout523 net528 vssd1 vssd1 vccd1 vccd1 net523 sky130_fd_sc_hd__clkbuf_2
Xfanout534 _04395_ vssd1 vssd1 vccd1 vccd1 net534 sky130_fd_sc_hd__buf_2
XANTENNA__10053__Y _05026_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18548__CLK clknet_leaf_132_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout674_A _04393_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout545 net547 vssd1 vssd1 vccd1 vccd1 net545 sky130_fd_sc_hd__clkbuf_4
Xfanout556 _06651_ vssd1 vssd1 vccd1 vccd1 net556 sky130_fd_sc_hd__clkbuf_4
X_20025_ clknet_leaf_58_clk _00969_ net1471 vssd1 vssd1 vccd1 vccd1 ag2.body\[375\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__16499__S1 net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09836_ net1157 control.body\[923\] vssd1 vssd1 vccd1 vccd1 _04809_ sky130_fd_sc_hd__or2_1
Xfanout567 _06650_ vssd1 vssd1 vccd1 vccd1 net567 sky130_fd_sc_hd__buf_2
XANTENNA_fanout1002_X net1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout578 net579 vssd1 vssd1 vccd1 vccd1 net578 sky130_fd_sc_hd__buf_2
Xfanout589 net592 vssd1 vssd1 vccd1 vccd1 net589 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_119_1322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout462_X net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout841_A net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09767_ _04537_ _04599_ _04688_ vssd1 vssd1 vccd1 vccd1 _04740_ sky130_fd_sc_hd__o21a_2
XANTENNA__14823__A1 net994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14189__A net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14823__B2 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout939_A net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09698_ ag2.body\[69\] net1114 vssd1 vssd1 vccd1 vccd1 _04671_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_29_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11325__B net1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16608__S net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout727_X net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_1218 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16040__A3 net498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11660_ net753 net743 _06625_ _06632_ _06624_ vssd1 vssd1 vccd1 vccd1 _06633_ sky130_fd_sc_hd__a311o_1
XANTENNA__11044__C _05985_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10611_ net1087 control.body\[990\] vssd1 vssd1 vccd1 vccd1 _05584_ sky130_fd_sc_hd__xor2_1
X_11591_ obsg2.obstacleArray\[2\] obsg2.obstacleArray\[3\] obsg2.obstacleArray\[6\]
+ obsg2.obstacleArray\[7\] net1124 net513 vssd1 vssd1 vccd1 vccd1 _06564_ sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_115_clk clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_115_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_119_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_94_3204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13330_ net249 _07844_ _07845_ net1811 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[442\]
+ sky130_fd_sc_hd__a22o_1
X_10542_ ag2.body\[230\] net1085 vssd1 vssd1 vccd1 vccd1 _05515_ sky130_fd_sc_hd__nand2_1
XFILLER_0_91_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13261_ net257 _07817_ _07818_ net1756 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[400\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_134_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10473_ net1179 control.body\[1010\] vssd1 vssd1 vccd1 vccd1 _05446_ sky130_fd_sc_hd__xor2_1
XANTENNA__16343__S net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12212_ img_gen.control.current\[0\] _07183_ _07179_ net677 vssd1 vssd1 vccd1 vccd1
+ _07184_ sky130_fd_sc_hd__a2bb2o_1
X_15000_ control.body\[1006\] net153 _01551_ control.body\[998\] vssd1 vssd1 vccd1
+ vccd1 _00336_ sky130_fd_sc_hd__a22o_1
XANTENNA__09746__A net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13192_ net241 _07785_ _07786_ net1869 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[363\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11995__B net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15839__B1 _01644_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12143_ img_gen.tracker.frame\[504\] net617 vssd1 vssd1 vccd1 vccd1 _07115_ sky130_fd_sc_hd__or2_1
XANTENNA__16500__A1 net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_88_3008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12117__A2 net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_3019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16951_ ag2.body\[388\] net963 vssd1 vssd1 vccd1 vccd1 _02630_ sky130_fd_sc_hd__xor2_1
XANTENNA__17682__B net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12074_ img_gen.tracker.frame\[120\] net629 net556 img_gen.tracker.frame\[126\] vssd1
+ vssd1 vccd1 vccd1 _07046_ sky130_fd_sc_hd__a22o_1
XFILLER_0_47_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17056__A2 net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15902_ ag2.body\[192\] net129 _01651_ ag2.body\[184\] vssd1 vssd1 vccd1 vccd1 _01138_
+ sky130_fd_sc_hd__a22o_1
X_11025_ _05994_ _05995_ _05996_ _05997_ vssd1 vssd1 vccd1 vccd1 _05998_ sky130_fd_sc_hd__a22o_1
XFILLER_0_60_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19670_ clknet_leaf_134_clk _00614_ net1307 vssd1 vssd1 vccd1 vccd1 control.body\[724\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_95_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16882_ ag2.body\[20\] net958 vssd1 vssd1 vccd1 vccd1 _02561_ sky130_fd_sc_hd__xor2_1
XFILLER_0_95_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18621_ clknet_leaf_145_clk img_gen.tracker.next_frame\[59\] net1242 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[59\] sky130_fd_sc_hd__dfrtp_1
X_15833_ ag2.body\[259\] net175 net49 ag2.body\[251\] vssd1 vssd1 vccd1 vccd1 _01077_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__14099__A net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1129 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18552_ clknet_leaf_37_clk _00078_ net1351 vssd1 vssd1 vccd1 vccd1 control.divider.fsm.current_mode\[2\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__11628__A1 net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15764_ ag2.body\[325\] net214 _01636_ ag2.body\[317\] vssd1 vssd1 vccd1 vccd1 _01015_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__19883__RESET_B net1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10420__A net1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12976_ net2075 net646 _07684_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[249\]
+ sky130_fd_sc_hd__and3_1
XFILLER_0_34_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17503_ ag2.body\[233\] net735 net726 ag2.body\[234\] vssd1 vssd1 vccd1 vccd1 _03182_
+ sky130_fd_sc_hd__o22ai_1
X_14715_ net978 ag2.body\[339\] vssd1 vssd1 vccd1 vccd1 _08876_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_16_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18483_ net1515 net1509 vssd1 vssd1 vccd1 vccd1 _00014_ sky130_fd_sc_hd__or2_1
X_11927_ net566 _06898_ vssd1 vssd1 vccd1 vccd1 _06899_ sky130_fd_sc_hd__nand2_1
X_15695_ ag2.body\[376\] net137 _01628_ ag2.body\[368\] vssd1 vssd1 vccd1 vccd1 _00954_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_16_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17434_ ag2.body\[145\] net877 vssd1 vssd1 vccd1 vccd1 _03113_ sky130_fd_sc_hd__xor2_1
XFILLER_0_74_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14646_ net976 _04190_ ag2.body\[516\] net814 _08803_ vssd1 vssd1 vccd1 vccd1 _08807_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_86_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11858_ img_gen.tracker.frame\[229\] net623 net577 _06829_ vssd1 vssd1 vccd1 vccd1
+ _06830_ sky130_fd_sc_hd__o211a_1
XFILLER_0_131_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17365_ _03039_ _03041_ _03043_ _03005_ vssd1 vssd1 vccd1 vccd1 _03044_ sky130_fd_sc_hd__or4b_1
Xclkbuf_leaf_106_clk clknet_4_10__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_106_clk
+ sky130_fd_sc_hd__clkbuf_8
X_10809_ net1206 control.body\[1089\] vssd1 vssd1 vccd1 vccd1 _05782_ sky130_fd_sc_hd__xor2_1
XANTENNA_19 _08509_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14577_ _08735_ _08736_ _08737_ _08734_ vssd1 vssd1 vccd1 vccd1 _08738_ sky130_fd_sc_hd__a211o_1
X_11789_ _06758_ _06760_ net569 vssd1 vssd1 vccd1 vccd1 _06761_ sky130_fd_sc_hd__mux2_1
XANTENNA__12347__A net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17516__B1 net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19104_ clknet_leaf_0_clk img_gen.tracker.next_frame\[542\] net1240 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[542\] sky130_fd_sc_hd__dfrtp_1
X_16316_ net369 _01982_ _01986_ net368 vssd1 vssd1 vccd1 vccd1 _01995_ sky130_fd_sc_hd__o211a_1
XFILLER_0_12_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13528_ net226 _07921_ _07922_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[563\]
+ sky130_fd_sc_hd__o21bai_1
XANTENNA__11800__A1 net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17296_ ag2.body\[345\] net734 vssd1 vssd1 vccd1 vccd1 _02975_ sky130_fd_sc_hd__nor2_1
XFILLER_0_82_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_2100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19035_ clknet_leaf_6_clk img_gen.tracker.next_frame\[473\] net1264 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[473\] sky130_fd_sc_hd__dfrtp_1
X_16247_ _01922_ _01925_ net369 vssd1 vssd1 vccd1 vccd1 _01926_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_557 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16253__S net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14562__A net1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13459_ net281 _07894_ _07895_ net1709 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[521\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA_max_cap358_X net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_71_clk_A clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16178_ obsg2.obstacleArray\[52\] obsg2.obstacleArray\[53\] net424 vssd1 vssd1 vccd1
+ vccd1 _01857_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11564__B1 net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15129_ control.body\[880\] net107 _01566_ control.body\[872\] vssd1 vssd1 vccd1
+ vccd1 _00450_ sky130_fd_sc_hd__a22o_1
XFILLER_0_121_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12108__A2 net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13305__A1 net235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09943__X _04916_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12513__C net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19937_ clknet_leaf_47_clk _00881_ net1375 vssd1 vssd1 vccd1 vccd1 ag2.body\[463\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__11316__B1 _06288_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17047__A2 net864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_86_clk_A clknet_4_12__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19868_ clknet_leaf_94_clk _00812_ net1440 vssd1 vssd1 vccd1 vccd1 ag2.body\[522\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_120_1492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09621_ _04591_ _04592_ _04593_ vssd1 vssd1 vccd1 vccd1 _04594_ sky130_fd_sc_hd__or3_1
X_18819_ clknet_leaf_2_clk img_gen.tracker.next_frame\[257\] net1249 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[257\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__09822__C _04792_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19799_ clknet_leaf_128_clk _00743_ net1328 vssd1 vssd1 vccd1 vccd1 ag2.body\[597\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__16001__B net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14805__A1 net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14805__B2 net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1229 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09552_ net1119 control.body\[724\] vssd1 vssd1 vccd1 vccd1 _04525_ sky130_fd_sc_hd__xor2_1
XANTENNA__16936__B net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09483_ _04448_ _04450_ _04454_ _04455_ vssd1 vssd1 vccd1 vccd1 _04456_ sky130_fd_sc_hd__or4_1
XFILLER_0_52_1527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14737__A net1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout255_A net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18990__CLK clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18209__A net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_860 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_144_clk_A clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_24_clk_A clknet_4_6__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout422_A net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1164_A net1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_1472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20574_ clknet_leaf_106_clk _01432_ _00038_ vssd1 vssd1 vccd1 vccd1 sound_gen.dac1.dacCount\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__16191__C1 _01729_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout210_X net210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1331_A net1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout308_X net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09748__B1 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_39_clk_A clknet_4_5__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14903__C net66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout791_A net797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14191__B ag2.body\[163\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19496__CLK clknet_leaf_113_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17783__A net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13088__A net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1217_X net1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1307 net1309 vssd1 vssd1 vccd1 vccd1 net1307 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_121_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout320 _08060_ vssd1 vssd1 vccd1 vccd1 net320 sky130_fd_sc_hd__buf_2
XANTENNA__13847__A2 net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout677_X net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1318 net1320 vssd1 vssd1 vccd1 vccd1 net1318 sky130_fd_sc_hd__clkbuf_4
Xfanout331 _07424_ vssd1 vssd1 vccd1 vccd1 net331 sky130_fd_sc_hd__clkbuf_2
Xfanout1329 net1330 vssd1 vssd1 vccd1 vccd1 net1329 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_61_1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17038__A2 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout342 _07308_ vssd1 vssd1 vccd1 vccd1 net342 sky130_fd_sc_hd__clkbuf_4
Xfanout353 net354 vssd1 vssd1 vccd1 vccd1 net353 sky130_fd_sc_hd__buf_1
XFILLER_0_96_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout364 _02068_ vssd1 vssd1 vccd1 vccd1 net364 sky130_fd_sc_hd__buf_4
XANTENNA_fanout70_A net91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout375 _01740_ vssd1 vssd1 vccd1 vccd1 net375 sky130_fd_sc_hd__clkbuf_4
X_20008_ clknet_leaf_59_clk _00952_ net1471 vssd1 vssd1 vccd1 vccd1 ag2.body\[390\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__09920__B1 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout386 _06676_ vssd1 vssd1 vccd1 vccd1 net386 sky130_fd_sc_hd__clkbuf_4
Xfanout397 net400 vssd1 vssd1 vccd1 vccd1 net397 sky130_fd_sc_hd__clkbuf_4
X_09819_ _04632_ _04791_ vssd1 vssd1 vccd1 vccd1 _04792_ sky130_fd_sc_hd__or2_4
XFILLER_0_92_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17007__B net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout844_X net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1329 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11336__A net1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12830_ net675 _07616_ vssd1 vssd1 vccd1 vccd1 _07617_ sky130_fd_sc_hd__nor2_1
XANTENNA__11086__A2 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12761_ net329 _07479_ vssd1 vssd1 vccd1 vccd1 _07584_ sky130_fd_sc_hd__nand2_2
XANTENNA__16338__S net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14647__A net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11623__X _06596_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10294__B1 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14500_ net975 _04088_ _04089_ net1010 _08658_ vssd1 vssd1 vccd1 vccd1 _08661_ sky130_fd_sc_hd__a221o_1
XFILLER_0_56_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11712_ img_gen.tracker.frame\[326\] net619 vssd1 vssd1 vccd1 vccd1 _06684_ sky130_fd_sc_hd__or2_1
X_12692_ net344 _07421_ net329 vssd1 vssd1 vccd1 vccd1 _07551_ sky130_fd_sc_hd__and3_2
X_15480_ ag2.body\[568\] net112 _01605_ ag2.body\[560\] vssd1 vssd1 vccd1 vccd1 _00762_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_83_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11643_ obsg2.obstacleArray\[128\] obsg2.obstacleArray\[132\] net513 vssd1 vssd1
+ vccd1 vccd1 _06616_ sky130_fd_sc_hd__mux2_1
X_14431_ net1007 ag2.body\[559\] vssd1 vssd1 vccd1 vccd1 _08592_ sky130_fd_sc_hd__xor2_1
XFILLER_0_65_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17150_ ag2.body\[609\] net868 vssd1 vssd1 vccd1 vccd1 _02829_ sky130_fd_sc_hd__or2_1
XFILLER_0_65_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11574_ obsg2.obstacleArray\[80\] obsg2.obstacleArray\[84\] net514 vssd1 vssd1 vccd1
+ vccd1 _06547_ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14362_ net987 ag2.body\[601\] vssd1 vssd1 vccd1 vccd1 _08523_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_80_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18171__B1 net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16101_ _01778_ _01779_ net374 vssd1 vssd1 vccd1 vccd1 _01780_ sky130_fd_sc_hd__mux2_1
XFILLER_0_91_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11794__B1 net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10525_ net1058 control.body\[919\] vssd1 vssd1 vccd1 vccd1 _05498_ sky130_fd_sc_hd__xor2_1
XANTENNA__18713__CLK clknet_leaf_144_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13313_ _07490_ net304 vssd1 vssd1 vccd1 vccd1 _07839_ sky130_fd_sc_hd__nor2_1
X_14293_ net970 _04169_ ag2.body\[479\] net791 _08453_ vssd1 vssd1 vccd1 vccd1 _08454_
+ sky130_fd_sc_hd__a221o_1
X_17081_ ag2.body\[197\] net947 vssd1 vssd1 vccd1 vccd1 _02760_ sky130_fd_sc_hd__nand2_1
XFILLER_0_135_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16073__S net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14382__A net992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xmax_cap509 _06465_ vssd1 vssd1 vccd1 vccd1 net509 sky130_fd_sc_hd__buf_4
X_16032_ net539 _01681_ vssd1 vssd1 vccd1 vccd1 _01711_ sky130_fd_sc_hd__xor2_1
X_13244_ net259 net314 _07435_ _07810_ net1744 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[391\]
+ sky130_fd_sc_hd__a32o_1
X_10456_ _05425_ _05426_ _05427_ _05428_ vssd1 vssd1 vccd1 vccd1 _05429_ sky130_fd_sc_hd__a22o_1
XANTENNA__10349__B2 ag2.body\[288\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12614__B net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13175_ net667 _07778_ vssd1 vssd1 vccd1 vccd1 _07779_ sky130_fd_sc_hd__nor2_1
X_10387_ net1160 control.body\[1059\] vssd1 vssd1 vccd1 vccd1 _05360_ sky130_fd_sc_hd__xor2_1
XANTENNA__10415__A _05301_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12126_ img_gen.tracker.frame\[528\] net613 net596 img_gen.tracker.frame\[531\] _07097_
+ vssd1 vssd1 vccd1 vccd1 _07098_ sky130_fd_sc_hd__o221a_1
X_17983_ obsg2.obstacleArray\[16\] _03602_ net533 vssd1 vssd1 vccd1 vccd1 _01267_
+ sky130_fd_sc_hd__o21a_1
XANTENNA__17029__A2 net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19722_ clknet_leaf_128_clk _00666_ net1308 vssd1 vssd1 vccd1 vccd1 control.body\[664\]
+ sky130_fd_sc_hd__dfrtp_1
X_12057_ img_gen.tracker.frame\[84\] net630 net595 img_gen.tracker.frame\[93\] vssd1
+ vssd1 vccd1 vccd1 _07029_ sky130_fd_sc_hd__a22o_1
X_16934_ ag2.body\[521\] net873 vssd1 vssd1 vccd1 vccd1 _02613_ sky130_fd_sc_hd__nand2_1
XFILLER_0_74_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16237__B1 net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11008_ net1182 control.body\[1082\] vssd1 vssd1 vccd1 vccd1 _05981_ sky130_fd_sc_hd__xnor2_1
XANTENNA__15767__A_N _04897_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19653_ clknet_leaf_134_clk _00597_ net1308 vssd1 vssd1 vccd1 vccd1 control.body\[739\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11517__Y _06490_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16865_ _02541_ _02542_ _02543_ _02540_ vssd1 vssd1 vccd1 vccd1 _02544_ sky130_fd_sc_hd__a211o_1
XANTENNA__16788__A1 net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18604_ clknet_leaf_17_clk img_gen.tracker.next_frame\[42\] net1318 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[42\] sky130_fd_sc_hd__dfrtp_1
X_15816_ ag2.body\[275\] net205 _01642_ ag2.body\[267\] vssd1 vssd1 vccd1 vccd1 _01061_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__10150__A ag2.body\[56\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19584_ clknet_leaf_116_clk _00528_ net1385 vssd1 vssd1 vccd1 vccd1 control.body\[814\]
+ sky130_fd_sc_hd__dfrtp_1
X_16796_ net365 _02474_ vssd1 vssd1 vccd1 vccd1 _02475_ sky130_fd_sc_hd__nor2_1
XFILLER_0_88_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18535_ clknet_leaf_136_clk _00061_ net1300 vssd1 vssd1 vccd1 vccd1 img_gen.updater.commands.count\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_15747_ ag2.body\[342\] net217 _01634_ ag2.body\[334\] vssd1 vssd1 vccd1 vccd1 _01000_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_38_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12959_ net668 _07676_ vssd1 vssd1 vccd1 vccd1 _07677_ sky130_fd_sc_hd__nor2_1
XANTENNA__18029__A net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14557__A net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13461__A net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17201__A2 net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19369__CLK clknet_leaf_102_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18466_ _04261_ net737 net732 vssd1 vssd1 vccd1 vccd1 _03953_ sky130_fd_sc_hd__or3_1
X_15678_ ag2.body\[392\] net141 _01627_ ag2.body\[384\] vssd1 vssd1 vccd1 vccd1 _00938_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_114_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17417_ _03094_ _03095_ vssd1 vssd1 vccd1 vccd1 _03096_ sky130_fd_sc_hd__nand2b_1
XANTENNA__13180__B net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14629_ net1016 ag2.body\[470\] vssd1 vssd1 vccd1 vccd1 _08790_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_51_1571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14844__X _01515_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18397_ _03789_ _03873_ vssd1 vssd1 vccd1 vccd1 _03887_ sky130_fd_sc_hd__nor2_1
XFILLER_0_90_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10037__B1 _04416_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17348_ _03012_ _03014_ _03026_ vssd1 vssd1 vccd1 vccd1 _03027_ sky130_fd_sc_hd__mux2_1
XANTENNA__14971__B1 net51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11785__B1 net598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14292__A net1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17279_ ag2.body\[553\] net731 net689 ag2.body\[559\] _02957_ vssd1 vssd1 vccd1 vccd1
+ _02958_ sky130_fd_sc_hd__a221o_1
XFILLER_0_86_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19018_ clknet_leaf_6_clk img_gen.tracker.next_frame\[456\] net1246 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[456\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_wire478_X net478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14723__B1 _08883_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20290_ clknet_leaf_35_clk control.divider.next_count\[11\] net1350 vssd1 vssd1 vccd1
+ vccd1 control.divider.count\[11\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17268__A2 net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09673__X _04646_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08983_ ag2.body\[77\] vssd1 vssd1 vccd1 vccd1 _04008_ sky130_fd_sc_hd__inv_2
XANTENNA__12811__Y _07607_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1576 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11662__B1_N net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16012__A net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12540__A net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09604_ net1073 control.body\[638\] vssd1 vssd1 vccd1 vccd1 _04577_ sky130_fd_sc_hd__xor2_1
XFILLER_0_93_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09535_ control.body\[1026\] net1182 vssd1 vssd1 vccd1 vccd1 _04508_ sky130_fd_sc_hd__and2b_1
XANTENNA__17728__B1 net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14467__A net1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout258_X net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1379_A net1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09466_ ag2.body\[377\] net778 net754 ag2.body\[381\] vssd1 vssd1 vccd1 vccd1 _04439_
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_133_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14186__B ag2.body\[166\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09681__A2 net1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18736__CLK clknet_leaf_142_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09397_ net1641 _04344_ _04382_ vssd1 vssd1 vccd1 vccd1 _01404_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout425_X net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout804_A net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1167_X net1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20626_ sound_gen.dac1.dacCount\[4\] vssd1 vssd1 vccd1 vccd1 net13 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_34_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14962__B1 _01547_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17497__B net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11776__B1 net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20557_ clknet_leaf_105_clk _01422_ _00031_ vssd1 vssd1 vccd1 vccd1 sound_gen.osc1.stayCount\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_7_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12715__A net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10310_ _04603_ _04640_ _04572_ vssd1 vssd1 vccd1 vccd1 _05283_ sky130_fd_sc_hd__o21ai_2
XANTENNA__14714__B1 ag2.body\[342\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11290_ _06257_ _06258_ _06261_ _06262_ vssd1 vssd1 vccd1 vccd1 _06263_ sky130_fd_sc_hd__a22o_1
X_20488_ clknet_leaf_38_clk _01375_ net1354 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[124\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__11528__B1 net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout794_X net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10241_ ag2.body\[320\] net1236 vssd1 vssd1 vccd1 vccd1 _05214_ sky130_fd_sc_hd__or2_1
XFILLER_0_104_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17717__S net378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14930__A _05364_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16467__B1 net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09583__X _04556_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13817__Y _08114_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10172_ _05120_ _05130_ _05132_ _05144_ vssd1 vssd1 vccd1 vccd1 _05145_ sky130_fd_sc_hd__o31a_1
XANTENNA_fanout961_X net961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_3690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1104 net1106 vssd1 vssd1 vccd1 vccd1 net1104 sky130_fd_sc_hd__clkbuf_8
Xfanout1115 net1117 vssd1 vssd1 vccd1 vccd1 net1115 sky130_fd_sc_hd__buf_4
Xfanout1126 net1129 vssd1 vssd1 vccd1 vccd1 net1126 sky130_fd_sc_hd__clkbuf_4
XANTENNA__18208__A1 net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1137 net1143 vssd1 vssd1 vccd1 vccd1 net1137 sky130_fd_sc_hd__clkbuf_4
X_14980_ control.body\[1019\] net158 _01550_ control.body\[1011\] vssd1 vssd1 vccd1
+ vccd1 _00317_ sky130_fd_sc_hd__a22o_1
XANTENNA__10522__X _05495_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout150 net154 vssd1 vssd1 vccd1 vccd1 net150 sky130_fd_sc_hd__clkbuf_2
Xfanout1148 net1151 vssd1 vssd1 vccd1 vccd1 net1148 sky130_fd_sc_hd__buf_4
Xfanout1159 net1161 vssd1 vssd1 vccd1 vccd1 net1159 sky130_fd_sc_hd__clkbuf_4
Xfanout161 net162 vssd1 vssd1 vccd1 vccd1 net161 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_96_1240 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout172 net174 vssd1 vssd1 vccd1 vccd1 net172 sky130_fd_sc_hd__buf_2
X_13931_ ag2.body\[74\] net185 _08153_ ag2.body\[66\] vssd1 vssd1 vccd1 vccd1 _00155_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11926__S1 net1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout183 net219 vssd1 vssd1 vccd1 vccd1 net183 sky130_fd_sc_hd__buf_4
Xfanout194 net196 vssd1 vssd1 vccd1 vccd1 net194 sky130_fd_sc_hd__clkbuf_2
XANTENNA__10503__A1 _04446_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11066__A _06028_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16650_ obsg2.obstacleArray\[6\] net446 vssd1 vssd1 vccd1 vccd1 _02329_ sky130_fd_sc_hd__or2_1
XANTENNA__12600__D _07312_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13862_ net325 net323 vssd1 vssd1 vccd1 vccd1 _08136_ sky130_fd_sc_hd__or2_1
XFILLER_0_44_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15601_ ag2.body\[467\] net121 _01619_ ag2.body\[459\] vssd1 vssd1 vccd1 vccd1 _00869_
+ sky130_fd_sc_hd__a22o_1
X_12813_ net669 _07608_ vssd1 vssd1 vccd1 vccd1 _07609_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_2_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16581_ net396 _02259_ _02258_ net361 vssd1 vssd1 vccd1 vccd1 _02260_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_104_3483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14377__A net1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_240 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13793_ _08099_ vssd1 vssd1 vccd1 vccd1 _08100_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_104_3494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18320_ _03815_ vssd1 vssd1 vccd1 vccd1 _03816_ sky130_fd_sc_hd__inv_2
XFILLER_0_70_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__20369__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15532_ ag2.body\[535\] net159 _01610_ ag2.body\[527\] vssd1 vssd1 vccd1 vccd1 _00809_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_100_3358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12744_ net305 _07575_ vssd1 vssd1 vccd1 vccd1 _07576_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_100_3369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1588 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18251_ obsg2.obstacleArray\[122\] _03764_ net525 vssd1 vssd1 vccd1 vccd1 _01373_
+ sky130_fd_sc_hd__o21a_1
X_15463_ ag2.body\[585\] net90 _01603_ ag2.body\[577\] vssd1 vssd1 vccd1 vccd1 _00747_
+ sky130_fd_sc_hd__a22o_1
X_12675_ net339 net315 _07542_ vssd1 vssd1 vccd1 vccd1 _07543_ sky130_fd_sc_hd__nor3_2
X_17202_ ag2.body\[177\] net870 vssd1 vssd1 vccd1 vccd1 _02881_ sky130_fd_sc_hd__xor2_1
XFILLER_0_127_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14414_ net1031 ag2.body\[533\] vssd1 vssd1 vccd1 vccd1 _08575_ sky130_fd_sc_hd__xnor2_1
X_18182_ _03622_ net36 vssd1 vssd1 vccd1 vccd1 _03730_ sky130_fd_sc_hd__nor2_1
X_11626_ obsg2.obstacleArray\[47\] net631 net510 obsg2.obstacleArray\[43\] net1125
+ vssd1 vssd1 vccd1 vccd1 _06599_ sky130_fd_sc_hd__o221a_1
XANTENNA__14953__B1 _01546_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15479__Y _01605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15394_ net2229 net82 _01596_ net2360 vssd1 vssd1 vccd1 vccd1 _00685_ sky130_fd_sc_hd__a22o_1
XANTENNA__11767__B1 net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_117_3877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17133_ ag2.body\[518\] net942 vssd1 vssd1 vccd1 vccd1 _02812_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_117_3888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14345_ net817 ag2.body\[611\] ag2.body\[615\] net790 _08501_ vssd1 vssd1 vccd1 vccd1
+ _08506_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_117_3899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11557_ obsg2.obstacleArray\[64\] obsg2.obstacleArray\[68\] net513 vssd1 vssd1 vccd1
+ vccd1 _06530_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13508__A1 net250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_1386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17064_ ag2.body\[25\] net868 vssd1 vssd1 vccd1 vccd1 _02743_ sky130_fd_sc_hd__or2_1
X_10508_ net1230 control.body\[976\] vssd1 vssd1 vccd1 vccd1 _05481_ sky130_fd_sc_hd__xnor2_1
Xhold609 control.body\[773\] vssd1 vssd1 vccd1 vccd1 net2171 sky130_fd_sc_hd__dlygate4sd3_1
X_14276_ _08431_ _08434_ _08435_ _08436_ vssd1 vssd1 vccd1 vccd1 _08437_ sky130_fd_sc_hd__or4_2
X_11488_ net1197 net1078 vssd1 vssd1 vccd1 vccd1 _06461_ sky130_fd_sc_hd__xor2_2
X_16015_ _01692_ _01693_ _01690_ vssd1 vssd1 vccd1 vccd1 _01694_ sky130_fd_sc_hd__o21ai_1
XANTENNA__14181__A1 net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10439_ net1229 control.body\[928\] vssd1 vssd1 vccd1 vccd1 _05412_ sky130_fd_sc_hd__xnor2_1
X_13227_ net239 _07802_ _07803_ net1906 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[381\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_21_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18447__A1 _05075_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14181__B2 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11534__A3 net1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13158_ net667 _07770_ vssd1 vssd1 vccd1 vccd1 _07771_ sky130_fd_sc_hd__nor2_1
XFILLER_0_0_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17960__A_N net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12109_ net1215 net1190 img_gen.tracker.frame\[189\] vssd1 vssd1 vccd1 vccd1 _07081_
+ sky130_fd_sc_hd__and3_1
XANTENNA__13456__A net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17966_ net298 _03589_ vssd1 vssd1 vccd1 vccd1 _03590_ sky130_fd_sc_hd__nand2_1
X_13089_ net685 _07737_ vssd1 vssd1 vccd1 vccd1 _07738_ sky130_fd_sc_hd__nor2_1
XFILLER_0_85_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10799__B net1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19705_ clknet_leaf_136_clk _00649_ net1301 vssd1 vssd1 vccd1 vccd1 control.body\[695\]
+ sky130_fd_sc_hd__dfrtp_1
X_16917_ ag2.body\[562\] net859 vssd1 vssd1 vccd1 vccd1 _02596_ sky130_fd_sc_hd__xnor2_1
XANTENNA__12495__A1 net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17897_ net433 _02054_ vssd1 vssd1 vccd1 vccd1 _03533_ sky130_fd_sc_hd__nor2_4
XPHY_EDGE_ROW_108_Left_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14839__X _01510_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16848_ ag2.body\[172\] net960 vssd1 vssd1 vccd1 vccd1 _02527_ sky130_fd_sc_hd__or2_1
XANTENNA__19145__RESET_B net1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19636_ clknet_leaf_123_clk _00580_ net1405 vssd1 vssd1 vccd1 vccd1 control.body\[754\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_0_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19567_ clknet_leaf_116_clk _00511_ net1387 vssd1 vssd1 vccd1 vccd1 control.body\[829\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__15390__B net63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18759__CLK clknet_leaf_15_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16779_ _02389_ _02392_ net432 vssd1 vssd1 vccd1 vccd1 _02458_ sky130_fd_sc_hd__mux2_1
XANTENNA__14287__A net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13191__A net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09320_ _04312_ _04319_ _04320_ net272 net2348 vssd1 vssd1 vccd1 vccd1 _01436_ sky130_fd_sc_hd__a32o_1
X_18518_ net1512 net1506 vssd1 vssd1 vccd1 vccd1 _00049_ sky130_fd_sc_hd__or2_1
X_19498_ clknet_leaf_113_clk _00442_ net1401 vssd1 vssd1 vccd1 vccd1 control.body\[888\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11040__A_N net1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09251_ control.detect3.Q\[0\] vssd1 vssd1 vccd1 vccd1 _04276_ sky130_fd_sc_hd__inv_2
XFILLER_0_88_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15197__B1 _01573_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18449_ _04642_ _03834_ _03891_ _03937_ vssd1 vssd1 vccd1 vccd1 _03938_ sky130_fd_sc_hd__a211o_1
XANTENNA__11423__B control.body\[848\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09182_ ag2.body\[562\] vssd1 vssd1 vccd1 vccd1 _04207_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_117_Left_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20411_ clknet_leaf_32_clk _01298_ net1345 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[47\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__18206__B net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17489__A2 net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_133_4380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_721 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout120_A net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_133_4391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout218_A net219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_6__f_clk clknet_3_3_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_6__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_82_1306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16697__B1 net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_1328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20342_ clknet_leaf_140_clk _01233_ net1292 vssd1 vssd1 vccd1 vccd1 img_gen.updater.commands.rR1.rainbowRNG\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__20525__Q control.body_update.curr_length\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20273_ clknet_leaf_37_clk net4 net1353 vssd1 vssd1 vccd1 vccd1 control.button3.Q\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_101_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17764__C _02742_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_4__f_clk_X clknet_4_4__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1127_A net1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19915__RESET_B net1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout587_A net589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17661__A2 net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_1991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08966_ ag2.body\[49\] vssd1 vssd1 vccd1 vccd1 _03991_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_127_4184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_126_Left_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_127_4195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20260__Q ag2.body\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13085__B net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout375_X net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout754_A _04232_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1496_A net1499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_95_clk clknet_4_11__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_95_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_93_1424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10497__B1 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17413__A2 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20511__CLK clknet_leaf_113_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20473__RESET_B net1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout921_A net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout542_X net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11614__A net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_722 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09518_ net896 net900 net890 vssd1 vssd1 vccd1 vccd1 _04491_ sky130_fd_sc_hd__a21oi_2
X_10790_ _05753_ _05754_ _05758_ _05759_ _05755_ vssd1 vssd1 vccd1 vccd1 _05763_ sky130_fd_sc_hd__a221o_1
XFILLER_0_116_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_1491 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09449_ net920 net916 vssd1 vssd1 vccd1 vccd1 _04422_ sky130_fd_sc_hd__and2_1
XANTENNA__14484__X _08645_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout807_X net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_1187 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1451_X net1451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_135_Left_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17939__C net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_427 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12460_ _07284_ _07294_ _07418_ net687 vssd1 vssd1 vccd1 vccd1 img_gen.dcx sky130_fd_sc_hd__a22o_1
XFILLER_0_81_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_10_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11411_ _06378_ _06381_ _06382_ _06383_ vssd1 vssd1 vccd1 vccd1 _06384_ sky130_fd_sc_hd__or4_1
X_20609_ net1541 vssd1 vssd1 vccd1 vccd1 gpio_oeb[21] sky130_fd_sc_hd__buf_2
X_12391_ net1217 _07355_ vssd1 vssd1 vccd1 vccd1 _07356_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_10_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12410__A1 net1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11342_ ag2.body\[442\] net1178 vssd1 vssd1 vccd1 vccd1 _06315_ sky130_fd_sc_hd__xor2_1
X_14130_ net833 ag2.body\[369\] ag2.body\[370\] net826 _08290_ vssd1 vssd1 vccd1 vccd1
+ _08291_ sky130_fd_sc_hd__a221o_1
XFILLER_0_65_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_112_3730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_3741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17955__B net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_3752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11273_ ag2.body\[126\] net1090 vssd1 vssd1 vccd1 vccd1 _06246_ sky130_fd_sc_hd__or2_1
X_14061_ net832 ag2.body\[33\] ag2.body\[39\] net790 vssd1 vssd1 vccd1 vccd1 _08222_
+ sky130_fd_sc_hd__o22a_1
XANTENNA__15360__B1 _01592_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14793__A1_N net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14660__A net1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18132__A net41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13012_ _07701_ net262 _07699_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[268\]
+ sky130_fd_sc_hd__mux2_1
X_10224_ _05193_ _05194_ _05195_ _05196_ vssd1 vssd1 vccd1 vccd1 _05197_ sky130_fd_sc_hd__a22o_1
X_17820_ _03481_ _03484_ _03483_ vssd1 vssd1 vccd1 vccd1 _03486_ sky130_fd_sc_hd__a21oi_1
XANTENNA__17971__A net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10155_ _05121_ _05122_ _05126_ _05127_ vssd1 vssd1 vccd1 vccd1 _05128_ sky130_fd_sc_hd__a22o_1
XANTENNA__15112__B1 _01554_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14178__A1_N net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17652__A2 net715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16860__B1 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17751_ _02610_ _02611_ _03333_ vssd1 vssd1 vccd1 vccd1 _03430_ sky130_fd_sc_hd__o21a_1
Xhold6 control.button1.Q\[1\] vssd1 vssd1 vccd1 vccd1 net1568 sky130_fd_sc_hd__dlygate4sd3_1
X_10086_ net1075 control.body\[798\] vssd1 vssd1 vccd1 vccd1 _05059_ sky130_fd_sc_hd__or2_1
X_14963_ net2540 net159 _01547_ control.body\[1029\] vssd1 vssd1 vccd1 vccd1 _00303_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12477__A1 _07425_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_106_3545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_505 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_86_clk clknet_4_12__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_86_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_136_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16702_ obsg2.obstacleArray\[87\] net503 net493 obsg2.obstacleArray\[84\] vssd1 vssd1
+ vccd1 vccd1 _02381_ sky130_fd_sc_hd__a22o_1
XANTENNA__18901__CLK clknet_leaf_144_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_3556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13914_ ag2.body\[59\] net129 _08151_ ag2.body\[51\] vssd1 vssd1 vccd1 vccd1 _00140_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__10488__B1 net1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_106_3567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17682_ ag2.body\[478\] net937 vssd1 vssd1 vccd1 vccd1 _03361_ sky130_fd_sc_hd__xor2_1
XANTENNA__20191__CLK clknet_leaf_88_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14894_ net635 _01536_ vssd1 vssd1 vccd1 vccd1 _01540_ sky130_fd_sc_hd__and2b_2
XFILLER_0_76_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19421_ clknet_leaf_107_clk _00365_ net1434 vssd1 vssd1 vccd1 vccd1 control.body\[971\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16633_ net395 _02311_ net359 vssd1 vssd1 vccd1 vccd1 _02312_ sky130_fd_sc_hd__a21o_1
X_13845_ ag2.body\[9\] net127 _08133_ net1043 vssd1 vssd1 vccd1 vccd1 _00089_ sky130_fd_sc_hd__a22o_1
XFILLER_0_85_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__20143__RESET_B net1451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19352_ clknet_leaf_101_clk net2514 net1439 vssd1 vssd1 vccd1 vccd1 control.body\[1046\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_4_15__f_clk_X clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16564_ _02207_ _02242_ vssd1 vssd1 vccd1 vccd1 _02243_ sky130_fd_sc_hd__and2_1
X_13776_ _08071_ _08085_ _08087_ vssd1 vssd1 vccd1 vccd1 _00066_ sky130_fd_sc_hd__and3_1
X_10988_ _05952_ _05955_ _05957_ _05958_ vssd1 vssd1 vccd1 vccd1 _05961_ sky130_fd_sc_hd__or4_1
XFILLER_0_69_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_80_2752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18303_ net325 net323 _03798_ _03793_ net321 vssd1 vssd1 vccd1 vccd1 _03799_ sky130_fd_sc_hd__a311oi_2
XANTENNA__11243__B net1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15515_ _05303_ net65 vssd1 vssd1 vccd1 vccd1 _01609_ sky130_fd_sc_hd__and2_2
XTAP_TAPCELL_ROW_80_2763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12727_ net305 _07567_ vssd1 vssd1 vccd1 vccd1 _07568_ sky130_fd_sc_hd__nor2_1
X_19283_ clknet_leaf_98_clk _00227_ net1446 vssd1 vssd1 vccd1 vccd1 control.body\[1105\]
+ sky130_fd_sc_hd__dfrtp_1
X_16495_ net400 _02173_ _02172_ net367 vssd1 vssd1 vccd1 vccd1 _02174_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_119_3939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_2774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_939 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_2173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18234_ _03675_ net35 vssd1 vssd1 vccd1 vccd1 _03756_ sky130_fd_sc_hd__nor2_1
XFILLER_0_26_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_2184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14926__B1 _01543_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15446_ ag2.body\[602\] net86 _01601_ ag2.body\[594\] vssd1 vssd1 vccd1 vccd1 _00732_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_61_2195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12658_ net240 _07533_ _07534_ net1890 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[81\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_112_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18026__B net38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14554__B ag2.body\[67\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11609_ net505 _06580_ _06581_ net475 vssd1 vssd1 vccd1 vccd1 _06582_ sky130_fd_sc_hd__o31a_1
X_18165_ net518 _03721_ vssd1 vssd1 vccd1 vccd1 _01330_ sky130_fd_sc_hd__nor2_1
XANTENNA__19407__CLK clknet_leaf_103_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15002__Y _01552_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15377_ net2396 net82 _01594_ control.body\[660\] vssd1 vssd1 vccd1 vccd1 _00670_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12355__A net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12589_ _07431_ _07494_ net644 vssd1 vssd1 vccd1 vccd1 _07496_ sky130_fd_sc_hd__o21a_1
XFILLER_0_128_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_10_clk clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_10_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_105_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17116_ ag2.body\[536\] net739 net735 ag2.body\[537\] vssd1 vssd1 vccd1 vccd1 _02795_
+ sky130_fd_sc_hd__a2bb2o_1
X_14328_ _08487_ _08488_ vssd1 vssd1 vccd1 vccd1 _08489_ sky130_fd_sc_hd__nand2_1
XFILLER_0_83_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18096_ net44 _03679_ vssd1 vssd1 vccd1 vccd1 _03680_ sky130_fd_sc_hd__nor2_1
XFILLER_0_40_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16143__A2 net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_2692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold406 img_gen.tracker.frame\[105\] vssd1 vssd1 vccd1 vccd1 net1968 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10963__A1 _05922_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold417 img_gen.tracker.frame\[503\] vssd1 vssd1 vccd1 vccd1 net1979 sky130_fd_sc_hd__dlygate4sd3_1
Xhold428 img_gen.tracker.frame\[180\] vssd1 vssd1 vccd1 vccd1 net1990 sky130_fd_sc_hd__dlygate4sd3_1
X_17047_ _04087_ net864 net933 _04089_ _02723_ vssd1 vssd1 vccd1 vccd1 _02726_ sky130_fd_sc_hd__a221o_1
Xhold439 img_gen.tracker.frame\[342\] vssd1 vssd1 vccd1 vccd1 net2001 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12505__D net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16261__S net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14259_ net1004 _04003_ ag2.body\[74\] net829 vssd1 vssd1 vccd1 vccd1 _08420_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_74_2567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_1346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_74_2578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_74_2589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout908 control.body_update.curr_length\[4\] vssd1 vssd1 vccd1 vccd1 net908 sky130_fd_sc_hd__buf_4
XANTENNA__11912__B1 net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout919 net920 vssd1 vssd1 vccd1 vccd1 net919 sky130_fd_sc_hd__buf_4
XFILLER_0_29_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13186__A net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16300__C1 _01918_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10603__A net1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_14__f_clk clknet_3_7_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_14__leaf_clk
+ sky130_fd_sc_hd__clkbuf_16
X_18998_ clknet_leaf_2_clk img_gen.tracker.next_frame\[436\] net1248 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[436\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__13665__B1 net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17949_ net380 net462 net495 net490 vssd1 vssd1 vccd1 vccd1 _03577_ sky130_fd_sc_hd__and4_2
Xclkbuf_leaf_77_clk clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_77_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_20_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10322__B net1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1490 net1492 vssd1 vssd1 vccd1 vccd1 net1490 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_75_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09884__A2 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1608 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19619_ clknet_leaf_119_clk _00563_ net1391 vssd1 vssd1 vccd1 vccd1 control.body\[769\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11691__A2 net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16944__B net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09303_ sound_gen.osc1.count\[3\] _04321_ vssd1 vssd1 vccd1 vccd1 _04323_ sky130_fd_sc_hd__and2_1
XANTENNA__11153__B net1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16367__C1 net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_135_4431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16436__S net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14745__A net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_4442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout335_A _07423_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_135_4453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1077_A net1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09839__A net1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_3_Right_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09234_ img_gen.control.current\[1\] vssd1 vssd1 vccd1 vccd1 _04259_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_131_4306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_4317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10992__B net1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_4328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11440__Y _06413_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_1534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09165_ ag2.body\[515\] vssd1 vssd1 vccd1 vccd1 _04190_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_20_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout502_A _01708_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_1556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_983 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1244_A net1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09096_ ag2.body\[342\] vssd1 vssd1 vccd1 vccd1 _04121_ sky130_fd_sc_hd__inv_2
XFILLER_0_4_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20325_ clknet_4_7__leaf_clk _01221_ net1377 vssd1 vssd1 vccd1 vccd1 ag2.body\[6\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_114_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16171__S net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15342__B1 _01590_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14480__A net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1032_X net1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16024__X _01703_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold940 control.body\[1027\] vssd1 vssd1 vccd1 vccd1 net2502 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1411_A net1415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_90_3070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12156__B1 net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold951 control.body\[1046\] vssd1 vssd1 vccd1 vccd1 net2513 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_4246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_3081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold962 control.body\[774\] vssd1 vssd1 vccd1 vccd1 net2524 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20256_ clknet_leaf_70_clk _01200_ net1497 vssd1 vssd1 vccd1 vccd1 ag2.body\[142\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_129_4257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold973 control.body\[971\] vssd1 vssd1 vccd1 vccd1 net2535 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_4268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold984 control.body\[692\] vssd1 vssd1 vccd1 vccd1 net2546 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout871_A net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout492_X net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_1474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold995 control.body\[763\] vssd1 vssd1 vccd1 vccd1 net2557 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_53_1928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_1496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20187_ clknet_leaf_88_clk _01131_ net1454 vssd1 vssd1 vccd1 vccd1 ag2.body\[201\]
+ sky130_fd_sc_hd__dfrtp_4
X_09998_ net1144 control.body\[731\] vssd1 vssd1 vccd1 vccd1 _04971_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_34_1349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09724__D net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08949_ ag2.body\[7\] vssd1 vssd1 vccd1 vccd1 _03974_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_4_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_68_clk clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_68_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__14853__C1 _08574_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout757_X net757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1499_X net1499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09580__Y _04553_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11960_ _06723_ _06931_ vssd1 vssd1 vccd1 vccd1 _06932_ sky130_fd_sc_hd__and2_1
X_10911_ _05871_ _05883_ _05855_ _05869_ vssd1 vssd1 vccd1 vccd1 _05884_ sky130_fd_sc_hd__o211ai_1
XANTENNA__17015__B net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15948__A2 net195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11891_ net470 _06862_ _06856_ net436 vssd1 vssd1 vccd1 vccd1 _06863_ sky130_fd_sc_hd__o211a_1
XANTENNA__11682__A2 net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13630_ net2190 _07992_ _07994_ vssd1 vssd1 vccd1 vccd1 control.divider.next_count\[10\]
+ sky130_fd_sc_hd__a21oi_1
X_10842_ ag2.body\[46\] net1074 vssd1 vssd1 vccd1 vccd1 _05815_ sky130_fd_sc_hd__xor2_1
XANTENNA_fanout36_X net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11063__B net1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12631__A1 net225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13561_ ssdec1.in\[3\] _07932_ _07940_ _07941_ _07936_ vssd1 vssd1 vccd1 vccd1 net18
+ sky130_fd_sc_hd__o32a_1
XANTENNA__16346__S net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10773_ ag2.body\[219\] net1164 vssd1 vssd1 vccd1 vccd1 _05746_ sky130_fd_sc_hd__xor2_1
XANTENNA__14655__A net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18127__A net38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15300_ _04968_ _01581_ vssd1 vssd1 vccd1 vccd1 _01586_ sky130_fd_sc_hd__and2b_2
X_12512_ net575 net555 vssd1 vssd1 vccd1 vccd1 _07452_ sky130_fd_sc_hd__nand2_1
X_16280_ net420 _01958_ _01957_ net370 vssd1 vssd1 vccd1 vccd1 _01959_ sky130_fd_sc_hd__a211o_1
X_13492_ net230 _07908_ _07909_ net1789 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[540\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_125_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_97_3268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_97_3279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_114_3803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15231_ net2567 net96 _01577_ control.body\[787\] vssd1 vssd1 vccd1 vccd1 _00541_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_114_3814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17966__A net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12443_ net625 _06525_ _07379_ vssd1 vssd1 vccd1 vccd1 _07404_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_1_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1312 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15162_ net2201 net98 _01569_ control.body\[854\] vssd1 vssd1 vccd1 vccd1 _00480_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_133_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16125__A2 net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12374_ _07282_ _07330_ _07339_ _07300_ vssd1 vssd1 vccd1 vccd1 net21 sky130_fd_sc_hd__a22o_1
XANTENNA__19837__RESET_B net1414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16756__S0 net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17322__B2 net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14113_ net1015 ag2.body\[574\] vssd1 vssd1 vccd1 vccd1 _08274_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_132_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11325_ ag2.body\[554\] net1172 vssd1 vssd1 vccd1 vccd1 _06298_ sky130_fd_sc_hd__xor2_1
X_19970_ clknet_leaf_62_clk _00914_ net1470 vssd1 vssd1 vccd1 vccd1 ag2.body\[416\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__16081__S net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15093_ _04553_ net58 vssd1 vssd1 vccd1 vccd1 _01563_ sky130_fd_sc_hd__nor2_2
XANTENNA__12903__A net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20557__CLK clknet_leaf_105_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14044_ net997 ag2.body\[184\] vssd1 vssd1 vccd1 vccd1 _08205_ sky130_fd_sc_hd__xor2_1
X_18921_ clknet_leaf_145_clk img_gen.tracker.next_frame\[359\] net1253 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[359\] sky130_fd_sc_hd__dfrtp_1
X_11256_ net1202 control.body\[769\] vssd1 vssd1 vccd1 vccd1 _06229_ sky130_fd_sc_hd__xor2_1
XFILLER_0_120_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_108_3607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10207_ net750 control.body\[998\] control.body\[999\] net745 _05179_ vssd1 vssd1
+ vccd1 vccd1 _05180_ sky130_fd_sc_hd__a221o_1
XFILLER_0_101_790 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11187_ _04054_ net1224 net1081 _04058_ _06158_ vssd1 vssd1 vccd1 vccd1 _06160_ sky130_fd_sc_hd__a221o_2
XANTENNA__11113__A1_N net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18852_ clknet_leaf_18_clk img_gen.tracker.next_frame\[290\] net1324 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[290\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_108_3618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_3629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17803_ net969 net948 net939 net931 vssd1 vssd1 vccd1 vccd1 _03473_ sky130_fd_sc_hd__a31o_1
X_10138_ net1226 control.body\[816\] vssd1 vssd1 vccd1 vccd1 _05111_ sky130_fd_sc_hd__xor2_1
XANTENNA__11238__B net1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18783_ clknet_leaf_12_clk img_gen.tracker.next_frame\[221\] net1286 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[221\] sky130_fd_sc_hd__dfrtp_1
X_15995_ net1628 control.body_update.direction\[1\] net223 vssd1 vssd1 vccd1 vccd1
+ _01207_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_59_clk clknet_4_13__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_59_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__14844__C1 _01489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17734_ _03235_ _03236_ _03239_ _02917_ vssd1 vssd1 vccd1 vccd1 _03413_ sky130_fd_sc_hd__o31a_1
X_10069_ net1049 control.body\[719\] vssd1 vssd1 vccd1 vccd1 _05042_ sky130_fd_sc_hd__or2_1
X_14946_ net2298 net173 _01545_ net2420 vssd1 vssd1 vccd1 vccd1 _00288_ sky130_fd_sc_hd__a22o_1
XFILLER_0_82_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_86_2950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17665_ _03336_ _03339_ _03342_ _03343_ vssd1 vssd1 vccd1 vccd1 _03344_ sky130_fd_sc_hd__or4b_1
XTAP_TAPCELL_ROW_82_2814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_2360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15939__A2 net195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14877_ control.body\[1104\] net181 _01538_ control.body\[1096\] vssd1 vssd1 vccd1
+ vccd1 _00226_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_82_2825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_2371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16616_ obsg2.obstacleArray\[40\] obsg2.obstacleArray\[41\] net442 vssd1 vssd1 vccd1
+ vccd1 _02295_ sky130_fd_sc_hd__mux2_1
X_19404_ clknet_leaf_103_clk _00348_ net1431 vssd1 vssd1 vccd1 vccd1 control.body\[986\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11254__A net1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13828_ _04276_ control.detect3.Q\[1\] _08111_ _08113_ _08114_ vssd1 vssd1 vccd1
+ vccd1 _08125_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_58_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_63_2235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17596_ net925 net924 _03011_ _03025_ _03274_ vssd1 vssd1 vccd1 vccd1 _03275_ sky130_fd_sc_hd__o311a_1
XFILLER_0_106_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_63_2246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_2257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16547_ net390 _02218_ net361 _02225_ vssd1 vssd1 vccd1 vccd1 _02226_ sky130_fd_sc_hd__a211o_1
XFILLER_0_85_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19335_ clknet_leaf_103_clk net2168 net1431 vssd1 vssd1 vccd1 vccd1 control.body\[1061\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_31_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16349__C1 _01918_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13759_ _08075_ vssd1 vssd1 vccd1 vccd1 _08076_ sky130_fd_sc_hd__inv_2
XFILLER_0_50_1636 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14565__A net1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17010__B1 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19266_ clknet_leaf_71_clk _00210_ net1503 vssd1 vssd1 vccd1 vccd1 ag2.body\[129\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_116_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_14_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09659__A net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16478_ obsg2.obstacleArray\[32\] obsg2.obstacleArray\[33\] net452 vssd1 vssd1 vccd1
+ vccd1 _02157_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_14_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18217_ obsg2.obstacleArray\[105\] _03747_ net524 vssd1 vssd1 vccd1 vccd1 _01356_
+ sky130_fd_sc_hd__o21a_1
XANTENNA__11701__B _06644_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15429_ ag2.body\[619\] net84 _01599_ ag2.body\[611\] vssd1 vssd1 vccd1 vccd1 _00717_
+ sky130_fd_sc_hd__a22o_1
X_19197_ clknet_leaf_53_clk _00141_ net1455 vssd1 vssd1 vccd1 vccd1 ag2.body\[60\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_83_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_76_2629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_819 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18148_ net47 _03574_ _03704_ obsg2.obstacleArray\[71\] vssd1 vssd1 vccd1 vccd1 _03713_
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_14_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10936__A1 net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold203 img_gen.tracker.frame\[465\] vssd1 vssd1 vccd1 vccd1 net1765 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__19864__Q ag2.body\[534\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10317__B net1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold214 img_gen.tracker.frame\[171\] vssd1 vssd1 vccd1 vccd1 net1776 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_48_1576 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18947__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18079_ net42 _03668_ vssd1 vssd1 vccd1 vccd1 _03669_ sky130_fd_sc_hd__nor2_1
Xhold225 img_gen.tracker.frame\[410\] vssd1 vssd1 vccd1 vccd1 net1787 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12813__A net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold236 img_gen.tracker.frame\[417\] vssd1 vssd1 vccd1 vccd1 net1798 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12138__B1 net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold247 img_gen.tracker.frame\[222\] vssd1 vssd1 vccd1 vccd1 net1809 sky130_fd_sc_hd__dlygate4sd3_1
Xhold258 img_gen.tracker.frame\[411\] vssd1 vssd1 vccd1 vccd1 net1820 sky130_fd_sc_hd__dlygate4sd3_1
X_20110_ clknet_leaf_80_clk _01054_ net1487 vssd1 vssd1 vccd1 vccd1 ag2.body\[284\]
+ sky130_fd_sc_hd__dfrtp_4
X_09921_ ag2.body\[316\] net764 net1066 _04108_ vssd1 vssd1 vccd1 vccd1 _04894_ sky130_fd_sc_hd__a22o_1
Xhold269 img_gen.tracker.frame\[162\] vssd1 vssd1 vccd1 vccd1 net1831 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12689__A1 net238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout705 _04267_ vssd1 vssd1 vccd1 vccd1 net705 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12532__B net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20041_ clknet_leaf_67_clk _00985_ net1473 vssd1 vssd1 vccd1 vccd1 ag2.body\[359\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_106_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout716 _04265_ vssd1 vssd1 vccd1 vccd1 net716 sky130_fd_sc_hd__buf_4
Xfanout727 net729 vssd1 vssd1 vccd1 vccd1 net727 sky130_fd_sc_hd__buf_4
XANTENNA__19160__RESET_B net1403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09852_ net1161 control.body\[971\] vssd1 vssd1 vccd1 vccd1 _04825_ sky130_fd_sc_hd__xor2_1
Xfanout738 _04262_ vssd1 vssd1 vccd1 vccd1 net738 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_124_4110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13347__C _07813_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout749 _04233_ vssd1 vssd1 vccd1 vccd1 net749 sky130_fd_sc_hd__clkbuf_4
XANTENNA__16939__B net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14008__A1_N net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09783_ net1161 control.body\[947\] vssd1 vssd1 vccd1 vccd1 _04756_ sky130_fd_sc_hd__xor2_1
XANTENNA__10052__B net1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout285_A _07335_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_1530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11113__B2 net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12861__A1 net240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout452_A net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_1438 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1194_A net1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_137_4504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_137_4515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_46_1721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout240_X net240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14475__A net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1361_A net1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout717_A _04265_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_27_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout338_X net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17001__B1 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_42_1618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1459_A net1461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09217_ control.body\[794\] vssd1 vssd1 vccd1 vccd1 _04242_ sky130_fd_sc_hd__inv_2
XANTENNA__17786__A net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout505_X net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10508__A net1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11315__C_N _04985_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_3121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_994 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_3132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11719__A3 _06671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09148_ ag2.body\[480\] vssd1 vssd1 vccd1 vccd1 _04173_ sky130_fd_sc_hd__inv_2
XANTENNA__19930__RESET_B net1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_3143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10927__A1 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10227__B net1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09079_ ag2.body\[313\] vssd1 vssd1 vccd1 vccd1 _04104_ sky130_fd_sc_hd__inv_2
XFILLER_0_130_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12129__B1 net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1414_X net1414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11110_ net1085 control.body\[1102\] vssd1 vssd1 vccd1 vccd1 _06083_ sky130_fd_sc_hd__nand2b_1
X_20308_ clknet_leaf_70_clk net1572 net1497 vssd1 vssd1 vccd1 vccd1 obsmode.sOBSMODE.pb_2
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_13_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12090_ img_gen.tracker.frame\[291\] net612 net595 img_gen.tracker.frame\[297\] _07061_
+ vssd1 vssd1 vccd1 vccd1 _07062_ sky130_fd_sc_hd__a221o_1
XFILLER_0_130_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16689__X _02368_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout874_X net874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold770 control.body\[674\] vssd1 vssd1 vccd1 vccd1 net2332 sky130_fd_sc_hd__dlygate4sd3_1
Xhold781 control.body\[705\] vssd1 vssd1 vccd1 vccd1 net2343 sky130_fd_sc_hd__dlygate4sd3_1
Xhold792 control.body\[940\] vssd1 vssd1 vccd1 vccd1 net2354 sky130_fd_sc_hd__dlygate4sd3_1
X_11041_ net779 control.body\[1041\] _06012_ _06013_ net895 vssd1 vssd1 vccd1 vccd1
+ _06014_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_60_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20239_ clknet_leaf_69_clk _01183_ net1496 vssd1 vssd1 vccd1 vccd1 ag2.body\[157\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_9_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17952__C net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19102__CLK clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11058__B net1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_1349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14800_ net1020 ag2.body\[294\] vssd1 vssd1 vccd1 vccd1 _01471_ sky130_fd_sc_hd__or2_1
X_15780_ ag2.body\[307\] net208 _01638_ ag2.body\[299\] vssd1 vssd1 vccd1 vccd1 _01029_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__09751__B net1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12992_ net665 _07691_ vssd1 vssd1 vccd1 vccd1 _07692_ sky130_fd_sc_hd__nor2_1
XFILLER_0_98_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16006__A_N net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14731_ net993 ag2.body\[113\] vssd1 vssd1 vccd1 vccd1 _08892_ sky130_fd_sc_hd__nand2_1
XFILLER_0_73_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13273__B _07460_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11943_ img_gen.tracker.frame\[136\] net599 vssd1 vssd1 vccd1 vccd1 _06915_ sky130_fd_sc_hd__or2_1
XANTENNA__19252__CLK clknet_leaf_75_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16043__A1 net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17450_ _03125_ _03126_ _03127_ _03128_ vssd1 vssd1 vccd1 vccd1 _03129_ sky130_fd_sc_hd__or4_1
XANTENNA__17240__B1 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14662_ net1010 ag2.body\[527\] vssd1 vssd1 vccd1 vccd1 _08823_ sky130_fd_sc_hd__xor2_1
X_11874_ img_gen.tracker.frame\[250\] net581 net543 img_gen.tracker.frame\[247\] _06845_
+ vssd1 vssd1 vccd1 vccd1 _06846_ sky130_fd_sc_hd__o221a_1
XANTENNA__17791__A1 net1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17791__B2 net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16401_ obsg2.obstacleArray\[110\] obsg2.obstacleArray\[111\] net452 vssd1 vssd1
+ vccd1 vccd1 _02080_ sky130_fd_sc_hd__mux2_1
X_13613_ control.divider.count\[4\] _07958_ net220 vssd1 vssd1 vccd1 vccd1 _07984_
+ sky130_fd_sc_hd__o21ai_1
X_17381_ ag2.body\[492\] net962 vssd1 vssd1 vccd1 vccd1 _03060_ sky130_fd_sc_hd__nand2_1
XANTENNA__12604__A1 net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12065__C1 net468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10825_ _04433_ _04758_ net641 vssd1 vssd1 vccd1 vccd1 _05798_ sky130_fd_sc_hd__o21ai_4
X_14593_ net1033 ag2.body\[309\] vssd1 vssd1 vccd1 vccd1 _08754_ sky130_fd_sc_hd__xor2_1
XFILLER_0_95_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19120_ clknet_leaf_141_clk img_gen.tracker.next_frame\[558\] net1294 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[558\] sky130_fd_sc_hd__dfrtp_1
X_16332_ _02009_ _02010_ net418 vssd1 vssd1 vccd1 vccd1 _02011_ sky130_fd_sc_hd__mux2_1
XFILLER_0_113_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13544_ _06624_ _06632_ vssd1 vssd1 vccd1 vccd1 _07929_ sky130_fd_sc_hd__nand2_1
XANTENNA__11958__A3 _06929_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11812__C1 net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09481__B1 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10756_ net1131 control.body\[892\] vssd1 vssd1 vccd1 vccd1 _05729_ sky130_fd_sc_hd__or2_1
XFILLER_0_36_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14357__A1 net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19051_ clknet_leaf_10_clk img_gen.tracker.next_frame\[489\] net1273 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[489\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__14357__B2 net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16263_ obsg2.obstacleArray\[50\] obsg2.obstacleArray\[51\] net405 vssd1 vssd1 vccd1
+ vccd1 _01942_ sky130_fd_sc_hd__mux2_1
X_13475_ net308 _07595_ vssd1 vssd1 vccd1 vccd1 _07902_ sky130_fd_sc_hd__nor2_1
X_10687_ ag2.body\[146\] net1185 vssd1 vssd1 vccd1 vccd1 _05660_ sky130_fd_sc_hd__xor2_1
XFILLER_0_10_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18002_ _03540_ _03569_ vssd1 vssd1 vccd1 vccd1 _03616_ sky130_fd_sc_hd__nor2_1
XANTENNA__09766__X _04739_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15214_ control.body\[812\] net93 _01575_ net2504 vssd1 vssd1 vccd1 vccd1 _00526_
+ sky130_fd_sc_hd__a22o_1
X_12426_ _06505_ _06556_ _06558_ vssd1 vssd1 vccd1 vccd1 _07388_ sky130_fd_sc_hd__nand3b_1
X_16194_ obsg2.obstacleArray\[47\] net430 net376 _01872_ vssd1 vssd1 vccd1 vccd1 _01873_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_22_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_806 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15145_ net2529 net106 _01567_ control.body\[871\] vssd1 vssd1 vccd1 vccd1 _00465_
+ sky130_fd_sc_hd__a22o_1
X_12357_ _07291_ _07322_ _07323_ _07292_ vssd1 vssd1 vccd1 vccd1 _07324_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_121_841 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12633__A net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11308_ ag2.body\[276\] net1137 vssd1 vssd1 vccd1 vccd1 _06281_ sky130_fd_sc_hd__xor2_1
X_19953_ clknet_leaf_45_clk _00897_ net1382 vssd1 vssd1 vccd1 vccd1 ag2.body\[447\]
+ sky130_fd_sc_hd__dfrtp_4
X_15076_ net2661 net148 _01561_ net2473 vssd1 vssd1 vccd1 vccd1 _00402_ sky130_fd_sc_hd__a22o_1
X_12288_ img_gen.updater.commands.mode\[2\] img_gen.control.current\[1\] img_gen.control.current\[0\]
+ _04388_ vssd1 vssd1 vccd1 vccd1 _07258_ sky130_fd_sc_hd__or4_1
XANTENNA__17059__B1 net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09536__A1 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14027_ net798 ag2.body\[30\] ag2.body\[28\] net811 vssd1 vssd1 vccd1 vccd1 _08188_
+ sky130_fd_sc_hd__a2bb2o_1
X_18904_ clknet_leaf_144_clk img_gen.tracker.next_frame\[342\] net1251 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[342\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__09536__B2 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10153__A ag2.body\[59\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11239_ ag2.body\[193\] net1208 vssd1 vssd1 vccd1 vccd1 _06212_ sky130_fd_sc_hd__or2_1
XANTENNA__11879__C1 net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19884_ clknet_leaf_86_clk _00828_ net1462 vssd1 vssd1 vccd1 vccd1 ag2.body\[506\]
+ sky130_fd_sc_hd__dfrtp_4
X_18835_ clknet_leaf_4_clk img_gen.tracker.next_frame\[273\] net1260 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[273\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_69_2422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_2433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09661__B net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15978_ net1043 _08119_ vssd1 vssd1 vccd1 vccd1 _01663_ sky130_fd_sc_hd__and2_1
XFILLER_0_93_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18766_ clknet_leaf_16_clk img_gen.tracker.next_frame\[204\] net1315 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[204\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_2308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17717_ _03394_ _03395_ net378 vssd1 vssd1 vccd1 vccd1 _03396_ sky130_fd_sc_hd__mux2_1
XANTENNA__13183__B net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14929_ control.body\[1071\] net167 _01543_ net2338 vssd1 vssd1 vccd1 vccd1 _00273_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_65_2319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18697_ clknet_leaf_29_clk img_gen.tracker.next_frame\[135\] net1335 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[135\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_8_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17231__B1 net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10854__B1 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17648_ ag2.body\[36\] net959 vssd1 vssd1 vccd1 vccd1 _03327_ sky130_fd_sc_hd__xor2_1
XANTENNA__17782__A1 net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19745__CLK clknet_leaf_131_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12056__C1 net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17579_ ag2.body\[343\] net934 vssd1 vssd1 vccd1 vccd1 _03258_ sky130_fd_sc_hd__nand2_1
X_19318_ clknet_leaf_105_clk _00262_ net1433 vssd1 vssd1 vccd1 vccd1 control.body\[1076\]
+ sky130_fd_sc_hd__dfrtp_1
X_20590_ net1522 vssd1 vssd1 vccd1 vccd1 gpio_oeb[2] sky130_fd_sc_hd__buf_2
XFILLER_0_85_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_462 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19249_ clknet_leaf_75_clk _00193_ net1482 vssd1 vssd1 vccd1 vccd1 ag2.body\[112\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_27_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09002_ ag2.body\[119\] vssd1 vssd1 vccd1 vccd1 _04027_ sky130_fd_sc_hd__inv_2
XFILLER_0_42_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15838__B net59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18214__B net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_154 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout200_A net218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11582__A1 _06511_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19125__CLK clknet_leaf_141_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13859__B1 _08134_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout502 _01708_ vssd1 vssd1 vccd1 vccd1 net502 sky130_fd_sc_hd__clkbuf_4
X_09904_ ag2.body\[131\] net1165 vssd1 vssd1 vccd1 vccd1 _04877_ sky130_fd_sc_hd__xor2_1
XANTENNA__14520__A1 net1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout513 net515 vssd1 vssd1 vccd1 vccd1 net513 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_6_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout524 net528 vssd1 vssd1 vccd1 vccd1 net524 sky130_fd_sc_hd__buf_2
XANTENNA__14520__B2 net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1207_A net1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20024_ clknet_leaf_58_clk _00968_ net1471 vssd1 vssd1 vccd1 vccd1 ag2.body\[374\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__09852__A net1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout546 net547 vssd1 vssd1 vccd1 vccd1 net546 sky130_fd_sc_hd__clkbuf_4
XANTENNA_input5_A gpio_in[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09835_ net1157 control.body\[923\] vssd1 vssd1 vccd1 vccd1 _04808_ sky130_fd_sc_hd__nand2_1
Xfanout557 _06651_ vssd1 vssd1 vccd1 vccd1 net557 sky130_fd_sc_hd__buf_2
XANTENNA__18262__A2 _03533_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout568 net573 vssd1 vssd1 vccd1 vccd1 net568 sky130_fd_sc_hd__clkbuf_4
XANTENNA__16021__Y _01700_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout579 net582 vssd1 vssd1 vccd1 vccd1 net579 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout667_A net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout288_X net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10350__X _05323_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17470__B1 net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09766_ _04728_ _04733_ _04738_ _04539_ vssd1 vssd1 vccd1 vccd1 _04739_ sky130_fd_sc_hd__or4b_2
XANTENNA__13087__A1 net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14189__B ag2.body\[160\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout834_A net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09697_ ag2.body\[69\] net1114 vssd1 vssd1 vccd1 vccd1 _04670_ sky130_fd_sc_hd__nand2_1
XFILLER_0_90_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17222__B1 net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1197_X net1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14587__A1 net845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14587__B2 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout622_X net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10610_ net1181 control.body\[986\] vssd1 vssd1 vccd1 vccd1 _05583_ sky130_fd_sc_hd__xor2_1
X_11590_ obsg2.obstacleArray\[0\] obsg2.obstacleArray\[1\] obsg2.obstacleArray\[4\]
+ obsg2.obstacleArray\[5\] net1124 net513 vssd1 vssd1 vccd1 vccd1 _06563_ sky130_fd_sc_hd__mux4_1
XANTENNA__12062__A2 net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_94_3205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10541_ ag2.body\[231\] net1061 vssd1 vssd1 vccd1 vccd1 _05514_ sky130_fd_sc_hd__or2_1
XANTENNA__16624__S net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13260_ net236 _07817_ _07818_ net1834 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[399\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_126_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout991_X net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10472_ net1204 control.body\[1009\] vssd1 vssd1 vccd1 vccd1 _05445_ sky130_fd_sc_hd__xor2_1
XFILLER_0_32_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17289__B1 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12211_ _07182_ net465 img_gen.control.current\[1\] vssd1 vssd1 vccd1 vccd1 _07183_
+ sky130_fd_sc_hd__and3b_1
XFILLER_0_103_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13191_ net675 _07785_ vssd1 vssd1 vccd1 vccd1 _07786_ sky130_fd_sc_hd__nor2_1
XANTENNA__12453__A net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12142_ img_gen.tracker.frame\[522\] net544 _07113_ net571 vssd1 vssd1 vccd1 vccd1
+ _07114_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_88_3009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16950_ ag2.body\[387\] net718 net697 ag2.body\[390\] _02628_ vssd1 vssd1 vccd1 vccd1
+ _02629_ sky130_fd_sc_hd__a221o_1
X_12073_ img_gen.tracker.frame\[102\] net556 _07044_ net572 vssd1 vssd1 vccd1 vccd1
+ _07045_ sky130_fd_sc_hd__a211o_1
X_11024_ ag2.body\[595\] net1147 vssd1 vssd1 vccd1 vccd1 _05997_ sky130_fd_sc_hd__or2_1
X_15901_ _05543_ net55 vssd1 vssd1 vccd1 vccd1 _01651_ sky130_fd_sc_hd__nor2_2
X_16881_ ag2.body\[19\] net848 vssd1 vssd1 vccd1 vccd1 _02560_ sky130_fd_sc_hd__xor2_1
XANTENNA__11876__A2 net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13284__A net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15832_ ag2.body\[258\] net201 net49 ag2.body\[250\] vssd1 vssd1 vccd1 vccd1 _01076_
+ sky130_fd_sc_hd__a22o_1
X_18620_ clknet_leaf_145_clk img_gen.tracker.next_frame\[58\] net1241 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[58\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__18642__CLK clknet_leaf_131_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19768__CLK clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15763_ ag2.body\[324\] net215 _01636_ ag2.body\[316\] vssd1 vssd1 vccd1 vccd1 _01014_
+ sky130_fd_sc_hd__a22o_1
X_18551_ clknet_leaf_132_clk _00077_ net1297 vssd1 vssd1 vccd1 vccd1 ag2.y\[3\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__12825__A1 net240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12975_ net341 _07502_ vssd1 vssd1 vccd1 vccd1 _07684_ sky130_fd_sc_hd__or2_1
XFILLER_0_63_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14714_ net1003 _04118_ ag2.body\[342\] net803 vssd1 vssd1 vccd1 vccd1 _08875_ sky130_fd_sc_hd__a22o_1
XANTENNA__17043__X _02722_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17502_ _03176_ _03177_ _03180_ vssd1 vssd1 vccd1 vccd1 _03181_ sky130_fd_sc_hd__a21o_1
XFILLER_0_87_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18482_ net1515 net1509 vssd1 vssd1 vccd1 vccd1 _00013_ sky130_fd_sc_hd__or2_1
X_11926_ img_gen.tracker.frame\[289\] img_gen.tracker.frame\[292\] img_gen.tracker.frame\[295\]
+ img_gen.tracker.frame\[298\] net1216 net1191 vssd1 vssd1 vccd1 vccd1 _06898_ sky130_fd_sc_hd__mux4_1
X_15694_ _04430_ net64 vssd1 vssd1 vccd1 vccd1 _01628_ sky130_fd_sc_hd__and2_2
XTAP_TAPCELL_ROW_16_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16567__A2 net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17433_ ag2.body\[144\] net741 net855 _04041_ _03111_ vssd1 vssd1 vccd1 vccd1 _03112_
+ sky130_fd_sc_hd__a221o_1
X_14645_ net820 ag2.body\[515\] ag2.body\[519\] net794 vssd1 vssd1 vccd1 vccd1 _08806_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_131_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14578__B2 net1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11857_ img_gen.tracker.frame\[232\] net608 net591 img_gen.tracker.frame\[238\] vssd1
+ vssd1 vccd1 vccd1 _06829_ sky130_fd_sc_hd__o22a_1
XFILLER_0_83_820 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12589__B1 net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11532__A net1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17364_ _03035_ _03036_ _03040_ _03016_ _03038_ vssd1 vssd1 vccd1 vccd1 _03043_ sky130_fd_sc_hd__a221o_1
X_10808_ _05670_ _05775_ _05780_ _05765_ vssd1 vssd1 vccd1 vccd1 _05781_ sky130_fd_sc_hd__o31a_2
XFILLER_0_126_911 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14576_ net1032 ag2.body\[493\] vssd1 vssd1 vccd1 vccd1 _08737_ sky130_fd_sc_hd__xor2_1
XANTENNA__10385__C_N _05347_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11788_ img_gen.tracker.frame\[350\] net615 net542 img_gen.tracker.frame\[356\] _06759_
+ vssd1 vssd1 vccd1 vccd1 _06760_ sky130_fd_sc_hd__o221a_1
XFILLER_0_125_410 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16315_ net415 _01991_ _01993_ net371 vssd1 vssd1 vccd1 vccd1 _01994_ sky130_fd_sc_hd__a211o_1
X_19103_ clknet_leaf_0_clk img_gen.tracker.next_frame\[541\] net1240 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[541\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13527_ img_gen.tracker.frame\[563\] net657 _07921_ vssd1 vssd1 vccd1 vccd1 _07922_
+ sky130_fd_sc_hd__and3_1
X_17295_ ag2.body\[348\] net966 vssd1 vssd1 vccd1 vccd1 _02974_ sky130_fd_sc_hd__or2_1
X_10739_ ag2.body\[503\] net1064 vssd1 vssd1 vccd1 vccd1 _05712_ sky130_fd_sc_hd__xor2_1
XANTENNA__10148__A ag2.body\[58\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19148__CLK clknet_leaf_51_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_2101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09496__X _04469_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19034_ clknet_leaf_6_clk img_gen.tracker.next_frame\[472\] net1264 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[472\] sky130_fd_sc_hd__dfrtp_1
X_16246_ _01923_ _01924_ net415 vssd1 vssd1 vccd1 vccd1 _01925_ sky130_fd_sc_hd__mux2_1
X_13458_ net256 _07894_ _07895_ net1592 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[520\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_70_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12409_ net748 _06630_ vssd1 vssd1 vccd1 vccd1 _07372_ sky130_fd_sc_hd__or2_1
XFILLER_0_45_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16177_ obsg2.obstacleArray\[55\] net430 net376 _01855_ vssd1 vssd1 vccd1 vccd1 _01856_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_49_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13389_ net229 _07868_ _07869_ net1988 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[477\]
+ sky130_fd_sc_hd__a22o_1
X_15128_ _05634_ net58 vssd1 vssd1 vccd1 vccd1 _01566_ sky130_fd_sc_hd__nor2_2
XFILLER_0_121_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12513__D net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19936_ clknet_leaf_47_clk _00880_ net1375 vssd1 vssd1 vccd1 vccd1 ag2.body\[462\]
+ sky130_fd_sc_hd__dfrtp_4
X_15059_ control.body\[945\] net149 _01559_ net2245 vssd1 vssd1 vccd1 vccd1 _00387_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__18050__A net43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire635_A _04633_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18244__A2 net37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19867_ clknet_leaf_95_clk _00811_ net1440 vssd1 vssd1 vccd1 vccd1 ag2.body\[521\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_128_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_1471 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17452__B1 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09620_ net783 control.body\[800\] control.body\[801\] net777 _04588_ vssd1 vssd1
+ vccd1 vccd1 _04593_ sky130_fd_sc_hd__a221o_1
X_18818_ clknet_leaf_5_clk img_gen.tracker.next_frame\[256\] net1249 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[256\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__10611__A net1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13069__A1 net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19798_ clknet_leaf_127_clk _00742_ net1330 vssd1 vssd1 vccd1 vccd1 ag2.body\[596\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__14805__A2 ag2.body\[288\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09551_ net1170 control.body\[722\] vssd1 vssd1 vccd1 vccd1 _04524_ sky130_fd_sc_hd__xor2_1
XFILLER_0_91_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18749_ clknet_leaf_143_clk img_gen.tracker.next_frame\[187\] net1257 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[187\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__12816__A1 net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_1506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09482_ ag2.body\[465\] net782 net1055 _04167_ vssd1 vssd1 vccd1 vccd1 _04455_ sky130_fd_sc_hd__a22o_1
XFILLER_0_17_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14569__A1 net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14569__B2 net1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_872 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout150_A net154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11442__A net1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1241 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12044__A2 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13241__A1 net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_533 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19593__RESET_B net1386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11161__B net1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20573_ clknet_leaf_106_clk _01431_ _00037_ vssd1 vssd1 vccd1 vccd1 sound_gen.dac1.dacCount\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_34_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16444__S net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout415_A net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1157_A net1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09847__A net1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17256__A2_N net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14741__A1 net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14741__B2 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1324_A net1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_468 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13088__B _07567_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17783__B net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout784_A net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20080__RESET_B net1492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1308 net1309 vssd1 vssd1 vccd1 vccd1 net1308 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout1112_X net1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout310 net311 vssd1 vssd1 vccd1 vccd1 net310 sky130_fd_sc_hd__buf_2
XFILLER_0_121_1257 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout321 track.nextHighScore\[5\] vssd1 vssd1 vccd1 vccd1 net321 sky130_fd_sc_hd__buf_2
Xfanout1319 net1320 vssd1 vssd1 vccd1 vccd1 net1319 sky130_fd_sc_hd__clkbuf_4
Xfanout332 net333 vssd1 vssd1 vccd1 vccd1 net332 sky130_fd_sc_hd__buf_2
Xfanout343 net344 vssd1 vssd1 vccd1 vccd1 net343 sky130_fd_sc_hd__clkbuf_4
Xfanout354 _01702_ vssd1 vssd1 vccd1 vccd1 net354 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout951_A net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11858__A2 net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout365 _02068_ vssd1 vssd1 vccd1 vccd1 net365 sky130_fd_sc_hd__clkbuf_4
X_20007_ clknet_leaf_59_clk _00951_ net1467 vssd1 vssd1 vccd1 vccd1 ag2.body\[389\]
+ sky130_fd_sc_hd__dfrtp_4
Xfanout376 net379 vssd1 vssd1 vccd1 vccd1 net376 sky130_fd_sc_hd__buf_4
XANTENNA__17443__B1 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout387 net388 vssd1 vssd1 vccd1 vccd1 net387 sky130_fd_sc_hd__buf_2
X_09818_ net917 net922 net913 net909 vssd1 vssd1 vccd1 vccd1 _04791_ sky130_fd_sc_hd__a211o_4
Xfanout398 net400 vssd1 vssd1 vccd1 vccd1 net398 sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_fanout63_A _08131_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09749_ _04716_ _04717_ _04720_ _04721_ vssd1 vssd1 vccd1 vccd1 _04722_ sky130_fd_sc_hd__or4b_1
XANTENNA__10240__B net1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout837_X net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12760_ net284 _07582_ _07583_ net1900 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[134\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_97_967 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11711_ img_gen.tracker.frame\[323\] net585 net546 img_gen.tracker.frame\[320\] _06682_
+ vssd1 vssd1 vccd1 vccd1 _06683_ sky130_fd_sc_hd__o221a_1
XFILLER_0_96_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12691_ net285 _07549_ _07550_ net1971 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[98\]
+ sky130_fd_sc_hd__a22o_1
X_14430_ net832 ag2.body\[553\] ag2.body\[555\] net817 _08590_ vssd1 vssd1 vccd1 vccd1
+ _08591_ sky130_fd_sc_hd__a221o_1
X_11642_ net505 _06613_ _06614_ net759 vssd1 vssd1 vccd1 vccd1 _06615_ sky130_fd_sc_hd__a211o_1
XFILLER_0_83_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13232__A1 net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12035__A2 net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10239__Y _05212_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16862__B net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11071__B net1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14361_ net1015 ag2.body\[606\] vssd1 vssd1 vccd1 vccd1 _08522_ sky130_fd_sc_hd__xnor2_1
X_11573_ obsg2.obstacleArray\[86\] net631 vssd1 vssd1 vccd1 vccd1 _06546_ sky130_fd_sc_hd__or2_1
XANTENNA__19263__RESET_B net1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16354__S net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10896__D_N _05857_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20148__CLK clknet_leaf_98_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14663__A net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16100_ obsg2.obstacleArray\[80\] obsg2.obstacleArray\[81\] net428 vssd1 vssd1 vccd1
+ vccd1 _01779_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13312_ net1935 net647 _07837_ _07838_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[431\]
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_134_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17080_ ag2.body\[196\] net962 vssd1 vssd1 vccd1 vccd1 _02759_ sky130_fd_sc_hd__or2_1
X_10524_ net1180 control.body\[914\] vssd1 vssd1 vccd1 vccd1 _05497_ sky130_fd_sc_hd__xor2_1
X_14292_ net1015 ag2.body\[478\] vssd1 vssd1 vccd1 vccd1 _08453_ sky130_fd_sc_hd__xor2_1
XFILLER_0_80_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16721__A2 net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11498__S net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16031_ _01678_ _01682_ vssd1 vssd1 vccd1 vccd1 _01710_ sky130_fd_sc_hd__xnor2_1
XANTENNA__20168__RESET_B net1480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13243_ net238 net314 _07435_ _07810_ net2077 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[390\]
+ sky130_fd_sc_hd__a32o_1
XANTENNA__13279__A net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10455_ ag2.body\[450\] net1176 vssd1 vssd1 vccd1 vccd1 _05428_ sky130_fd_sc_hd__nand2_1
XFILLER_0_106_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09476__B net1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12183__A net1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11546__A1 net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12614__C net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13174_ net341 _07607_ vssd1 vssd1 vccd1 vccd1 _07778_ sky130_fd_sc_hd__nor2_1
X_10386_ _04604_ _05340_ _05345_ _05358_ vssd1 vssd1 vccd1 vccd1 _05359_ sky130_fd_sc_hd__o31a_1
XFILLER_0_62_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_1591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10415__B _05335_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16485__A1 net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_43_clk_X clknet_leaf_43_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12125_ img_gen.tracker.frame\[537\] net579 net541 img_gen.tracker.frame\[534\] vssd1
+ vssd1 vccd1 vccd1 _07097_ sky130_fd_sc_hd__o22a_1
XANTENNA__12470__X _07425_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17982_ net351 _03539_ net39 vssd1 vssd1 vccd1 vccd1 _03602_ sky130_fd_sc_hd__and3_1
XANTENNA__12415__A_N net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19590__CLK clknet_leaf_118_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19721_ clknet_leaf_132_clk _00665_ net1303 vssd1 vssd1 vccd1 vccd1 control.body\[679\]
+ sky130_fd_sc_hd__dfrtp_1
X_12056_ img_gen.tracker.frame\[78\] net555 _07027_ net575 vssd1 vssd1 vccd1 vccd1
+ _07028_ sky130_fd_sc_hd__a211oi_1
X_16933_ ag2.body\[521\] net873 vssd1 vssd1 vccd1 vccd1 _02612_ sky130_fd_sc_hd__or2_1
XANTENNA__12630__B net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16102__B net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16237__A1 net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11007_ _04425_ net635 vssd1 vssd1 vccd1 vccd1 _05980_ sky130_fd_sc_hd__nand2_1
X_19652_ clknet_leaf_133_clk net2483 net1308 vssd1 vssd1 vccd1 vccd1 control.body\[738\]
+ sky130_fd_sc_hd__dfrtp_1
X_16864_ ag2.body\[200\] net739 net952 _04065_ vssd1 vssd1 vccd1 vccd1 _02543_ sky130_fd_sc_hd__a22o_1
X_18603_ clknet_leaf_16_clk img_gen.tracker.next_frame\[41\] net1320 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[41\] sky130_fd_sc_hd__dfrtp_1
X_15815_ ag2.body\[274\] net205 _01642_ ag2.body\[266\] vssd1 vssd1 vccd1 vccd1 _01060_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11246__B net1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16795_ _02075_ _02473_ _02472_ vssd1 vssd1 vccd1 vccd1 _02474_ sky130_fd_sc_hd__a21oi_1
X_19583_ clknet_leaf_117_clk _00527_ net1385 vssd1 vssd1 vccd1 vccd1 control.body\[813\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10150__B net1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15746_ ag2.body\[341\] net211 _01634_ ag2.body\[333\] vssd1 vssd1 vccd1 vccd1 _00999_
+ sky130_fd_sc_hd__a22o_1
X_18534_ clknet_leaf_136_clk _00060_ net1300 vssd1 vssd1 vccd1 vccd1 img_gen.updater.commands.count\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_90_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_967 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12958_ _07490_ _07639_ vssd1 vssd1 vccd1 vccd1 _07676_ sky130_fd_sc_hd__nor2_1
XANTENNA__14557__B ag2.body\[65\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1602 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11909_ img_gen.tracker.frame\[376\] net608 net549 img_gen.tracker.frame\[379\] _06880_
+ vssd1 vssd1 vccd1 vccd1 _06881_ sky130_fd_sc_hd__o221a_1
X_18465_ _04261_ net737 _03952_ vssd1 vssd1 vccd1 vccd1 _01423_ sky130_fd_sc_hd__a21oi_1
X_15677_ _06399_ net58 vssd1 vssd1 vccd1 vccd1 _01627_ sky130_fd_sc_hd__nor2_4
XANTENNA__19202__Q ag2.body\[65\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12889_ net267 _07643_ _07644_ net1963 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[202\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_8_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14628_ net842 ag2.body\[464\] ag2.body\[466\] net825 _08788_ vssd1 vssd1 vccd1 vccd1
+ _08789_ sky130_fd_sc_hd__a221o_1
X_17416_ ag2.body\[280\] net740 net719 ag2.body\[283\] vssd1 vssd1 vccd1 vccd1 _03095_
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_114_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_1512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18396_ _03791_ _03883_ _03884_ _03885_ _03789_ vssd1 vssd1 vccd1 vccd1 _03886_ sky130_fd_sc_hd__o311a_1
XANTENNA__13223__A1 net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12026__A2 net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17347_ net926 ag2.body\[6\] vssd1 vssd1 vccd1 vccd1 _03026_ sky130_fd_sc_hd__nand2_1
XFILLER_0_7_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10037__B2 _04944_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14559_ net986 _04000_ _04001_ net1023 vssd1 vssd1 vccd1 vccd1 _08720_ sky130_fd_sc_hd__a22o_1
XANTENNA__15021__X _01555_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17278_ net723 ag2.body\[554\] _04203_ net869 vssd1 vssd1 vccd1 vccd1 _02957_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_71_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14292__B ag2.body\[478\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16229_ _01905_ _01906_ vssd1 vssd1 vccd1 vccd1 _01908_ sky130_fd_sc_hd__or2_1
XFILLER_0_12_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19017_ clknet_leaf_1_clk img_gen.tracker.next_frame\[455\] net1246 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[455\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14860__X _01531_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10606__A net1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_1490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18465__A2 net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10325__B net1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17673__B1 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08982_ ag2.body\[76\] vssd1 vssd1 vccd1 vccd1 _04007_ sky130_fd_sc_hd__inv_2
XFILLER_0_80_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19919_ clknet_leaf_52_clk _00863_ net1456 vssd1 vssd1 vccd1 vccd1 ag2.body\[477\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__16012__B net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09603_ net1047 control.body\[639\] vssd1 vssd1 vccd1 vccd1 _04576_ sky130_fd_sc_hd__xor2_1
XANTENNA__11156__B net1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout365_A _02068_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14748__A net1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09534_ net787 control.body\[1024\] control.body\[1028\] net761 vssd1 vssd1 vccd1
+ vccd1 _04507_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_91_1352 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13462__A1 net235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10995__B net1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09465_ _04133_ net1234 net1139 _04136_ _04437_ vssd1 vssd1 vccd1 vccd1 _04438_ sky130_fd_sc_hd__a221o_1
XFILLER_0_91_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout532_A net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11172__A net1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12017__A2 net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09396_ sound_gen.osc1.stayCount\[5\] _04344_ net271 vssd1 vssd1 vccd1 vccd1 _04382_
+ sky130_fd_sc_hd__o21ai_1
XANTENNA__14411__B1 net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15579__A _04429_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20625_ sound_gen.dac1.dacCount\[3\] vssd1 vssd1 vccd1 vccd1 net12 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_47_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout418_X net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1062_X net1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1441_A net1442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09577__A net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_785 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20556_ clknet_leaf_105_clk _01421_ _00030_ vssd1 vssd1 vccd1 vccd1 sound_gen.osc1.stayCount\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__16703__A2 net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12715__B _07561_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout999_A net1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13099__A net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14714__A1 net1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14714__B2 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15911__B1 _01652_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20487_ clknet_leaf_37_clk _01374_ net1351 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[123\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__11528__A1 net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10240_ ag2.body\[320\] net1236 vssd1 vssd1 vccd1 vccd1 _05213_ sky130_fd_sc_hd__nand2_1
XANTENNA__18456__A2 _04791_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10235__B net1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout787_X net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14930__B net59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16467__A1 net403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17944__D net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17664__B1 net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10171_ _05133_ _05142_ _05143_ vssd1 vssd1 vccd1 vccd1 _05144_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_110_3680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_3691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_110_Right_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1105 net1106 vssd1 vssd1 vccd1 vccd1 net1105 sky130_fd_sc_hd__buf_2
XANTENNA__10751__A2 _05703_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1116 net1117 vssd1 vssd1 vccd1 vccd1 net1116 sky130_fd_sc_hd__buf_4
XFILLER_0_121_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1127 net1129 vssd1 vssd1 vccd1 vccd1 net1127 sky130_fd_sc_hd__buf_4
XANTENNA__18208__A2 _03566_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout954_X net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout140 net141 vssd1 vssd1 vccd1 vccd1 net140 sky130_fd_sc_hd__buf_2
Xfanout1138 net1139 vssd1 vssd1 vccd1 vccd1 net1138 sky130_fd_sc_hd__buf_4
XFILLER_0_22_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1149 net1151 vssd1 vssd1 vccd1 vccd1 net1149 sky130_fd_sc_hd__buf_2
Xfanout151 net154 vssd1 vssd1 vccd1 vccd1 net151 sky130_fd_sc_hd__buf_2
XANTENNA__17416__B1 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout162 net183 vssd1 vssd1 vccd1 vccd1 net162 sky130_fd_sc_hd__clkbuf_2
X_13930_ ag2.body\[73\] net186 _08153_ ag2.body\[65\] vssd1 vssd1 vccd1 vccd1 _00154_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__10251__A net1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout173 net174 vssd1 vssd1 vccd1 vccd1 net173 sky130_fd_sc_hd__buf_2
XANTENNA__17960__C net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout184 net187 vssd1 vssd1 vccd1 vccd1 net184 sky130_fd_sc_hd__buf_2
Xfanout195 net196 vssd1 vssd1 vccd1 vccd1 net195 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout66_X net66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16857__B net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13861_ net325 net323 vssd1 vssd1 vccd1 vccd1 _08135_ sky130_fd_sc_hd__nor2_1
XFILLER_0_134_1404 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15600_ ag2.body\[466\] net121 _01619_ ag2.body\[458\] vssd1 vssd1 vccd1 vccd1 _00868_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_92_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12812_ net307 _07607_ vssd1 vssd1 vccd1 vccd1 _07608_ sky130_fd_sc_hd__nor2_1
XANTENNA__15442__A2 net90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16580_ obsg2.obstacleArray\[112\] obsg2.obstacleArray\[113\] net443 vssd1 vssd1
+ vccd1 vccd1 _02259_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_2_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13453__A1 net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13792_ img_gen.updater.commands.count\[14\] img_gen.updater.commands.count\[13\]
+ _08091_ vssd1 vssd1 vccd1 vccd1 _08099_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_2_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_3484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_3495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_1414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_70_clk_A clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15531_ ag2.body\[534\] net157 _01610_ ag2.body\[526\] vssd1 vssd1 vccd1 vccd1 _00808_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11464__B1 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12743_ net334 _07467_ vssd1 vssd1 vccd1 vccd1 _07575_ sky130_fd_sc_hd__or2_1
XFILLER_0_70_1436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_3359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12178__A net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18250_ _03691_ net35 vssd1 vssd1 vccd1 vccd1 _03764_ sky130_fd_sc_hd__nor2_1
X_15462_ ag2.body\[584\] net90 _01603_ ag2.body\[576\] vssd1 vssd1 vccd1 vccd1 _00746_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__17688__B net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12008__A2 net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12674_ net435 net467 _06671_ _07452_ vssd1 vssd1 vccd1 vccd1 _07542_ sky130_fd_sc_hd__or4_4
XFILLER_0_60_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17201_ _04054_ net884 net949 _04057_ _02875_ vssd1 vssd1 vccd1 vccd1 _02880_ sky130_fd_sc_hd__a221o_1
X_14413_ _08563_ _08567_ _08569_ _08573_ vssd1 vssd1 vccd1 vccd1 _08574_ sky130_fd_sc_hd__or4_2
XANTENNA__20349__RESET_B net1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18181_ net519 _03729_ vssd1 vssd1 vccd1 vccd1 _01338_ sky130_fd_sc_hd__nor2_1
X_11625_ obsg2.obstacleArray\[42\] net633 net509 obsg2.obstacleArray\[46\] net759
+ vssd1 vssd1 vccd1 vccd1 _06598_ sky130_fd_sc_hd__o221a_1
XFILLER_0_25_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15393_ net2226 net80 _01596_ net2526 vssd1 vssd1 vccd1 vccd1 _00684_ sky130_fd_sc_hd__a22o_1
XANTENNA__14393__A net1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_85_clk_A clknet_4_12__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17132_ ag2.body\[518\] net942 vssd1 vssd1 vccd1 vccd1 _02811_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_117_3878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_1481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16155__A0 obsg2.obstacleArray\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14344_ net1026 ag2.body\[613\] vssd1 vssd1 vccd1 vccd1 _08505_ sky130_fd_sc_hd__xor2_1
X_11556_ _06528_ vssd1 vssd1 vccd1 vccd1 _06529_ sky130_fd_sc_hd__inv_2
XANTENNA__18830__CLK clknet_leaf_141_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_3889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17063_ _02736_ _02738_ _02741_ vssd1 vssd1 vccd1 vccd1 _02742_ sky130_fd_sc_hd__or3_2
X_10507_ net1133 control.body\[980\] vssd1 vssd1 vccd1 vccd1 _05480_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_69_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14275_ _08428_ _08429_ _08432_ _08433_ vssd1 vssd1 vccd1 vccd1 _08436_ sky130_fd_sc_hd__a22o_1
XFILLER_0_123_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11487_ net1197 net1078 vssd1 vssd1 vccd1 vccd1 _06460_ sky130_fd_sc_hd__and2_1
XFILLER_0_46_1630 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16014_ net732 net860 net882 vssd1 vssd1 vccd1 vccd1 _01693_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_21_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13226_ net675 _07802_ vssd1 vssd1 vccd1 vccd1 _07803_ sky130_fd_sc_hd__nor2_1
XFILLER_0_110_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10438_ _05407_ _05408_ _05409_ _05410_ _05406_ vssd1 vssd1 vccd1 vccd1 _05411_ sky130_fd_sc_hd__o221a_1
XFILLER_0_104_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_438 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16458__A1 net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18980__CLK clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09934__B net1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13157_ _07501_ net327 net336 vssd1 vssd1 vccd1 vccd1 _07770_ sky130_fd_sc_hd__and3b_1
XFILLER_0_85_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12641__A net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10369_ net767 control.body\[763\] control.body\[764\] net762 _05341_ vssd1 vssd1
+ vccd1 vccd1 _05342_ sky130_fd_sc_hd__o221ai_1
XFILLER_0_42_1549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_143_clk_A clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12108_ img_gen.tracker.frame\[171\] net610 net555 img_gen.tracker.frame\[174\] _07079_
+ vssd1 vssd1 vccd1 vccd1 _07080_ sky130_fd_sc_hd__a221o_1
X_17965_ net380 _01713_ net490 vssd1 vssd1 vccd1 vccd1 _03589_ sky130_fd_sc_hd__and3_1
X_13088_ net343 _07567_ vssd1 vssd1 vccd1 vccd1 _07737_ sky130_fd_sc_hd__nor2_1
XANTENNA_clkbuf_leaf_23_clk_A clknet_4_6__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19704_ clknet_leaf_135_clk net2273 net1301 vssd1 vssd1 vccd1 vccd1 control.body\[694\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11257__A net1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17407__B1 net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12039_ img_gen.tracker.frame\[12\] net629 net556 img_gen.tracker.frame\[18\] vssd1
+ vssd1 vccd1 vccd1 _07011_ sky130_fd_sc_hd__a22o_1
X_16916_ _02593_ _02594_ _02591_ _02592_ vssd1 vssd1 vccd1 vccd1 _02595_ sky130_fd_sc_hd__a211o_1
XANTENNA__17958__A1 net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17896_ net2174 _03531_ _03532_ _03519_ vssd1 vssd1 vccd1 vccd1 _01250_ sky130_fd_sc_hd__a22o_1
X_19635_ clknet_leaf_123_clk _00579_ net1406 vssd1 vssd1 vccd1 vccd1 control.body\[753\]
+ sky130_fd_sc_hd__dfrtp_1
X_16847_ ag2.body\[172\] net961 vssd1 vssd1 vccd1 vccd1 _02526_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_0_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19566_ clknet_leaf_115_clk net2462 net1388 vssd1 vssd1 vccd1 vccd1 control.body\[828\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13444__A1 net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_38_clk_A clknet_4_5__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16778_ obsg2.obstacleArray\[27\] net503 net488 obsg2.obstacleArray\[26\] _02456_
+ vssd1 vssd1 vccd1 vccd1 _02457_ sky130_fd_sc_hd__a221o_1
XANTENNA__10258__A1 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1634 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18517_ net1512 net1506 vssd1 vssd1 vccd1 vccd1 _00048_ sky130_fd_sc_hd__or2_1
X_15729_ ag2.body\[358\] net200 _01632_ ag2.body\[350\] vssd1 vssd1 vccd1 vccd1 _00984_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__14855__X _01526_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19497_ clknet_leaf_113_clk _00441_ net1399 vssd1 vssd1 vccd1 vccd1 control.body\[903\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_1678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09250_ img_gen.updater.commands.count\[16\] vssd1 vssd1 vccd1 vccd1 _04275_ sky130_fd_sc_hd__inv_2
X_18448_ _03835_ _03935_ _03936_ vssd1 vssd1 vccd1 vccd1 _03937_ sky130_fd_sc_hd__and3_1
XFILLER_0_34_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17598__B net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09181_ ag2.body\[561\] vssd1 vssd1 vccd1 vccd1 _04206_ sky130_fd_sc_hd__inv_2
XFILLER_0_8_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18379_ net323 _03801_ track.nextHighScore\[1\] vssd1 vssd1 vccd1 vccd1 _03869_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_29_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20410_ clknet_leaf_30_clk _01297_ net1357 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[46\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_16_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_133_4370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16146__B1 net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_133_4381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_133_4392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20341_ clknet_leaf_140_clk _01232_ net1297 vssd1 vssd1 vccd1 vccd1 img_gen.updater.commands.rR1.rainbowRNG\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_47_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout113_A net114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20272_ clknet_leaf_42_clk net1585 net1373 vssd1 vssd1 vccd1 vccd1 control.button4.Q\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10055__B net1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18222__B net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1022_A net1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08965_ ag2.body\[47\] vssd1 vssd1 vccd1 vccd1 _03990_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout482_A net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_1992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_4185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16958__A ag2.body\[291\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11167__A net1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_4196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10071__A net1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09887__B1 net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_1889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18071__B1 net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11694__B1 net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16169__S net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14478__A net1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19829__CLK clknet_leaf_124_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout747_A _04234_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13382__A _07542_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16621__B2 net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1489_A net1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09517_ net1076 control.body\[838\] vssd1 vssd1 vccd1 vccd1 _04490_ sky130_fd_sc_hd__xor2_1
XFILLER_0_56_1280 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13986__A2 net214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16693__A net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_734 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18374__A1 _07181_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout914_A net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09807__D_N _04772_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09859__X _04832_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09448_ net910 net914 vssd1 vssd1 vccd1 vccd1 _04421_ sky130_fd_sc_hd__and2_4
XFILLER_0_52_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20442__RESET_B net1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09578__Y _04551_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout702_X net702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09379_ sound_gen.osc1.stayCount\[14\] _04365_ net271 vssd1 vssd1 vccd1 vccd1 _04374_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_81_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11410_ _06374_ _06377_ _06379_ _06380_ vssd1 vssd1 vccd1 vccd1 _06383_ sky130_fd_sc_hd__or4_1
X_20608_ net1540 vssd1 vssd1 vccd1 vccd1 gpio_oeb[20] sky130_fd_sc_hd__buf_2
XFILLER_0_90_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12390_ _07292_ _07296_ vssd1 vssd1 vccd1 vccd1 _07355_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_10_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16688__A1 net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11341_ net891 _04239_ _04423_ _04428_ _04686_ vssd1 vssd1 vccd1 vccd1 _06314_ sky130_fd_sc_hd__o41a_4
XFILLER_0_132_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20539_ clknet_leaf_106_clk _01404_ _00013_ vssd1 vssd1 vccd1 vccd1 sound_gen.osc1.stayCount\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_34_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_112_3731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_3742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17955__C net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_112_3753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_788 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1263 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14060_ net824 ag2.body\[34\] _03986_ net1006 vssd1 vssd1 vccd1 vccd1 _08221_ sky130_fd_sc_hd__o22a_1
X_11272_ ag2.body\[126\] net1090 vssd1 vssd1 vccd1 vccd1 _06245_ sky130_fd_sc_hd__nand2_1
XFILLER_0_123_1127 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12174__A1 net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13011_ img_gen.tracker.frame\[268\] net654 vssd1 vssd1 vccd1 vccd1 _07701_ sky130_fd_sc_hd__and2_1
X_10223_ ag2.body\[567\] net1052 vssd1 vssd1 vccd1 vccd1 _05196_ sky130_fd_sc_hd__or2_1
XANTENNA__09754__B net1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17971__B _01713_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10154_ ag2.body\[59\] net1155 vssd1 vssd1 vccd1 vccd1 _05127_ sky130_fd_sc_hd__or2_1
X_17750_ _03156_ net389 _02501_ vssd1 vssd1 vccd1 vccd1 _03429_ sky130_fd_sc_hd__a21oi_2
X_14962_ net2617 net172 _01547_ control.body\[1028\] vssd1 vssd1 vccd1 vccd1 _00302_
+ sky130_fd_sc_hd__a22o_1
Xhold7 control.divider.synch.Q\[0\] vssd1 vssd1 vccd1 vccd1 net1569 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__20336__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10085_ net1075 control.body\[798\] vssd1 vssd1 vccd1 vccd1 _05058_ sky130_fd_sc_hd__nand2_1
XFILLER_0_57_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16701_ obsg2.obstacleArray\[82\] net489 net485 obsg2.obstacleArray\[81\] _02379_
+ vssd1 vssd1 vccd1 vccd1 _02380_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_106_3546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_106_3557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13913_ ag2.body\[58\] net129 _08151_ ag2.body\[50\] vssd1 vssd1 vccd1 vccd1 _00139_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_106_3568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16079__S net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17681_ _03356_ _03357_ _03358_ _03359_ vssd1 vssd1 vccd1 vccd1 _03360_ sky130_fd_sc_hd__or4_1
X_14893_ control.body\[1103\] net179 _01539_ net2199 vssd1 vssd1 vccd1 vccd1 _00241_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_57_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19420_ clknet_leaf_111_clk net2219 net1434 vssd1 vssd1 vccd1 vccd1 control.body\[970\]
+ sky130_fd_sc_hd__dfrtp_1
X_16632_ obsg2.obstacleArray\[60\] obsg2.obstacleArray\[61\] net444 vssd1 vssd1 vccd1
+ vccd1 _02311_ sky130_fd_sc_hd__mux2_1
X_13844_ ag2.body\[8\] net127 _08133_ net1044 vssd1 vssd1 vccd1 vccd1 _00088_ sky130_fd_sc_hd__a22o_1
XFILLER_0_76_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_1077 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__20486__CLK clknet_leaf_37_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19351_ clknet_leaf_101_clk net2438 net1439 vssd1 vssd1 vccd1 vccd1 control.body\[1045\]
+ sky130_fd_sc_hd__dfrtp_1
X_16563_ net350 _02206_ vssd1 vssd1 vccd1 vccd1 _02242_ sky130_fd_sc_hd__or2_1
X_13775_ _08086_ vssd1 vssd1 vccd1 vccd1 _08087_ sky130_fd_sc_hd__inv_2
XFILLER_0_71_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10987_ _05950_ _05951_ _05953_ _05954_ _05959_ vssd1 vssd1 vccd1 vccd1 _05960_ sky130_fd_sc_hd__a221o_1
XANTENNA__17168__A2 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18302_ track.nextHighScore\[1\] net326 vssd1 vssd1 vccd1 vccd1 _03798_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_80_2753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15514_ ag2.body\[551\] net155 _01608_ ag2.body\[543\] vssd1 vssd1 vccd1 vccd1 _00793_
+ sky130_fd_sc_hd__a22o_1
X_12726_ _07313_ net335 vssd1 vssd1 vccd1 vccd1 _07567_ sky130_fd_sc_hd__or2_2
XFILLER_0_57_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16494_ obsg2.obstacleArray\[24\] obsg2.obstacleArray\[25\] net459 vssd1 vssd1 vccd1
+ vccd1 _02173_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_80_2764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19282_ clknet_leaf_97_clk _00226_ net1450 vssd1 vssd1 vccd1 vccd1 control.body\[1104\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__17640__A2_N ag2.body\[167\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_2775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14835__B _01503_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18233_ obsg2.obstacleArray\[113\] _03755_ net527 vssd1 vssd1 vccd1 vccd1 _01364_
+ sky130_fd_sc_hd__o21a_1
XANTENNA__10660__A1 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15445_ ag2.body\[601\] net86 _01601_ ag2.body\[593\] vssd1 vssd1 vccd1 vccd1 _00731_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_61_2174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17211__B net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12657_ net677 _07533_ vssd1 vssd1 vccd1 vccd1 _07534_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_61_2185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_2196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09929__B _04661_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11608_ obsg2.obstacleArray\[31\] net632 net514 obsg2.obstacleArray\[27\] net1126
+ vssd1 vssd1 vccd1 vccd1 _06581_ sky130_fd_sc_hd__o221a_1
XFILLER_0_81_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18164_ _03600_ net37 obsg2.obstacleArray\[79\] vssd1 vssd1 vccd1 vccd1 _03721_ sky130_fd_sc_hd__a21oi_1
X_15376_ control.body\[667\] net69 _01594_ net2268 vssd1 vssd1 vccd1 vccd1 _00669_
+ sky130_fd_sc_hd__a22o_1
X_12588_ net336 _07494_ vssd1 vssd1 vccd1 vccd1 _07495_ sky130_fd_sc_hd__nor2_2
XFILLER_0_26_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16679__A1 net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14327_ net998 _04160_ ag2.body\[449\] net835 _08481_ vssd1 vssd1 vccd1 vccd1 _08488_
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_0_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17115_ ag2.body\[543\] net932 vssd1 vssd1 vccd1 vccd1 _02794_ sky130_fd_sc_hd__xor2_1
X_18095_ net351 _03610_ vssd1 vssd1 vccd1 vccd1 _03679_ sky130_fd_sc_hd__or2_1
X_11539_ obsg2.obstacleArray\[96\] obsg2.obstacleArray\[97\] obsg2.obstacleArray\[100\]
+ obsg2.obstacleArray\[101\] net1123 net510 vssd1 vssd1 vccd1 vccd1 _06512_ sky130_fd_sc_hd__mux4_1
XANTENNA__10156__A ag2.body\[62\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14851__A _08509_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_2693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold407 img_gen.tracker.frame\[284\] vssd1 vssd1 vccd1 vccd1 net1969 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__18323__A _04947_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_1303 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10963__A2 _05935_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold418 img_gen.tracker.frame\[560\] vssd1 vssd1 vccd1 vccd1 net1980 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17046_ ag2.body\[258\] net729 net695 ag2.body\[263\] _02724_ vssd1 vssd1 vccd1 vccd1
+ _02725_ sky130_fd_sc_hd__a221o_1
X_14258_ net986 _04005_ _04010_ net1013 vssd1 vssd1 vccd1 vccd1 _08419_ sky130_fd_sc_hd__a22o_1
Xhold429 img_gen.tracker.frame\[349\] vssd1 vssd1 vccd1 vccd1 net1991 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_74_2568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12165__A1 net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_2579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_1358 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17628__B1 net697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13209_ net676 _07794_ vssd1 vssd1 vccd1 vccd1 _07795_ sky130_fd_sc_hd__nor2_1
XFILLER_0_0_433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14189_ net998 ag2.body\[160\] vssd1 vssd1 vccd1 vccd1 _08350_ sky130_fd_sc_hd__or2_1
XFILLER_0_81_1384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12371__A net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout909 net910 vssd1 vssd1 vccd1 vccd1 net909 sky130_fd_sc_hd__clkbuf_4
X_18997_ clknet_leaf_2_clk img_gen.tracker.next_frame\[435\] net1248 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[435\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_104_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18726__CLK clknet_leaf_142_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15654__A2 net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17948_ net517 _03576_ vssd1 vssd1 vccd1 vccd1 _01258_ sky130_fd_sc_hd__nor2_1
XANTENNA__13665__A1 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1480 net1484 vssd1 vssd1 vccd1 vccd1 net1480 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_20_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1491 net1492 vssd1 vssd1 vccd1 vccd1 net1491 sky130_fd_sc_hd__buf_2
X_17879_ obsg2.obstacleCount\[3\] _04397_ vssd1 vssd1 vccd1 vccd1 _03519_ sky130_fd_sc_hd__or2_4
XFILLER_0_45_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11137__D _04470_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16603__B2 net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19618_ clknet_leaf_123_clk _00562_ net1407 vssd1 vssd1 vccd1 vccd1 control.body\[768\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_75_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13417__A1 net236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11434__B net1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19549_ clknet_leaf_115_clk _00493_ net1387 vssd1 vssd1 vccd1 vccd1 control.body\[843\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14223__A1_N net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09302_ _04321_ vssd1 vssd1 vccd1 vccd1 _04322_ sky130_fd_sc_hd__inv_2
XFILLER_0_53_1464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11979__B2 net564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_4432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16906__A2 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_135_4443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09233_ obsg2.obstacleArray\[1\] vssd1 vssd1 vccd1 vccd1 _04258_ sky130_fd_sc_hd__inv_2
XFILLER_0_8_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_4454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_1527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout230_A net233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_4307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12546__A net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_4318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_759 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11450__A net1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout328_A net331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_4329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_20_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09164_ ag2.body\[514\] vssd1 vssd1 vccd1 vccd1 _04189_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_20_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16960__B net955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_40_1557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09095_ ag2.body\[340\] vssd1 vssd1 vccd1 vccd1 _04120_ sky130_fd_sc_hd__inv_2
XFILLER_0_114_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10066__A net1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1237_A net1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20324_ clknet_leaf_43_clk _01220_ net1379 vssd1 vssd1 vccd1 vccd1 ag2.body\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__19501__CLK clknet_leaf_113_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold930 control.body\[975\] vssd1 vssd1 vccd1 vccd1 net2492 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_3060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold941 control.body\[881\] vssd1 vssd1 vccd1 vccd1 net2503 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout697_A net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_3071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold952 _00296_ vssd1 vssd1 vccd1 vccd1 net2514 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__17619__B1 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_4247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_3082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15893__A2 net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold963 control.body\[1031\] vssd1 vssd1 vccd1 vccd1 net2525 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13377__A _07539_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20255_ clknet_leaf_68_clk _01199_ net1498 vssd1 vssd1 vccd1 vccd1 ag2.body\[141\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_129_4258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold974 control.body\[932\] vssd1 vssd1 vccd1 vccd1 net2536 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1404_A net1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20359__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_4269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1025_X net1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold985 sound_gen.osc1.stayCount\[23\] vssd1 vssd1 vccd1 vccd1 net2547 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11903__A1 net438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_1475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold996 _00573_ vssd1 vssd1 vccd1 vccd1 net2558 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_53_1929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09572__A2 net1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_1486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20186_ clknet_leaf_88_clk _01130_ net1454 vssd1 vssd1 vccd1 vccd1 ag2.body\[200\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_38_1497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09997_ net1096 control.body\[733\] vssd1 vssd1 vccd1 vccd1 _04970_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout485_X net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout864_A net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10513__B net1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08948_ net1012 vssd1 vssd1 vccd1 vccd1 _03973_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_4_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09590__A net1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_826 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17398__A2 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1244 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10910_ _05875_ _05876_ _05877_ _05882_ vssd1 vssd1 vccd1 vccd1 _05883_ sky130_fd_sc_hd__or4_2
X_11890_ net576 _06861_ _06859_ vssd1 vssd1 vccd1 vccd1 _06862_ sky130_fd_sc_hd__a21oi_1
XANTENNA__13408__A1 net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_3410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16694__Y _02373_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11344__B net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10841_ ag2.body\[47\] net1048 vssd1 vssd1 vccd1 vccd1 _05814_ sky130_fd_sc_hd__xor2_1
XFILLER_0_79_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18347__A1 _04420_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14081__A1 net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14081__B2 net980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13840__A net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13560_ ssdec1.in\[2\] ssdec1.in\[0\] vssd1 vssd1 vccd1 vccd1 _07941_ sky130_fd_sc_hd__nor2_1
X_10772_ _05741_ _05742_ _05743_ _05744_ vssd1 vssd1 vccd1 vccd1 _05745_ sky130_fd_sc_hd__or4_1
X_12511_ net226 _07450_ _07451_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[17\]
+ sky130_fd_sc_hd__o21bai_1
XANTENNA__16453__S0 net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17031__B net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13491_ net666 _07908_ vssd1 vssd1 vccd1 vccd1 _07909_ sky130_fd_sc_hd__nor2_1
XFILLER_0_81_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_97_3269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15230_ control.body\[794\] net96 _01577_ net2235 vssd1 vssd1 vccd1 vccd1 _00540_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_136_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_114_3804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12442_ _06658_ _07255_ _07287_ _07402_ vssd1 vssd1 vccd1 vccd1 _07403_ sky130_fd_sc_hd__or4_1
XFILLER_0_63_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_114_3815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_1660 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16870__B net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15161_ control.body\[861\] net98 _01569_ control.body\[853\] vssd1 vssd1 vccd1 vccd1
+ _00479_ sky130_fd_sc_hd__a22o_1
XFILLER_0_133_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12373_ img_gen.updater.commands.rR1.rainbowRNG\[9\] _07319_ _07334_ _07338_ _07297_
+ vssd1 vssd1 vccd1 vccd1 _07339_ sky130_fd_sc_hd__a221o_1
XFILLER_0_1_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12743__X _07575_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_872 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__08940__Y _03965_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18143__A net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16756__S1 net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19181__CLK clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14112_ net1025 ag2.body\[573\] vssd1 vssd1 vccd1 vccd1 _08273_ sky130_fd_sc_hd__xor2_1
XFILLER_0_107_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11324_ ag2.body\[556\] net1132 vssd1 vssd1 vccd1 vccd1 _06297_ sky130_fd_sc_hd__xor2_1
X_15092_ control.body\[927\] net147 _01562_ net2358 vssd1 vssd1 vccd1 vccd1 _00417_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_65_1368 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12147__A1 _07105_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17982__A net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14043_ _08192_ _08201_ _08202_ _08203_ vssd1 vssd1 vccd1 vccd1 _08204_ sky130_fd_sc_hd__or4_1
X_18920_ clknet_leaf_145_clk img_gen.tracker.next_frame\[358\] net1253 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[358\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_103_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11255_ net1151 control.body\[771\] vssd1 vssd1 vccd1 vccd1 _06228_ sky130_fd_sc_hd__or2_1
XFILLER_0_120_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10158__B1 net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12191__A net1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19877__RESET_B net1415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10206_ net1107 control.body\[997\] vssd1 vssd1 vccd1 vccd1 _05179_ sky130_fd_sc_hd__xor2_1
X_18851_ clknet_leaf_18_clk img_gen.tracker.next_frame\[289\] net1319 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[289\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__11519__B net1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_108_3608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11186_ _04056_ net1176 net1056 _04059_ _06154_ vssd1 vssd1 vccd1 vccd1 _06159_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_108_3619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17802_ net696 _03470_ _03472_ vssd1 vssd1 vccd1 vccd1 _01217_ sky130_fd_sc_hd__a21oi_1
X_10137_ net1130 control.body\[820\] vssd1 vssd1 vccd1 vccd1 _05110_ sky130_fd_sc_hd__xor2_1
X_18782_ clknet_leaf_12_clk img_gen.tracker.next_frame\[220\] net1285 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[220\] sky130_fd_sc_hd__dfrtp_1
X_15994_ net1755 control.body_update.direction\[0\] net223 vssd1 vssd1 vccd1 vccd1
+ _01206_ sky130_fd_sc_hd__mux2_1
XANTENNA__18899__CLK clknet_leaf_144_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14844__B1 _08783_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17733_ _02725_ _02731_ _03411_ _02578_ vssd1 vssd1 vccd1 vccd1 _03412_ sky130_fd_sc_hd__o211a_2
X_10068_ net1049 control.body\[719\] vssd1 vssd1 vccd1 vccd1 _05041_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_13_Right_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14945_ control.body\[1053\] net174 _01545_ net2303 vssd1 vssd1 vccd1 vccd1 _00287_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__17206__B net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11180__A_N net1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17389__A2 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17664_ ag2.body\[108\] net713 net708 ag2.body\[109\] _03335_ vssd1 vssd1 vccd1 vccd1
+ _03343_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_82_2815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14876_ _04859_ _01536_ vssd1 vssd1 vccd1 vccd1 _01538_ sky130_fd_sc_hd__and2b_2
XTAP_TAPCELL_ROW_67_2361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_67_2372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19403_ clknet_leaf_103_clk _00347_ net1431 vssd1 vssd1 vccd1 vccd1 control.body\[985\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09005__A ag2.body\[122\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16615_ obsg2.obstacleArray\[43\] net449 net390 _02293_ vssd1 vssd1 vccd1 vccd1 _02294_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_98_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20364__RESET_B net1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13827_ _04270_ _08110_ vssd1 vssd1 vccd1 vccd1 _08124_ sky130_fd_sc_hd__or2_2
X_17595_ net926 net924 _03013_ vssd1 vssd1 vccd1 vccd1 _03274_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_63_2236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_2247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_1150 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_2258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19334_ clknet_leaf_103_clk net2469 net1432 vssd1 vssd1 vccd1 vccd1 control.body\[1060\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09499__X _04472_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16546_ obsg2.obstacleArray\[97\] net449 net394 _02224_ vssd1 vssd1 vccd1 vccd1 _02225_
+ sky130_fd_sc_hd__o211a_1
X_13758_ img_gen.updater.commands.count\[4\] img_gen.updater.commands.count\[3\] _08068_
+ vssd1 vssd1 vccd1 vccd1 _08075_ sky130_fd_sc_hd__and3_1
XFILLER_0_50_1648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_1571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12709_ net305 _07558_ vssd1 vssd1 vccd1 vccd1 _07559_ sky130_fd_sc_hd__nor2_1
X_19265_ clknet_leaf_71_clk _00209_ net1503 vssd1 vssd1 vccd1 vccd1 ag2.body\[128\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_14_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11830__B1 net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16477_ obsg2.obstacleArray\[34\] obsg2.obstacleArray\[35\] net452 vssd1 vssd1 vccd1
+ vccd1 _02156_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_14_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12366__A net241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09659__B net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13689_ net899 net434 _08030_ _08022_ vssd1 vssd1 vccd1 vccd1 track.nextCurrScore\[6\]
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_14_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18216_ _03658_ net40 vssd1 vssd1 vccd1 vccd1 _03747_ sky130_fd_sc_hd__nor2_1
XANTENNA__20356__Q obsg2.obstacleCount\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15428_ ag2.body\[618\] net84 _01599_ ag2.body\[610\] vssd1 vssd1 vccd1 vccd1 _00716_
+ sky130_fd_sc_hd__a22o_1
X_19196_ clknet_leaf_53_clk _00140_ net1455 vssd1 vssd1 vccd1 vccd1 ag2.body\[59\]
+ sky130_fd_sc_hd__dfrtp_4
XPHY_EDGE_ROW_22_Right_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11701__C _06671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11189__A2 net1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18147_ net529 _03712_ vssd1 vssd1 vccd1 vccd1 _01321_ sky130_fd_sc_hd__and2_1
XFILLER_0_5_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15359_ control.body\[684\] net75 _01592_ net2377 vssd1 vssd1 vccd1 vccd1 _00654_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_14_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11594__C1 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10936__A2 _04982_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold204 img_gen.tracker.frame\[186\] vssd1 vssd1 vccd1 vccd1 net1766 sky130_fd_sc_hd__dlygate4sd3_1
Xhold215 img_gen.tracker.frame\[360\] vssd1 vssd1 vccd1 vccd1 net1777 sky130_fd_sc_hd__dlygate4sd3_1
X_18078_ net300 _03597_ vssd1 vssd1 vccd1 vccd1 _03668_ sky130_fd_sc_hd__nand2_1
Xhold226 img_gen.tracker.frame\[404\] vssd1 vssd1 vccd1 vccd1 net1788 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_48_1588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold237 img_gen.tracker.frame\[511\] vssd1 vssd1 vccd1 vccd1 net1799 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_61_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09920_ ag2.body\[313\] net781 net752 ag2.body\[318\] _04892_ vssd1 vssd1 vccd1 vccd1
+ _04893_ sky130_fd_sc_hd__a221o_1
XANTENNA__13197__A net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold248 img_gen.tracker.frame\[535\] vssd1 vssd1 vccd1 vccd1 net1810 sky130_fd_sc_hd__dlygate4sd3_1
X_17029_ _04145_ net953 net701 ag2.body\[406\] _02707_ vssd1 vssd1 vccd1 vccd1 _02708_
+ sky130_fd_sc_hd__a221o_1
Xhold259 img_gen.tracker.frame\[515\] vssd1 vssd1 vccd1 vccd1 net1821 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20040_ clknet_leaf_68_clk _00984_ net1494 vssd1 vssd1 vccd1 vccd1 ag2.body\[358\]
+ sky130_fd_sc_hd__dfrtp_4
Xfanout706 net708 vssd1 vssd1 vccd1 vccd1 net706 sky130_fd_sc_hd__buf_4
XFILLER_0_21_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout717 _04265_ vssd1 vssd1 vccd1 vccd1 net717 sky130_fd_sc_hd__buf_4
X_09851_ net1205 _04249_ control.body\[975\] net745 _04823_ vssd1 vssd1 vccd1 vccd1
+ _04824_ sky130_fd_sc_hd__a221o_1
XANTENNA__11429__B net1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout728 net729 vssd1 vssd1 vccd1 vccd1 net728 sky130_fd_sc_hd__buf_4
XANTENNA__11897__B1 net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_4100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_1480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10333__B net1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_4111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout739 net741 vssd1 vssd1 vccd1 vccd1 net739 sky130_fd_sc_hd__buf_4
XANTENNA__15627__A2 net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09782_ net1087 control.body\[950\] vssd1 vssd1 vccd1 vccd1 _04755_ sky130_fd_sc_hd__or2_1
XFILLER_0_77_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_31_Right_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout180_A net182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout278_A net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11445__A net1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16955__B net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_137_4505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19054__CLK clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16447__S net456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_137_4516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout445_A _02214_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15260__B1 net50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18329__A1 net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14756__A net1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_46_1722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13660__A net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1187_A net1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_46_1733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12074__B1 net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_27_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12547__Y _07472_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__20031__CLK clknet_leaf_66_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout612_A _06475_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_23_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15012__B1 _01553_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout233_X net233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_40_Right_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1354_A net1355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_23_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09216_ control.body\[775\] vssd1 vssd1 vccd1 vccd1 _04241_ sky130_fd_sc_hd__inv_2
XFILLER_0_9_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17786__B net1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16760__B1 net489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_3122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09147_ ag2.body\[479\] vssd1 vssd1 vccd1 vccd1 _04172_ sky130_fd_sc_hd__inv_2
XFILLER_0_126_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout400_X net400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16182__S net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_3133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_3144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1142_X net1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_308 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17304__A2 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09585__A net1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09078_ ag2.body\[312\] vssd1 vssd1 vccd1 vccd1 _04103_ sky130_fd_sc_hd__inv_2
XANTENNA__16512__B1 net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout981_A net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_544 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20307_ clknet_leaf_70_clk net1563 net1499 vssd1 vssd1 vccd1 vccd1 obsmode.sOBSMODE.pb_1
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__15866__A2 net161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1244 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold760 control.body\[719\] vssd1 vssd1 vccd1 vccd1 net2322 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10524__A net1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19970__RESET_B net1470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout93_A net100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold771 control.body\[655\] vssd1 vssd1 vccd1 vccd1 net2333 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09872__X _04845_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold782 control.body\[988\] vssd1 vssd1 vccd1 vccd1 net2344 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__18265__B1 net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11040_ net1085 control.body\[1046\] vssd1 vssd1 vccd1 vccd1 _06013_ sky130_fd_sc_hd__nand2b_1
X_20238_ clknet_leaf_65_clk _01182_ net1476 vssd1 vssd1 vccd1 vccd1 ag2.body\[156\]
+ sky130_fd_sc_hd__dfrtp_4
Xhold793 control.body\[838\] vssd1 vssd1 vccd1 vccd1 net2355 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11888__B1 net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout867_X net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10243__B net1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16276__C1 _01912_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15618__A2 net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17952__D net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13835__A net677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20169_ clknet_leaf_95_clk _01113_ net1441 vssd1 vssd1 vccd1 vccd1 ag2.body\[231\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_137_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17026__B net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12991_ net341 _07512_ vssd1 vssd1 vccd1 vccd1 _07691_ sky130_fd_sc_hd__nor2_1
XFILLER_0_137_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11355__A net1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14730_ net845 ag2.body\[112\] ag2.body\[119\] net796 _08890_ vssd1 vssd1 vccd1 vccd1
+ _08891_ sky130_fd_sc_hd__a221o_1
XFILLER_0_98_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_807 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11942_ _06911_ _06913_ net574 vssd1 vssd1 vccd1 vccd1 _06914_ sky130_fd_sc_hd__mux2_1
XANTENNA__16579__B1 net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13273__C _07813_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13841__Y _08131_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14661_ net1021 ag2.body\[526\] vssd1 vssd1 vccd1 vccd1 _08822_ sky130_fd_sc_hd__or2_1
X_11873_ img_gen.tracker.frame\[241\] net615 net598 img_gen.tracker.frame\[244\] vssd1
+ vssd1 vccd1 vccd1 _06845_ sky130_fd_sc_hd__o22a_1
XANTENNA__16357__S net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13612_ _07958_ net220 _07983_ vssd1 vssd1 vccd1 vccd1 control.divider.next_count\[3\]
+ sky130_fd_sc_hd__and3b_1
X_16400_ _02077_ _02078_ net403 vssd1 vssd1 vccd1 vccd1 _02079_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10824_ _05791_ _05792_ _05793_ _05796_ vssd1 vssd1 vccd1 vccd1 _05797_ sky130_fd_sc_hd__or4_1
X_14592_ net829 ag2.body\[82\] _08745_ _08752_ vssd1 vssd1 vccd1 vccd1 _08753_ sky130_fd_sc_hd__a211o_1
X_17380_ ag2.body\[492\] net962 vssd1 vssd1 vccd1 vccd1 _03059_ sky130_fd_sc_hd__or2_1
XANTENNA__19547__CLK clknet_leaf_115_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_931 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18852__RESET_B net1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16331_ obsg2.obstacleArray\[76\] obsg2.obstacleArray\[77\] net406 vssd1 vssd1 vccd1
+ vccd1 _02010_ sky130_fd_sc_hd__mux2_1
X_13543_ net2045 net655 _07927_ _07928_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[572\]
+ sky130_fd_sc_hd__a31o_1
XANTENNA__17977__A net45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10755_ net1131 control.body\[892\] vssd1 vssd1 vccd1 vccd1 _05728_ sky130_fd_sc_hd__nand2_1
XANTENNA__12186__A net1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15003__B1 _01552_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16262_ _01939_ _01940_ net418 vssd1 vssd1 vccd1 vccd1 _01941_ sky130_fd_sc_hd__mux2_1
XANTENNA__20524__CLK clknet_leaf_93_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19050_ clknet_leaf_10_clk img_gen.tracker.next_frame\[488\] net1275 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[488\] sky130_fd_sc_hd__dfrtp_1
X_13474_ net276 _07900_ _07901_ net1752 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[530\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_129_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10686_ ag2.body\[150\] net1088 vssd1 vssd1 vccd1 vccd1 _05659_ sky130_fd_sc_hd__or2_1
X_18001_ obsg2.obstacleArray\[21\] _03615_ net533 vssd1 vssd1 vccd1 vccd1 _01272_
+ sky130_fd_sc_hd__o21a_1
X_15213_ net2578 net92 _01575_ control.body\[803\] vssd1 vssd1 vccd1 vccd1 _00525_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_10_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12425_ _06556_ _06558_ _06505_ vssd1 vssd1 vccd1 vccd1 _07387_ sky130_fd_sc_hd__a21bo_1
XANTENNA__18571__CLK clknet_leaf_15_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16193_ obsg2.obstacleArray\[46\] net421 vssd1 vssd1 vccd1 vccd1 _01872_ sky130_fd_sc_hd__or2_1
XFILLER_0_22_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11576__C1 net1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15144_ net2633 net107 _01567_ control.body\[870\] vssd1 vssd1 vccd1 vccd1 _00464_
+ sky130_fd_sc_hd__a22o_1
X_12356_ _07251_ _06506_ vssd1 vssd1 vccd1 vccd1 _07323_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_51_976 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_2040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_853 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11591__A2 obsg2.obstacleArray\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11307_ ag2.body\[275\] net1164 vssd1 vssd1 vccd1 vccd1 _06280_ sky130_fd_sc_hd__xor2_1
X_19952_ clknet_leaf_45_clk _00896_ net1379 vssd1 vssd1 vccd1 vccd1 ag2.body\[446\]
+ sky130_fd_sc_hd__dfrtp_4
X_15075_ _04552_ _04586_ net65 vssd1 vssd1 vccd1 vccd1 _01561_ sky130_fd_sc_hd__and3_2
XFILLER_0_26_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12287_ net687 _07246_ _07255_ _07230_ vssd1 vssd1 vccd1 vccd1 _07257_ sky130_fd_sc_hd__o31a_1
XANTENNA__10434__A net1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14026_ net798 ag2.body\[30\] _03985_ net1006 vssd1 vssd1 vccd1 vccd1 _08187_ sky130_fd_sc_hd__a22o_1
X_18903_ clknet_leaf_144_clk img_gen.tracker.next_frame\[341\] net1251 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[341\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__11249__B net1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11238_ ag2.body\[193\] net1208 vssd1 vssd1 vccd1 vccd1 _06211_ sky130_fd_sc_hd__nand2_1
X_19883_ clknet_leaf_84_clk _00827_ net1483 vssd1 vssd1 vccd1 vccd1 ag2.body\[505\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__11879__B1 net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10153__B net1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16267__C1 net368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18834_ clknet_leaf_4_clk img_gen.tracker.next_frame\[272\] net1263 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[272\] sky130_fd_sc_hd__dfrtp_1
X_11169_ net1050 control.body\[783\] vssd1 vssd1 vccd1 vccd1 _06142_ sky130_fd_sc_hd__or2_1
XFILLER_0_93_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_69_2423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_2434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18765_ clknet_leaf_16_clk img_gen.tracker.next_frame\[203\] net1318 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[203\] sky130_fd_sc_hd__dfrtp_1
X_15977_ _01659_ _01662_ ag2.body\[0\] vssd1 vssd1 vccd1 vccd1 _01202_ sky130_fd_sc_hd__mux2_1
XANTENNA__14293__A1 net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14293__B2 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19205__Q ag2.body\[68\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17716_ obsg2.obstacleArray\[138\] obsg2.obstacleArray\[139\] net426 vssd1 vssd1
+ vccd1 vccd1 _03395_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_65_2309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1261 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14928_ control.body\[1070\] net170 _01543_ net2184 vssd1 vssd1 vccd1 vccd1 _00272_
+ sky130_fd_sc_hd__a22o_1
X_18696_ clknet_leaf_11_clk img_gen.tracker.next_frame\[134\] net1281 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[134\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_72_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17647_ ag2.body\[37\] net946 vssd1 vssd1 vccd1 vccd1 _03326_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_8_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14859_ _08165_ _08171_ _08403_ vssd1 vssd1 vccd1 vccd1 _01530_ sky130_fd_sc_hd__o21a_1
XPHY_EDGE_ROW_11_Left_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14576__A net1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15242__B1 _01578_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17782__A2 net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13480__A net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_931 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17578_ ag2.body\[341\] net954 vssd1 vssd1 vccd1 vccd1 _03257_ sky130_fd_sc_hd__xor2_1
XANTENNA__15793__A1 ag2.body\[303\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16990__B1 net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15793__B2 ag2.body\[295\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19317_ clknet_leaf_104_clk _00261_ net1433 vssd1 vssd1 vccd1 vccd1 control.body\[1075\]
+ sky130_fd_sc_hd__dfrtp_1
X_16529_ _01700_ _02207_ vssd1 vssd1 vccd1 vccd1 _02208_ sky130_fd_sc_hd__nor2_1
XANTENNA__11712__B net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18914__CLK clknet_leaf_142_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10609__A net1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_0_clk_X clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19248_ clknet_leaf_84_clk _00192_ net1481 vssd1 vssd1 vccd1 vccd1 ag2.body\[111\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_2_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16742__B1 net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09001_ ag2.body\[112\] vssd1 vssd1 vccd1 vccd1 _04026_ sky130_fd_sc_hd__inv_2
XFILLER_0_61_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19179_ clknet_leaf_20_clk _00123_ net1365 vssd1 vssd1 vccd1 vccd1 ag2.body\[42\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_131_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12824__A net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11567__C1 net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_35_1401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18247__B1 net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09903_ _04863_ _04870_ _04875_ _04858_ _04831_ vssd1 vssd1 vccd1 vccd1 _04876_ sky130_fd_sc_hd__o32a_1
XTAP_TAPCELL_ROW_6_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout503 _01708_ vssd1 vssd1 vccd1 vccd1 net503 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_6_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11159__B net1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout514 net515 vssd1 vssd1 vccd1 vccd1 net514 sky130_fd_sc_hd__clkbuf_4
Xfanout525 net528 vssd1 vssd1 vccd1 vccd1 net525 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_6_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16258__C1 net369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout395_A net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1547 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12531__A1 net283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20023_ clknet_leaf_58_clk _00967_ net1471 vssd1 vssd1 vccd1 vccd1 ag2.body\[373\]
+ sky130_fd_sc_hd__dfrtp_4
X_09834_ net1107 control.body\[925\] vssd1 vssd1 vccd1 vccd1 _04807_ sky130_fd_sc_hd__nand2_1
Xfanout547 net553 vssd1 vssd1 vccd1 vccd1 net547 sky130_fd_sc_hd__clkbuf_4
XANTENNA__16849__A1_N net704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18262__A3 net48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1102_A net1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout558 net559 vssd1 vssd1 vccd1 vccd1 net558 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_96_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout569 net570 vssd1 vssd1 vccd1 vccd1 net569 sky130_fd_sc_hd__buf_2
XANTENNA__16273__A2 net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09765_ _04734_ _04735_ _04736_ _04737_ vssd1 vssd1 vccd1 vccd1 _04738_ sky130_fd_sc_hd__or4_1
XANTENNA__14284__A1 net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout562_A net567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout183_X net183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14284__B2 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11175__A net1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15481__B1 _01605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09696_ net641 _04493_ vssd1 vssd1 vccd1 vccd1 _04669_ sky130_fd_sc_hd__nor2_1
XFILLER_0_83_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout350_X net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10845__B2 net1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14486__A net1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1092_X net1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout827_A net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout448_X net448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20547__CLK clknet_leaf_105_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12047__B1 net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16981__B1 net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15784__B2 ag2.body\[303\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12598__A1 net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_3320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18594__CLK clknet_leaf_13_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout615_X net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1357_X net1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10540_ ag2.body\[231\] net1061 vssd1 vssd1 vccd1 vccd1 _05513_ sky130_fd_sc_hd__nand2_1
XANTENNA__16733__B1 net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10238__B net1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13465__B_N _07486_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10471_ net1084 control.body\[1014\] vssd1 vssd1 vccd1 vccd1 _05444_ sky130_fd_sc_hd__xor2_1
XFILLER_0_134_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11558__C1 net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12210_ img_gen.updater.commands.mode\[1\] img_gen.updater.commands.mode\[0\] img_gen.updater.commands.mode\[2\]
+ vssd1 vssd1 vccd1 vccd1 _07182_ sky130_fd_sc_hd__and3b_1
X_13190_ net383 _07615_ vssd1 vssd1 vccd1 vccd1 _07785_ sky130_fd_sc_hd__nor2_1
XFILLER_0_60_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout984_X net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16497__C1 _02076_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12770__A1 net235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12141_ img_gen.tracker.frame\[516\] net620 net583 img_gen.tracker.frame\[525\] _07112_
+ vssd1 vssd1 vccd1 vccd1 _07113_ sky130_fd_sc_hd__o221a_1
XFILLER_0_103_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11069__B net1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12072_ img_gen.tracker.frame\[96\] net629 net611 img_gen.tracker.frame\[99\] _07043_
+ vssd1 vssd1 vccd1 vccd1 _07044_ sky130_fd_sc_hd__a221o_1
Xhold590 control.body\[1117\] vssd1 vssd1 vccd1 vccd1 net2152 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1051 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11637__X _06610_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15900_ ag2.body\[207\] net133 _01650_ ag2.body\[199\] vssd1 vssd1 vccd1 vccd1 _01137_
+ sky130_fd_sc_hd__a22o_1
X_11023_ ag2.body\[595\] net1147 vssd1 vssd1 vccd1 vccd1 _05996_ sky130_fd_sc_hd__nand2_1
XANTENNA__09762__B net1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16880_ ag2.body\[22\] net937 vssd1 vssd1 vccd1 vccd1 _02559_ sky130_fd_sc_hd__xor2_1
XANTENNA__13284__B _07827_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15831_ ag2.body\[257\] net204 net49 ag2.body\[249\] vssd1 vssd1 vccd1 vccd1 _01075_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__10701__B net1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14948__X _01546_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18550_ clknet_leaf_132_clk _00076_ net1297 vssd1 vssd1 vccd1 vccd1 ag2.y\[2\] sky130_fd_sc_hd__dfrtp_1
X_15762_ ag2.body\[323\] net215 _01636_ ag2.body\[315\] vssd1 vssd1 vccd1 vccd1 _01013_
+ sky130_fd_sc_hd__a22o_1
X_12974_ net279 _07681_ _07682_ net1692 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[248\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_137_1457 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16595__B net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17501_ ag2.body\[236\] net965 vssd1 vssd1 vccd1 vccd1 _03180_ sky130_fd_sc_hd__xor2_1
X_14713_ net993 _04119_ ag2.body\[340\] net816 _08873_ vssd1 vssd1 vccd1 vccd1 _08874_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_115_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11925_ img_gen.tracker.frame\[310\] net591 net551 img_gen.tracker.frame\[307\] vssd1
+ vssd1 vccd1 vccd1 _06897_ sky130_fd_sc_hd__o22ai_1
X_18481_ net1515 net1509 vssd1 vssd1 vccd1 vccd1 _00012_ sky130_fd_sc_hd__or2_1
X_15693_ ag2.body\[391\] net137 _01616_ ag2.body\[383\] vssd1 vssd1 vccd1 vccd1 _00953_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__16087__S net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14027__B2 net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17432_ ag2.body\[150\] net701 net693 ag2.body\[151\] vssd1 vssd1 vccd1 vccd1 _03111_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_16_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14644_ ag2.body\[519\] net794 net984 _04189_ vssd1 vssd1 vccd1 vccd1 _08805_ sky130_fd_sc_hd__a2bb2o_1
X_11856_ img_gen.tracker.frame\[235\] net552 vssd1 vssd1 vccd1 vccd1 _06828_ sky130_fd_sc_hd__or2_1
XANTENNA__16972__B1 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12589__A1 _07431_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10807_ _05776_ _05777_ _05778_ _05779_ vssd1 vssd1 vccd1 vccd1 _05780_ sky130_fd_sc_hd__or4_1
X_17363_ _03007_ _03032_ vssd1 vssd1 vccd1 vccd1 _03042_ sky130_fd_sc_hd__xnor2_1
X_14575_ net973 ag2.body\[491\] vssd1 vssd1 vccd1 vccd1 _08736_ sky130_fd_sc_hd__or2_1
XFILLER_0_83_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11787_ img_gen.tracker.frame\[353\] net598 net580 img_gen.tracker.frame\[359\] vssd1
+ vssd1 vccd1 vccd1 _06759_ sky130_fd_sc_hd__o22a_1
XANTENNA__10429__A net1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13250__A2 net648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17516__A2 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19102_ clknet_leaf_0_clk img_gen.tracker.next_frame\[540\] net1240 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[540\] sky130_fd_sc_hd__dfrtp_1
X_16314_ obsg2.obstacleArray\[109\] net413 _01992_ net418 vssd1 vssd1 vccd1 vccd1
+ _01993_ sky130_fd_sc_hd__o211a_1
XFILLER_0_83_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11261__A1 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10738_ ag2.body\[496\] net1233 vssd1 vssd1 vccd1 vccd1 _05711_ sky130_fd_sc_hd__xor2_1
XFILLER_0_27_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13526_ net2091 net655 _07921_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[562\]
+ sky130_fd_sc_hd__and3_1
XFILLER_0_125_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17294_ ag2.body\[348\] net966 vssd1 vssd1 vccd1 vccd1 _02973_ sky130_fd_sc_hd__nand2_1
XANTENNA__11261__B2 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10148__B net1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11959__S net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19033_ clknet_leaf_6_clk img_gen.tracker.next_frame\[471\] net1264 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[471\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_58_2102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16245_ obsg2.obstacleArray\[46\] obsg2.obstacleArray\[47\] net404 vssd1 vssd1 vccd1
+ vccd1 _01924_ sky130_fd_sc_hd__mux2_1
X_13457_ net235 _07894_ _07895_ net1613 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[519\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__09937__B net1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10669_ net1227 _04245_ control.body\[887\] net746 _05636_ vssd1 vssd1 vccd1 vccd1
+ _05642_ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_124_Right_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15020__A _04551_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12408_ _06626_ _06628_ _07351_ _07370_ vssd1 vssd1 vccd1 vccd1 _07371_ sky130_fd_sc_hd__a31o_1
X_16176_ obsg2.obstacleArray\[54\] net424 vssd1 vssd1 vccd1 vccd1 _01855_ sky130_fd_sc_hd__or2_1
X_13388_ net670 _07868_ vssd1 vssd1 vccd1 vccd1 _07869_ sky130_fd_sc_hd__nor2_1
XFILLER_0_80_1405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_1536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16488__C1 net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11564__A2 net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15955__A _05237_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15127_ net2662 net104 _01565_ control.body\[887\] vssd1 vssd1 vccd1 vccd1 _00449_
+ sky130_fd_sc_hd__a22o_1
X_12339_ net435 _07305_ vssd1 vssd1 vccd1 vccd1 _07306_ sky130_fd_sc_hd__and2_2
XANTENNA__18331__A net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09509__A2 net1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19935_ clknet_leaf_47_clk _00879_ net1375 vssd1 vssd1 vccd1 vccd1 ag2.body\[461\]
+ sky130_fd_sc_hd__dfrtp_4
X_15058_ net2575 net149 _01559_ net2291 vssd1 vssd1 vccd1 vccd1 _00386_ sky130_fd_sc_hd__a22o_1
XFILLER_0_103_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11316__A2 _06276_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14009_ net837 ag2.body\[505\] ag2.body\[508\] net814 _08169_ vssd1 vssd1 vccd1 vccd1
+ _08170_ sky130_fd_sc_hd__a221o_1
XANTENNA__13475__A net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19866_ clknet_leaf_95_clk _00810_ net1440 vssd1 vssd1 vccd1 vccd1 ag2.body\[520\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_128_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18817_ clknet_leaf_2_clk img_gen.tracker.next_frame\[255\] net1249 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[255\] sky130_fd_sc_hd__dfrtp_1
X_19797_ clknet_leaf_128_clk _00741_ net1328 vssd1 vssd1 vccd1 vccd1 ag2.body\[595\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__15463__B1 _01603_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09550_ net1217 control.body\[720\] vssd1 vssd1 vccd1 vccd1 _04523_ sky130_fd_sc_hd__xor2_1
X_18748_ clknet_leaf_143_clk img_gen.tracker.next_frame\[186\] net1256 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[186\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_95_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09481_ ag2.body\[470\] net748 net744 ag2.body\[471\] vssd1 vssd1 vccd1 vccd1 _04454_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_76_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18679_ clknet_leaf_27_clk img_gen.tracker.next_frame\[117\] net1339 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[117\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_884 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout143_A net144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09687__X _04660_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16715__B1 net482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20572_ clknet_leaf_106_clk _01430_ _00036_ vssd1 vssd1 vccd1 vccd1 sound_gen.dac1.dacCount\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__18180__A2 _03703_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_293 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10058__B net1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16191__A1 _01743_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout310_A net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout408_A _01902_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1052_A net1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11004__A1 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09748__A2 net788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12201__B1 net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11004__B2 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12752__A1 net236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15865__A _05517_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17783__C net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1317_A net1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout300 net301 vssd1 vssd1 vccd1 vccd1 net300 sky130_fd_sc_hd__buf_2
Xfanout311 _07429_ vssd1 vssd1 vccd1 vccd1 net311 sky130_fd_sc_hd__clkbuf_4
Xfanout1309 net1310 vssd1 vssd1 vccd1 vccd1 net1309 sky130_fd_sc_hd__buf_2
XANTENNA_fanout777_A net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12504__A1 net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout322 track.nextHighScore\[5\] vssd1 vssd1 vccd1 vccd1 net322 sky130_fd_sc_hd__buf_1
XFILLER_0_121_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10361__X _05334_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout333 _07423_ vssd1 vssd1 vccd1 vccd1 net333 sky130_fd_sc_hd__buf_2
Xfanout344 _07308_ vssd1 vssd1 vccd1 vccd1 net344 sky130_fd_sc_hd__buf_2
XANTENNA_fanout1105_X net1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout355 _01699_ vssd1 vssd1 vccd1 vccd1 net355 sky130_fd_sc_hd__buf_2
XANTENNA__19392__CLK clknet_leaf_102_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout366 _02067_ vssd1 vssd1 vccd1 vccd1 net366 sky130_fd_sc_hd__buf_4
XFILLER_0_103_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20006_ clknet_leaf_59_clk _00950_ net1472 vssd1 vssd1 vccd1 vccd1 ag2.body\[388\]
+ sky130_fd_sc_hd__dfrtp_4
Xfanout377 net379 vssd1 vssd1 vccd1 vccd1 net377 sky130_fd_sc_hd__buf_2
XANTENNA__09920__A2 net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09817_ net769 control.body\[1051\] control.body\[1053\] net755 _04789_ vssd1 vssd1
+ vccd1 vccd1 _04790_ sky130_fd_sc_hd__o221a_1
XANTENNA__14257__A1 net815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1456 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout388 _06675_ vssd1 vssd1 vccd1 vccd1 net388 sky130_fd_sc_hd__buf_2
XANTENNA_fanout944_A net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout399 net400 vssd1 vssd1 vccd1 vccd1 net399 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout565_X net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14257__B2 net802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15454__B1 _01602_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09748_ ag2.body\[352\] net788 net763 ag2.body\[356\] _04714_ vssd1 vssd1 vccd1 vccd1
+ _04721_ sky130_fd_sc_hd__o221a_1
XANTENNA_fanout56_A net62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout732_X net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09679_ _04648_ _04649_ _04650_ _04651_ vssd1 vssd1 vccd1 vccd1 _04652_ sky130_fd_sc_hd__a22o_1
XANTENNA__14009__A1 net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16983__X _02662_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14009__B2 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15206__B1 _01574_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_979 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11710_ img_gen.tracker.frame\[314\] net619 net607 img_gen.tracker.frame\[317\] vssd1
+ vssd1 vccd1 vccd1 _06682_ sky130_fd_sc_hd__o22a_1
XANTENNA__10294__A2 net1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12690_ net259 _07549_ _07550_ net2098 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[97\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_90_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11352__B net1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11641_ obsg2.obstacleArray\[135\] net632 net513 obsg2.obstacleArray\[131\] net507
+ vssd1 vssd1 vccd1 vccd1 _06614_ sky130_fd_sc_hd__o221a_1
XFILLER_0_65_865 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14360_ _08517_ _08518_ _08519_ _08520_ vssd1 vssd1 vccd1 vccd1 _08521_ sky130_fd_sc_hd__or4_2
XFILLER_0_108_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09597__X _04570_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11572_ net504 _06544_ _06543_ net475 vssd1 vssd1 vccd1 vccd1 _06545_ sky130_fd_sc_hd__o211a_1
XANTENNA__08942__A ag2.body\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16706__B1 net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18135__B net41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13311_ net225 _07837_ vssd1 vssd1 vccd1 vccd1 _07838_ sky130_fd_sc_hd__nor2_1
XFILLER_0_107_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11794__A2 net587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10523_ _05419_ _05449_ _05473_ _05495_ vssd1 vssd1 vccd1 vccd1 _05496_ sky130_fd_sc_hd__or4_1
X_14291_ net996 ag2.body\[472\] vssd1 vssd1 vccd1 vccd1 _08452_ sky130_fd_sc_hd__xor2_1
XANTENNA__09757__B net1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10536__X _05509_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16030_ _01678_ _01682_ vssd1 vssd1 vccd1 vccd1 _01709_ sky130_fd_sc_hd__xor2_4
X_13242_ _07434_ _07807_ net651 vssd1 vssd1 vccd1 vccd1 _07810_ sky130_fd_sc_hd__o21a_1
X_10454_ ag2.body\[450\] net1176 vssd1 vssd1 vccd1 vccd1 _05427_ sky130_fd_sc_hd__or2_1
XANTENNA__13279__B _07825_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12614__D _07508_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13173_ net277 _07775_ _07776_ net1715 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[353\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_131_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19232__RESET_B net1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10385_ _05352_ _05357_ _05347_ vssd1 vssd1 vccd1 vccd1 _05358_ sky130_fd_sc_hd__or3b_4
XFILLER_0_42_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18151__A net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12124_ img_gen.tracker.frame\[540\] net613 net579 img_gen.tracker.frame\[549\] _07094_
+ vssd1 vssd1 vccd1 vccd1 _07096_ sky130_fd_sc_hd__o221a_1
XANTENNA__19735__CLK clknet_leaf_132_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17981_ obsg2.obstacleArray\[15\] _03601_ net523 vssd1 vssd1 vccd1 vccd1 _01266_
+ sky130_fd_sc_hd__o21a_1
X_19720_ clknet_leaf_132_clk _00664_ net1305 vssd1 vssd1 vccd1 vccd1 control.body\[678\]
+ sky130_fd_sc_hd__dfrtp_1
X_16932_ _02602_ _02603_ _02604_ _02605_ vssd1 vssd1 vccd1 vccd1 _02611_ sky130_fd_sc_hd__or4_1
XANTENNA__09492__B net1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12055_ img_gen.tracker.frame\[72\] net628 net610 img_gen.tracker.frame\[75\] _07026_
+ vssd1 vssd1 vccd1 vccd1 _07027_ sky130_fd_sc_hd__a221o_1
XANTENNA__20137__RESET_B net1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11006_ net786 control.body\[1080\] _04254_ net1136 _05978_ vssd1 vssd1 vccd1 vccd1
+ _05979_ sky130_fd_sc_hd__o221a_1
X_19651_ clknet_leaf_133_clk _00595_ net1308 vssd1 vssd1 vccd1 vccd1 control.body\[737\]
+ sky130_fd_sc_hd__dfrtp_1
X_16863_ ag2.body\[207\] net933 vssd1 vssd1 vccd1 vccd1 _02542_ sky130_fd_sc_hd__or2_1
XANTENNA__15445__B1 _01601_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16642__C1 net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18602_ clknet_leaf_17_clk img_gen.tracker.next_frame\[40\] net1320 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[40\] sky130_fd_sc_hd__dfrtp_1
X_15814_ ag2.body\[273\] net205 _01642_ ag2.body\[265\] vssd1 vssd1 vccd1 vccd1 _01059_
+ sky130_fd_sc_hd__a22o_1
X_19582_ clknet_leaf_118_clk net2505 net1388 vssd1 vssd1 vccd1 vccd1 control.body\[812\]
+ sky130_fd_sc_hd__dfrtp_1
X_16794_ obsg2.obstacleArray\[136\] obsg2.obstacleArray\[137\] obsg2.obstacleArray\[138\]
+ obsg2.obstacleArray\[139\] net456 net399 vssd1 vssd1 vccd1 vccd1 _02473_ sky130_fd_sc_hd__mux4_1
X_18533_ clknet_leaf_136_clk _00059_ net1298 vssd1 vssd1 vccd1 vccd1 img_gen.updater.commands.count\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_15745_ ag2.body\[340\] net217 _01634_ ag2.body\[332\] vssd1 vssd1 vccd1 vccd1 _00998_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_99_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12957_ net294 _07673_ _07674_ net1880 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[239\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_90_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18464_ net969 net883 _03951_ vssd1 vssd1 vccd1 vccd1 _03952_ sky130_fd_sc_hd__and3_1
XANTENNA__11482__A1 _06433_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11908_ net1215 net1190 img_gen.tracker.frame\[373\] vssd1 vssd1 vccd1 vccd1 _06880_
+ sky130_fd_sc_hd__or3_1
XFILLER_0_5_1614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19115__CLK clknet_leaf_141_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15676_ ag2.body\[407\] net142 _01626_ ag2.body\[399\] vssd1 vssd1 vccd1 vccd1 _00937_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_87_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12888_ net245 _07643_ _07644_ net1845 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[201\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_34_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17415_ ag2.body\[283\] net721 net699 ag2.body\[286\] vssd1 vssd1 vccd1 vccd1 _03094_
+ sky130_fd_sc_hd__a22o_1
X_14627_ net989 ag2.body\[465\] vssd1 vssd1 vccd1 vccd1 _08788_ sky130_fd_sc_hd__xor2_1
X_18395_ net326 _03791_ vssd1 vssd1 vccd1 vccd1 _03885_ sky130_fd_sc_hd__nand2_1
X_11839_ img_gen.tracker.frame\[494\] net617 net602 img_gen.tracker.frame\[497\] vssd1
+ vssd1 vccd1 vccd1 _06811_ sky130_fd_sc_hd__o22a_1
XANTENNA__14420__A1 net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14420__B2 net1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11234__A1 _04695_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10037__A2 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17346_ net926 _03017_ vssd1 vssd1 vccd1 vccd1 _03025_ sky130_fd_sc_hd__xor2_1
XFILLER_0_86_1603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09948__A net1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14558_ net802 ag2.body\[70\] ag2.body\[71\] net793 _08718_ vssd1 vssd1 vccd1 vccd1
+ _08719_ sky130_fd_sc_hd__a221o_1
XFILLER_0_83_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11785__A2 net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12982__A1 net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13509_ net276 _07914_ _07915_ net1924 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[551\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA_max_cap363_X net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10446__X _05419_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17277_ ag2.body\[556\] net962 vssd1 vssd1 vccd1 vccd1 _02956_ sky130_fd_sc_hd__or2_1
X_14489_ net821 ag2.body\[347\] ag2.body\[351\] net796 _08647_ vssd1 vssd1 vccd1 vccd1
+ _08650_ sky130_fd_sc_hd__a221o_1
XFILLER_0_109_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19016_ clknet_leaf_1_clk img_gen.tracker.next_frame\[454\] net1246 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[454\] sky130_fd_sc_hd__dfrtp_1
X_16228_ _01905_ _01906_ vssd1 vssd1 vccd1 vccd1 _01907_ sky130_fd_sc_hd__nor2_1
XFILLER_0_130_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12734__A1 net237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16159_ obsg2.obstacleArray\[26\] obsg2.obstacleArray\[27\] net428 vssd1 vssd1 vccd1
+ vccd1 _01838_ sky130_fd_sc_hd__mux2_1
XANTENNA__12661__X _07535_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18061__A net42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08981_ ag2.body\[75\] vssd1 vssd1 vccd1 vccd1 _04006_ sky130_fd_sc_hd__inv_2
XANTENNA__15684__B1 _01627_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11718__A net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19918_ clknet_leaf_55_clk _00862_ net1456 vssd1 vssd1 vccd1 vccd1 ag2.body\[476\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__09970__X _04943_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11437__B net1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19849_ clknet_leaf_93_clk _00793_ net1412 vssd1 vssd1 vccd1 vccd1 ag2.body\[551\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_120_1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14239__A1 net841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14239__B2 net799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09602_ net1120 control.body\[636\] vssd1 vssd1 vccd1 vccd1 _04575_ sky130_fd_sc_hd__xor2_1
XFILLER_0_74_1039 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09533_ net1182 control.body\[1026\] vssd1 vssd1 vccd1 vccd1 _04506_ sky130_fd_sc_hd__and2b_1
XFILLER_0_64_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout260_A net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17124__B net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17189__B1 net705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17728__A2 net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09464_ ag2.body\[376\] net784 net1177 _04134_ vssd1 vssd1 vccd1 vccd1 _04437_ sky130_fd_sc_hd__a22o_1
XFILLER_0_38_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09395_ net273 _04345_ _04381_ vssd1 vssd1 vccd1 vccd1 _01405_ sky130_fd_sc_hd__nor3_1
XANTENNA_fanout525_A net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16455__S _02076_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14411__A1 net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14764__A net1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10069__A net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1267_A net1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20624_ sound_gen.dac1.dacCount\[2\] vssd1 vssd1 vccd1 vccd1 net11 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_80_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11599__S net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11776__A2 net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12973__A1 net254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20555_ clknet_leaf_106_clk _01420_ _00029_ vssd1 vssd1 vccd1 vccd1 sound_gen.osc1.stayCount\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09577__B net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout313_X net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1055_X net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1434_A net1435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13099__B _07572_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20486_ clknet_leaf_37_clk _01373_ net1350 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[122\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_131_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_907 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout894_A control.body_update.curr_length\[7\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__12725__A1 net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16190__S net346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17113__B1 net727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1222_X net1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1575 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10736__B1 net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09593__A net1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_3670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10170_ _05134_ _05135_ _05136_ _05138_ vssd1 vssd1 vccd1 vccd1 _05143_ sky130_fd_sc_hd__or4_1
XFILLER_0_125_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_110_3681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout682_X net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_3692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11187__X _06160_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1106 ag2.x\[1\] vssd1 vssd1 vccd1 vccd1 net1106 sky130_fd_sc_hd__buf_4
XANTENNA__10751__A3 _05710_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1117 ag2.x\[1\] vssd1 vssd1 vccd1 vccd1 net1117 sky130_fd_sc_hd__buf_4
Xfanout130 net131 vssd1 vssd1 vccd1 vccd1 net130 sky130_fd_sc_hd__buf_2
XANTENNA__18208__A3 _03703_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10532__A net1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_6_0_clk_X clknet_3_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1128 net1129 vssd1 vssd1 vccd1 vccd1 net1128 sky130_fd_sc_hd__buf_4
Xfanout141 net144 vssd1 vssd1 vccd1 vccd1 net141 sky130_fd_sc_hd__buf_2
Xfanout1139 net1143 vssd1 vssd1 vccd1 vccd1 net1139 sky130_fd_sc_hd__clkbuf_8
XANTENNA__13150__A1 net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout152 net154 vssd1 vssd1 vccd1 vccd1 net152 sky130_fd_sc_hd__buf_2
XANTENNA__11347__B net1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout163 net165 vssd1 vssd1 vccd1 vccd1 net163 sky130_fd_sc_hd__buf_2
Xfanout174 net176 vssd1 vssd1 vccd1 vccd1 net174 sky130_fd_sc_hd__buf_2
Xfanout185 net187 vssd1 vssd1 vccd1 vccd1 net185 sky130_fd_sc_hd__buf_2
XANTENNA__17960__D net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout947_X net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14939__A net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout196 net218 vssd1 vssd1 vccd1 vccd1 net196 sky130_fd_sc_hd__buf_2
XANTENNA__13843__A _04647_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13860_ ag2.body\[23\] net116 _08134_ ag2.body\[15\] vssd1 vssd1 vccd1 vccd1 _00103_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_88_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19138__CLK clknet_leaf_132_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08937__A ag2.goodColl vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout59_X net59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1416 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12811_ net327 _07511_ vssd1 vssd1 vccd1 vccd1 _07607_ sky130_fd_sc_hd__nand2_2
XANTENNA__17034__B net954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13791_ net687 _08097_ _08096_ vssd1 vssd1 vccd1 vccd1 _08098_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_2_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_104_3485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11363__A net1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_3496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15530_ ag2.body\[533\] net157 _01610_ ag2.body\[525\] vssd1 vssd1 vccd1 vccd1 _00807_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_74_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12742_ net284 _07573_ _07574_ net1713 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[125\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__16927__B1 net691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17969__B net45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12178__B _07147_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16873__B net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_69_Right_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19288__CLK clknet_leaf_98_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11082__B net1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12673_ net289 _07540_ _07541_ net1827 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[89\]
+ sky130_fd_sc_hd__a22o_1
X_15461_ _05453_ net63 vssd1 vssd1 vccd1 vccd1 _01603_ sky130_fd_sc_hd__and2_2
XANTENNA__14674__A net1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08943__Y _03968_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17200_ _04058_ net941 net931 _04059_ _02874_ vssd1 vssd1 vccd1 vccd1 _02879_ sky130_fd_sc_hd__a221o_1
XANTENNA__11650__X _06623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14412_ net1008 _03974_ _08570_ _08571_ _08572_ vssd1 vssd1 vccd1 vccd1 _08573_ sky130_fd_sc_hd__a221o_1
X_11624_ obsg2.obstacleArray\[40\] obsg2.obstacleArray\[41\] obsg2.obstacleArray\[44\]
+ obsg2.obstacleArray\[45\] net1123 net510 vssd1 vssd1 vccd1 vccd1 _06597_ sky130_fd_sc_hd__mux4_1
X_18180_ _03619_ _03703_ obsg2.obstacleArray\[87\] vssd1 vssd1 vccd1 vccd1 _03729_
+ sky130_fd_sc_hd__a21oi_1
X_15392_ net2274 net80 _01596_ net2362 vssd1 vssd1 vccd1 vccd1 _00683_ sky130_fd_sc_hd__a22o_1
XANTENNA__18144__A2 _03566_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11767__A2 net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17131_ _02808_ _02809_ vssd1 vssd1 vccd1 vccd1 _02810_ sky130_fd_sc_hd__nand2_1
XANTENNA__17985__A net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16155__A1 obsg2.obstacleArray\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09487__B net1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11555_ _06509_ _06526_ vssd1 vssd1 vccd1 vccd1 _06528_ sky130_fd_sc_hd__xor2_2
XANTENNA__11810__B net597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14343_ net1034 ag2.body\[612\] vssd1 vssd1 vccd1 vccd1 _08504_ sky130_fd_sc_hd__xor2_1
XFILLER_0_135_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_117_3879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20184__Q ag2.body\[214\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10506_ net1087 control.body\[982\] vssd1 vssd1 vccd1 vccd1 _05479_ sky130_fd_sc_hd__xnor2_1
X_17062_ _02739_ _02740_ vssd1 vssd1 vccd1 vccd1 _02741_ sky130_fd_sc_hd__nand2_1
X_14274_ net818 ag2.body\[11\] ag2.body\[12\] net812 _08423_ vssd1 vssd1 vccd1 vccd1
+ _08435_ sky130_fd_sc_hd__a221o_1
XFILLER_0_52_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11486_ _04434_ _04469_ _04902_ _06458_ vssd1 vssd1 vccd1 vccd1 _06459_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_122_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16013_ _01685_ _01691_ vssd1 vssd1 vccd1 vccd1 _01692_ sky130_fd_sc_hd__nor2_1
X_13225_ _06821_ _07633_ vssd1 vssd1 vccd1 vccd1 _07802_ sky130_fd_sc_hd__and2_1
XFILLER_0_46_1642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10437_ net1083 control.body\[934\] vssd1 vssd1 vccd1 vccd1 _05410_ sky130_fd_sc_hd__and2_1
XFILLER_0_46_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_78_Right_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13156_ net277 _07767_ _07768_ net1931 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[344\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__20561__D toggle1.nextDisplayOut\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10368_ net1077 control.body\[766\] vssd1 vssd1 vccd1 vccd1 _05341_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_42_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10713__Y _05686_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17209__B net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12641__B _07523_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12107_ img_gen.tracker.frame\[168\] net627 net593 img_gen.tracker.frame\[177\] vssd1
+ vssd1 vccd1 vccd1 _07079_ sky130_fd_sc_hd__a22o_1
X_17964_ net518 _03588_ vssd1 vssd1 vccd1 vccd1 _01262_ sky130_fd_sc_hd__nor2_1
X_13087_ net290 _07734_ _07735_ net1805 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[308\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__10442__A _04586_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10299_ _05177_ _05206_ _05236_ _05271_ vssd1 vssd1 vccd1 vccd1 _05272_ sky130_fd_sc_hd__and4_1
XFILLER_0_97_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19703_ clknet_leaf_135_clk _00647_ net1301 vssd1 vssd1 vccd1 vccd1 control.body\[693\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12038_ net576 _07009_ vssd1 vssd1 vccd1 vccd1 _07010_ sky130_fd_sc_hd__nor2_1
X_16915_ ag2.body\[560\] net881 vssd1 vssd1 vccd1 vccd1 _02594_ sky130_fd_sc_hd__or2_1
XANTENNA__10161__B net1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17895_ net2175 _03531_ _03532_ _03521_ vssd1 vssd1 vccd1 vccd1 _01249_ sky130_fd_sc_hd__a22o_1
X_19634_ clknet_leaf_123_clk _00578_ net1406 vssd1 vssd1 vccd1 vccd1 control.body\[752\]
+ sky130_fd_sc_hd__dfrtp_1
X_16846_ ag2.body\[171\] net717 net704 ag2.body\[173\] _02524_ vssd1 vssd1 vccd1 vccd1
+ _02525_ sky130_fd_sc_hd__a221o_1
XANTENNA__09950__B net1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16091__B1 net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19565_ clknet_leaf_116_clk net2532 net1387 vssd1 vssd1 vccd1 vccd1 control.body\[827\]
+ sky130_fd_sc_hd__dfrtp_1
X_16777_ obsg2.obstacleArray\[24\] net493 net485 obsg2.obstacleArray\[25\] vssd1 vssd1
+ vccd1 vccd1 _02456_ sky130_fd_sc_hd__a22o_1
XFILLER_0_92_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13989_ ag2.body\[126\] net211 _08159_ ag2.body\[118\] vssd1 vssd1 vccd1 vccd1 _00207_
+ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_87_Right_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18516_ net1512 net1506 vssd1 vssd1 vccd1 vccd1 _00047_ sky130_fd_sc_hd__or2_1
X_15728_ ag2.body\[357\] net194 _01632_ ag2.body\[349\] vssd1 vssd1 vccd1 vccd1 _00983_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_73_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19496_ clknet_leaf_113_clk _00440_ net1399 vssd1 vssd1 vccd1 vccd1 control.body\[902\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_1646 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16918__B1 net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18447_ _05075_ _06173_ _03828_ vssd1 vssd1 vccd1 vccd1 _03936_ sky130_fd_sc_hd__o21ai_1
X_15659_ _06111_ net57 vssd1 vssd1 vccd1 vccd1 _01625_ sky130_fd_sc_hd__nor2_2
XFILLER_0_5_1444 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17591__B1 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_1370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18655__CLK clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09180_ ag2.body\[559\] vssd1 vssd1 vccd1 vccd1 _04205_ sky130_fd_sc_hd__inv_2
X_18378_ net2246 _08024_ _03866_ net464 _03868_ vssd1 vssd1 vccd1 vccd1 _01396_ sky130_fd_sc_hd__o221a_1
XFILLER_0_44_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17329_ net1043 net870 vssd1 vssd1 vccd1 vccd1 _03008_ sky130_fd_sc_hd__xor2_1
XFILLER_0_83_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_701 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_133_4371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_1444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_133_4382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09820__B2 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_133_4393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16697__A2 net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20340_ clknet_leaf_140_clk _01231_ net1292 vssd1 vssd1 vccd1 vccd1 img_gen.updater.commands.rR1.rainbowRNG\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_12_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17894__B2 _03523_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10336__B net1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_96_Right_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13928__A _04863_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20271_ clknet_leaf_38_clk net5 net1353 vssd1 vssd1 vccd1 vccd1 control.button4.Q\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10718__B1 net766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout106_A net107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13380__A1 net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09584__B1 _04553_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17119__B net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11448__A net1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08964_ ag2.body\[43\] vssd1 vssd1 vccd1 vccd1 _03989_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout1015_A net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_1993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_4186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16958__B net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_4197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_51_1868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09887__A1 net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13663__A net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09860__B net1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10497__A2 net1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_3_Left_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_32_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13382__B net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09639__A1 net1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19430__CLK clknet_leaf_111_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout263_X net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09639__B2 net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14632__B2 net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09516_ net1201 control.body\[833\] vssd1 vssd1 vccd1 vccd1 _04489_ sky130_fd_sc_hd__xor2_1
XFILLER_0_67_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_1292 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16693__B net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19924__RESET_B net1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09447_ net917 net921 vssd1 vssd1 vccd1 vccd1 _04420_ sky130_fd_sc_hd__nand2_4
XANTENNA__11997__A2 net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout430_X net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16185__S net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14494__A net1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1172_X net1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout528_X net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17582__B1 net878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout907_A net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09588__A net1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09378_ sound_gen.osc1.stayCount\[15\] _04366_ _04359_ net271 vssd1 vssd1 vccd1 vccd1
+ _01414_ sky130_fd_sc_hd__o211a_1
XANTENNA__19580__CLK clknet_leaf_118_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20607_ net1539 vssd1 vssd1 vccd1 vccd1 gpio_oeb[19] sky130_fd_sc_hd__buf_2
XANTENNA__11630__B net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16137__A1 net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15102__B net58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10527__A net1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_10_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_49_Left_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11340_ _06290_ _06300_ _06312_ _05856_ vssd1 vssd1 vccd1 vccd1 _06313_ sky130_fd_sc_hd__o22a_1
XANTENNA__20482__RESET_B net1356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20538_ clknet_leaf_107_clk _01403_ _00012_ vssd1 vssd1 vccd1 vccd1 sound_gen.osc1.stayCount\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__17885__A1 net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14699__A1 net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_3732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10246__B net1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14699__B2 net1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_3743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_112_3754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11271_ ag2.body\[125\] net1116 vssd1 vssd1 vccd1 vccd1 _06244_ sky130_fd_sc_hd__xor2_1
XANTENNA__20411__RESET_B net1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20469_ clknet_leaf_34_clk _01356_ net1346 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[105\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_127_1275 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16214__A net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13010_ net240 _07699_ _07700_ net2017 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[267\]
+ sky130_fd_sc_hd__a22o_1
X_10222_ ag2.body\[567\] net1052 vssd1 vssd1 vccd1 vccd1 _05195_ sky130_fd_sc_hd__nand2_1
XFILLER_0_123_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_759 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1274 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15648__B1 _01623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10153_ ag2.body\[59\] net1155 vssd1 vssd1 vccd1 vccd1 _05126_ sky130_fd_sc_hd__nand2_1
XANTENNA__17971__C net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16868__B net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16860__A2 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_115_clk_X clknet_leaf_115_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10084_ _05053_ _05054_ _05055_ _05056_ vssd1 vssd1 vccd1 vccd1 _05057_ sky130_fd_sc_hd__a22o_1
X_14961_ control.body\[1035\] net172 _01547_ control.body\[1027\] vssd1 vssd1 vccd1
+ vccd1 _00301_ sky130_fd_sc_hd__a22o_1
Xhold8 img_gen.control.button5.Q\[0\] vssd1 vssd1 vccd1 vccd1 net1570 sky130_fd_sc_hd__dlygate4sd3_1
X_16700_ obsg2.obstacleArray\[83\] net502 net494 obsg2.obstacleArray\[80\] vssd1 vssd1
+ vccd1 vccd1 _02379_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_58_Left_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13912_ ag2.body\[57\] net120 _08151_ ag2.body\[49\] vssd1 vssd1 vccd1 vccd1 _00138_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__09770__B net1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_3547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17680_ ag2.body\[477\] net705 net688 ag2.body\[479\] vssd1 vssd1 vccd1 vccd1 _03359_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__10488__A2 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_3558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14892_ net2582 net180 _01539_ net2325 vssd1 vssd1 vccd1 vccd1 _00240_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_106_3569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16631_ obsg2.obstacleArray\[63\] net450 net391 _02309_ vssd1 vssd1 vccd1 vccd1 _02310_
+ sky130_fd_sc_hd__o211a_1
X_13843_ _04647_ net56 vssd1 vssd1 vccd1 vccd1 _08133_ sky130_fd_sc_hd__nor2_2
XANTENNA__12189__A net1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_1089 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19350_ clknet_leaf_102_clk _00294_ net1429 vssd1 vssd1 vccd1 vccd1 control.body\[1044\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__20179__Q ag2.body\[209\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16562_ _02226_ net358 _02232_ _02240_ vssd1 vssd1 vccd1 vccd1 _02241_ sky130_fd_sc_hd__a31o_1
XFILLER_0_74_1381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13774_ img_gen.updater.commands.count\[8\] img_gen.updater.commands.count\[9\] _08082_
+ vssd1 vssd1 vccd1 vccd1 _08086_ sky130_fd_sc_hd__and3_1
X_10986_ net1172 control.body\[754\] vssd1 vssd1 vccd1 vccd1 _05959_ sky130_fd_sc_hd__xor2_1
XFILLER_0_85_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_84_2890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19923__CLK clknet_leaf_51_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18301_ _03792_ _03796_ vssd1 vssd1 vccd1 vccd1 _03797_ sky130_fd_sc_hd__nand2_1
X_15513_ ag2.body\[550\] net155 _01608_ ag2.body\[542\] vssd1 vssd1 vccd1 vccd1 _00792_
+ sky130_fd_sc_hd__a22o_1
X_12725_ net285 _07565_ _07566_ net1682 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[116\]
+ sky130_fd_sc_hd__a22o_1
X_19281_ clknet_leaf_97_clk net2144 net1451 vssd1 vssd1 vccd1 vccd1 control.body\[1119\]
+ sky130_fd_sc_hd__dfrtp_1
X_16493_ net402 _02171_ vssd1 vssd1 vccd1 vccd1 _02172_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_80_2754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17573__B1 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_2765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_80_2776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18232_ _03673_ net41 vssd1 vssd1 vccd1 vccd1 _03755_ sky130_fd_sc_hd__nor2_1
XANTENNA__14835__C _01504_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15444_ ag2.body\[600\] net86 _01601_ ag2.body\[592\] vssd1 vssd1 vccd1 vccd1 _00730_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_61_2175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12656_ net307 _07532_ vssd1 vssd1 vccd1 vccd1 _07533_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_61_2186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_2197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16108__B net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12937__A1 net246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11607_ obsg2.obstacleArray\[26\] net633 net509 obsg2.obstacleArray\[30\] net760
+ vssd1 vssd1 vccd1 vccd1 _06580_ sky130_fd_sc_hd__o221a_1
X_18163_ obsg2.obstacleArray\[78\] _03720_ net522 vssd1 vssd1 vccd1 vccd1 _01329_
+ sky130_fd_sc_hd__o21a_1
X_12587_ net327 _07493_ vssd1 vssd1 vccd1 vccd1 _07494_ sky130_fd_sc_hd__or2_2
XFILLER_0_5_729 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15375_ control.body\[666\] net69 _01594_ net2255 vssd1 vssd1 vccd1 vccd1 _00668_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__10948__B1 net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10437__A net1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_440 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09785__X _04758_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17114_ ag2.body\[542\] net942 vssd1 vssd1 vccd1 vccd1 _02793_ sky130_fd_sc_hd__xor2_1
XFILLER_0_68_1152 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14326_ net842 ag2.body\[448\] ag2.body\[454\] net800 _08486_ vssd1 vssd1 vccd1 vccd1
+ _08487_ sky130_fd_sc_hd__o221a_1
XFILLER_0_135_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18094_ net519 _03678_ vssd1 vssd1 vccd1 vccd1 _01302_ sky130_fd_sc_hd__nor2_1
XFILLER_0_111_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11538_ _06509_ _06510_ vssd1 vssd1 vccd1 vccd1 _06511_ sky130_fd_sc_hd__nand2_2
XFILLER_0_29_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10156__B net1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_2694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold408 img_gen.tracker.frame\[277\] vssd1 vssd1 vccd1 vccd1 net1970 sky130_fd_sc_hd__dlygate4sd3_1
X_17045_ ag2.body\[262\] net943 vssd1 vssd1 vccd1 vccd1 _02724_ sky130_fd_sc_hd__xor2_1
Xhold419 toggle1.bcd_tens\[1\] vssd1 vssd1 vccd1 vccd1 net1981 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__20152__RESET_B net1452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14257_ net815 ag2.body\[76\] ag2.body\[78\] net802 _08416_ vssd1 vssd1 vccd1 vccd1
+ _08418_ sky130_fd_sc_hd__a221o_1
XFILLER_0_106_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11469_ ag2.body\[490\] net1184 vssd1 vssd1 vccd1 vccd1 _06442_ sky130_fd_sc_hd__xor2_1
XFILLER_0_111_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_74_2569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09566__B1 net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13208_ _07624_ _07639_ vssd1 vssd1 vccd1 vccd1 _07794_ sky130_fd_sc_hd__nor2_1
XFILLER_0_0_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14188_ net999 ag2.body\[160\] vssd1 vssd1 vccd1 vccd1 _08349_ sky130_fd_sc_hd__nand2_1
XANTENNA__19208__Q ag2.body\[71\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12371__B net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11912__A2 net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16300__A1 _01912_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15103__A2 net183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13139_ net291 _07758_ _07759_ net1725 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[335\]
+ sky130_fd_sc_hd__a22o_1
X_18996_ clknet_leaf_0_clk img_gen.tracker.next_frame\[434\] net1244 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[434\] sky130_fd_sc_hd__dfrtp_1
X_17947_ net318 _03575_ obsg2.obstacleArray\[7\] vssd1 vssd1 vccd1 vccd1 _03576_ sky130_fd_sc_hd__a21oi_1
XANTENNA__19453__CLK clknet_leaf_111_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1470 net1478 vssd1 vssd1 vccd1 vccd1 net1470 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_75_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1481 net1482 vssd1 vssd1 vccd1 vccd1 net1481 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_20_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17878_ _04903_ _03458_ _04688_ vssd1 vssd1 vccd1 vccd1 _03518_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_122_4050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1492 net1493 vssd1 vssd1 vccd1 vccd1 net1492 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_75_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16829_ ag2.body\[228\] net711 net699 ag2.body\[230\] _02502_ vssd1 vssd1 vccd1 vccd1
+ _02508_ sky130_fd_sc_hd__a221o_1
X_19617_ clknet_leaf_120_clk _00561_ net1392 vssd1 vssd1 vccd1 vccd1 control.body\[783\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15811__B1 _01641_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19548_ clknet_leaf_115_clk _00492_ net1396 vssd1 vssd1 vccd1 vccd1 control.body\[842\]
+ sky130_fd_sc_hd__dfrtp_1
X_09301_ sound_gen.osc1.count\[2\] sound_gen.osc1.count\[1\] sound_gen.osc1.count\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04321_ sky130_fd_sc_hd__and3_1
XANTENNA__16367__A1 net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_757 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19479_ clknet_leaf_111_clk _00423_ net1424 vssd1 vssd1 vccd1 vccd1 control.body\[917\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17402__B net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_135_4433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09232_ control.body\[1101\] vssd1 vssd1 vccd1 vccd1 _04257_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_135_4444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_4455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_44_1661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_4308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12546__B net436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12928__A1 net290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_131_4319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09163_ ag2.body\[513\] vssd1 vssd1 vccd1 vccd1 _04188_ sky130_fd_sc_hd__inv_2
XFILLER_0_133_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_20_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09094_ ag2.body\[337\] vssd1 vssd1 vccd1 vccd1 _04119_ sky130_fd_sc_hd__inv_2
XFILLER_0_114_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20323_ clknet_leaf_46_clk _01219_ net1379 vssd1 vssd1 vccd1 vccd1 ag2.body\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold920 control.body\[738\] vssd1 vssd1 vccd1 vccd1 net2482 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_128_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16034__A net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_540 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1132_A net1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold931 control.body\[662\] vssd1 vssd1 vccd1 vccd1 net2493 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_90_3061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold942 control.body\[804\] vssd1 vssd1 vccd1 vccd1 net2504 sky130_fd_sc_hd__dlygate4sd3_1
X_20254_ clknet_leaf_70_clk _01198_ net1497 vssd1 vssd1 vccd1 vccd1 ag2.body\[140\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_90_3072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold953 control.body\[875\] vssd1 vssd1 vccd1 vccd1 net2515 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13377__B net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_129_4248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_3083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold964 control.body\[642\] vssd1 vssd1 vccd1 vccd1 net2526 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_129_4259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold975 control.body\[1012\] vssd1 vssd1 vccd1 vccd1 net2537 sky130_fd_sc_hd__dlygate4sd3_1
Xhold986 control.body\[707\] vssd1 vssd1 vccd1 vccd1 net2548 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold997 control.body\[692\] vssd1 vssd1 vccd1 vccd1 net2559 sky130_fd_sc_hd__dlygate4sd3_1
X_20185_ clknet_leaf_87_clk _01129_ net1460 vssd1 vssd1 vccd1 vccd1 ag2.body\[215\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_38_1487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09996_ net1096 control.body\[733\] vssd1 vssd1 vccd1 vccd1 _04969_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout1018_X net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08947_ net1016 vssd1 vssd1 vccd1 vccd1 _03972_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout380_X net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_4_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13393__A net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_84_clk_A clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10810__A net1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_1392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_1256 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_3400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_3411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10840_ _04632_ _05076_ vssd1 vssd1 vccd1 vccd1 _05813_ sky130_fd_sc_hd__nor2_2
XFILLER_0_94_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_99_clk_A clknet_4_11__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13840__B net223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17312__B net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12092__A1 net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10771_ ag2.body\[221\] net1114 vssd1 vssd1 vccd1 vccd1 _05744_ sky130_fd_sc_hd__xor2_1
XANTENNA__17555__B1 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout812_X net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_145_clk clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_145_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_109_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_142_clk_A clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12510_ img_gen.tracker.frame\[17\] net649 _07450_ vssd1 vssd1 vccd1 vccd1 _07451_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_48_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16453__S1 net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13490_ net328 _07505_ _07813_ vssd1 vssd1 vccd1 vccd1 _07908_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_118_3930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12441_ net748 net1045 _06630_ _07401_ vssd1 vssd1 vccd1 vccd1 _07402_ sky130_fd_sc_hd__o211a_1
XFILLER_0_129_1304 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_22_clk_A clknet_4_6__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_114_3805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_259 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19326__CLK clknet_leaf_103_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_985 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12372_ net263 net241 net289 _07320_ vssd1 vssd1 vccd1 vccd1 _07338_ sky130_fd_sc_hd__o31a_1
X_15160_ net2509 net105 _01569_ control.body\[852\] vssd1 vssd1 vccd1 vccd1 _00478_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_34_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15767__B _01631_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11323_ ag2.body\[552\] net1228 vssd1 vssd1 vccd1 vccd1 _06296_ sky130_fd_sc_hd__xor2_1
X_14111_ net1035 ag2.body\[572\] vssd1 vssd1 vccd1 vccd1 _08272_ sky130_fd_sc_hd__or2_1
XFILLER_0_133_884 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15091_ net2306 net147 _01562_ control.body\[918\] vssd1 vssd1 vccd1 vccd1 _00416_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__20303__CLK clknet_leaf_37_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_37_clk_A clknet_4_5__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14042_ net1039 _04181_ _04183_ net1011 _08195_ vssd1 vssd1 vccd1 vccd1 _08203_ sky130_fd_sc_hd__a221o_1
X_11254_ net1151 control.body\[771\] vssd1 vssd1 vccd1 vccd1 _06227_ sky130_fd_sc_hd__nand2_1
XANTENNA__17982__B _03539_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10158__A1 ag2.body\[60\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10158__B2 ag2.body\[63\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10704__B net1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10205_ net742 _04599_ net637 vssd1 vssd1 vccd1 vccd1 _05178_ sky130_fd_sc_hd__a21o_1
XFILLER_0_120_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18850_ clknet_leaf_16_clk img_gen.tracker.next_frame\[288\] net1321 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[288\] sky130_fd_sc_hd__dfrtp_1
X_11185_ ag2.body\[176\] net784 net782 ag2.body\[177\] vssd1 vssd1 vccd1 vccd1 _06158_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_66_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_3609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_66_Left_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17801_ _03288_ net940 net948 net969 vssd1 vssd1 vccd1 vccd1 _03472_ sky130_fd_sc_hd__and4b_1
XANTENNA__09781__A net1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10136_ _05105_ _05106_ _05107_ _05108_ _05104_ vssd1 vssd1 vccd1 vccd1 _05109_ sky130_fd_sc_hd__a221o_1
X_18781_ clknet_leaf_12_clk img_gen.tracker.next_frame\[219\] net1284 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[219\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_1107 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15993_ ag2.body\[3\] _01660_ _01661_ _01675_ vssd1 vssd1 vccd1 vccd1 _01205_ sky130_fd_sc_hd__a22o_1
XANTENNA__14844__A1 _08705_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17732_ _03256_ _03262_ _03355_ vssd1 vssd1 vccd1 vccd1 _03411_ sky130_fd_sc_hd__o21a_1
X_10067_ net1148 control.body\[715\] vssd1 vssd1 vccd1 vccd1 _05040_ sky130_fd_sc_hd__xor2_1
X_14944_ control.body\[1052\] net168 _01545_ control.body\[1044\] vssd1 vssd1 vccd1
+ vccd1 _00286_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_86_2941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17663_ _03337_ _03338_ _03341_ vssd1 vssd1 vccd1 vccd1 _03342_ sky130_fd_sc_hd__a21o_1
XANTENNA__10330__A1 control.body_update.curr_length\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14875_ net2143 net182 _01537_ control.body\[1111\] vssd1 vssd1 vccd1 vccd1 _00225_
+ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_4_5__f_clk_A clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_82_2816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19402_ clknet_leaf_103_clk _00346_ net1427 vssd1 vssd1 vccd1 vccd1 control.body\[984\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkload1_A clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_2362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16614_ obsg2.obstacleArray\[42\] net442 vssd1 vssd1 vccd1 vccd1 _02293_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_82_2827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_2373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13826_ _04270_ _08118_ _08122_ _08117_ vssd1 vssd1 vccd1 vccd1 _08123_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_82_2838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17594_ _03267_ _03272_ vssd1 vssd1 vccd1 vccd1 _03273_ sky130_fd_sc_hd__nand2_1
XFILLER_0_15_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_2237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19333_ clknet_leaf_100_clk _00277_ net1443 vssd1 vssd1 vccd1 vccd1 control.body\[1059\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_63_2248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16545_ obsg2.obstacleArray\[96\] net441 vssd1 vssd1 vccd1 vccd1 _02224_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_63_2259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_136_clk clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_136_clk
+ sky130_fd_sc_hd__clkbuf_8
X_13757_ img_gen.updater.commands.count\[3\] _08068_ img_gen.updater.commands.count\[4\]
+ vssd1 vssd1 vccd1 vccd1 _08074_ sky130_fd_sc_hd__a21o_1
XFILLER_0_35_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16349__B2 _01912_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10969_ net1205 control.body\[1001\] vssd1 vssd1 vccd1 vccd1 _05942_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_35_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_75_Left_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11551__A net1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19264_ clknet_leaf_74_clk _00208_ net1504 vssd1 vssd1 vccd1 vccd1 ag2.body\[127\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__17010__A2 net712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12708_ net333 _07442_ vssd1 vssd1 vccd1 vccd1 _07558_ sky130_fd_sc_hd__or2_2
X_16476_ obsg2.obstacleArray\[40\] obsg2.obstacleArray\[41\] net453 vssd1 vssd1 vccd1
+ vccd1 _02155_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13688_ _04945_ _08029_ vssd1 vssd1 vccd1 vccd1 _08031_ sky130_fd_sc_hd__nand2_2
XFILLER_0_127_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18215_ obsg2.obstacleArray\[104\] _03746_ net528 vssd1 vssd1 vccd1 vccd1 _01355_
+ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_14_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_1447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11270__B net1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15427_ ag2.body\[617\] net84 _01599_ ag2.body\[609\] vssd1 vssd1 vccd1 vccd1 _00715_
+ sky130_fd_sc_hd__a22o_1
X_19195_ clknet_leaf_53_clk _00139_ net1455 vssd1 vssd1 vccd1 vccd1 ag2.body\[58\]
+ sky130_fd_sc_hd__dfrtp_4
X_12639_ net604 net435 net467 net574 vssd1 vssd1 vccd1 vccd1 _07522_ sky130_fd_sc_hd__or4_1
XANTENNA__14862__A _01526_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15572__A2 net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18146_ net47 _03570_ _03704_ obsg2.obstacleArray\[70\] vssd1 vssd1 vccd1 vccd1 _03712_
+ sky130_fd_sc_hd__a31o_1
X_15358_ control.body\[683\] net75 _01592_ net2379 vssd1 vssd1 vccd1 vccd1 _00653_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_31_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15677__B net58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11594__B1 net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10936__A3 _05074_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14309_ net1007 ag2.body\[55\] vssd1 vssd1 vccd1 vccd1 _08470_ sky130_fd_sc_hd__or2_1
Xhold205 img_gen.tracker.frame\[178\] vssd1 vssd1 vccd1 vccd1 net1767 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09675__B net1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18077_ obsg2.obstacleArray\[45\] _03667_ net520 vssd1 vssd1 vccd1 vccd1 _01296_
+ sky130_fd_sc_hd__o21a_1
XANTENNA__19819__CLK clknet_leaf_124_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15289_ net2452 net88 _01584_ control.body\[742\] vssd1 vssd1 vccd1 vccd1 _00592_
+ sky130_fd_sc_hd__a22o_1
Xhold216 img_gen.tracker.frame\[495\] vssd1 vssd1 vccd1 vccd1 net1778 sky130_fd_sc_hd__dlygate4sd3_1
Xhold227 img_gen.tracker.frame\[540\] vssd1 vssd1 vccd1 vccd1 net1789 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13335__A1 net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold238 img_gen.tracker.frame\[478\] vssd1 vssd1 vccd1 vccd1 net1800 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12138__A2 net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17028_ ag2.body\[400\] net888 vssd1 vssd1 vccd1 vccd1 _02707_ sky130_fd_sc_hd__xor2_1
Xhold249 img_gen.tracker.frame\[442\] vssd1 vssd1 vccd1 vccd1 net1811 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_84_Left_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18274__A1 net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12532__D net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout707 net708 vssd1 vssd1 vccd1 vccd1 net707 sky130_fd_sc_hd__clkbuf_4
X_09850_ net779 control.body\[969\] _04250_ net1110 vssd1 vssd1 vccd1 vccd1 _04823_
+ sky130_fd_sc_hd__a22o_1
Xfanout718 _04265_ vssd1 vssd1 vccd1 vccd1 net718 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_124_4101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout729 _04264_ vssd1 vssd1 vccd1 vccd1 net729 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_42_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18843__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_4112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09691__A ag2.body\[68\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09781_ net1087 control.body\[950\] vssd1 vssd1 vccd1 vccd1 _04754_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_33_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18979_ clknet_leaf_8_clk img_gen.tracker.next_frame\[417\] net1265 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[417\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__10630__A net1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19587__RESET_B net1386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18993__CLK clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_137_4506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18329__A2 _04519_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_93_Left_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_46_1723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_138_Right_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_46_1734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_127_clk clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_127_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__17132__B net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16029__A net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1082_A ag2.x\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout438_A net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17001__A2 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_1303 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17071__A2_N net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11821__A1 net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09215_ control.body\[729\] vssd1 vssd1 vccd1 vccd1 _04240_ sky130_fd_sc_hd__inv_2
XFILLER_0_17_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout605_A net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout226_X net226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09146_ ag2.body\[478\] vssd1 vssd1 vccd1 vccd1 _04171_ sky130_fd_sc_hd__inv_2
XANTENNA__09778__B1 net1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_3123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_92_3134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_933 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19499__CLK clknet_leaf_113_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_873 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13388__A net670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09077_ ag2.body\[311\] vssd1 vssd1 vccd1 vccd1 _04102_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1514_A net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1135_X net1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12129__A2 net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20306_ clknet_leaf_70_clk net7 net1497 vssd1 vssd1 vccd1 vccd1 obsmode.sOBSMODE.sync
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_31_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_556 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold750 control.body\[960\] vssd1 vssd1 vccd1 vccd1 net2312 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout974_A ag2.randCord\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout595_X net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold761 control.body\[1086\] vssd1 vssd1 vccd1 vccd1 net2323 sky130_fd_sc_hd__dlygate4sd3_1
Xhold772 control.body\[901\] vssd1 vssd1 vccd1 vccd1 net2334 sky130_fd_sc_hd__dlygate4sd3_1
X_20237_ clknet_leaf_69_clk _01181_ net1496 vssd1 vssd1 vccd1 vccd1 ag2.body\[155\]
+ sky130_fd_sc_hd__dfrtp_4
Xhold783 control.body\[823\] vssd1 vssd1 vccd1 vccd1 net2345 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold794 control.body\[646\] vssd1 vssd1 vccd1 vccd1 net2356 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_1375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17307__B net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20168_ clknet_leaf_81_clk _01112_ net1480 vssd1 vssd1 vccd1 vccd1 ag2.body\[230\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA_fanout762_X net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09979_ net1062 control.body\[1119\] vssd1 vssd1 vccd1 vccd1 _04952_ sky130_fd_sc_hd__xnor2_1
XANTENNA__14826__A1 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16211__B net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18280__A4 _03579_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14826__B2 net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14012__A net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20099_ clknet_leaf_79_clk _01043_ net1486 vssd1 vssd1 vccd1 vccd1 ag2.body\[289\]
+ sky130_fd_sc_hd__dfrtp_4
X_12990_ net278 _07688_ _07689_ net1871 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[257\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_99_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11941_ img_gen.tracker.frame\[157\] net621 net548 img_gen.tracker.frame\[163\] _06912_
+ vssd1 vssd1 vccd1 vccd1 _06913_ sky130_fd_sc_hd__o221a_1
XFILLER_0_118_1049 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14660_ net1021 ag2.body\[526\] vssd1 vssd1 vccd1 vccd1 _08821_ sky130_fd_sc_hd__nand2_1
XANTENNA__17240__A2 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout41_X net41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11872_ net563 _06838_ _06840_ _06843_ vssd1 vssd1 vccd1 vccd1 _06844_ sky130_fd_sc_hd__a31o_1
XFILLER_0_135_1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08945__A net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13611_ control.divider.count\[2\] control.divider.count\[1\] control.divider.count\[0\]
+ control.divider.count\[3\] vssd1 vssd1 vccd1 vccd1 _07983_ sky130_fd_sc_hd__a31o_1
XFILLER_0_95_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_95_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12065__A1 net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10823_ net1112 _04255_ net635 _05794_ _05795_ vssd1 vssd1 vccd1 vccd1 _05796_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_138_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14591_ _08747_ _08749_ _08750_ _08751_ vssd1 vssd1 vccd1 vccd1 _08752_ sky130_fd_sc_hd__or4b_1
XPHY_EDGE_ROW_105_Right_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_118_clk clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_118_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_32_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12467__A net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16330_ obsg2.obstacleArray\[78\] obsg2.obstacleArray\[79\] net406 vssd1 vssd1 vccd1
+ vccd1 _02009_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13542_ net226 _07927_ vssd1 vssd1 vccd1 vccd1 _07928_ sky130_fd_sc_hd__nor2_1
XFILLER_0_137_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10754_ net785 control.body\[888\] _04247_ net1107 _05726_ vssd1 vssd1 vccd1 vccd1
+ _05727_ sky130_fd_sc_hd__a221o_1
XFILLER_0_32_1357 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09481__A2 net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16881__B net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16261_ obsg2.obstacleArray\[52\] obsg2.obstacleArray\[53\] net407 vssd1 vssd1 vccd1
+ vccd1 _01940_ sky130_fd_sc_hd__mux2_1
XANTENNA__18716__CLK clknet_leaf_144_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10685_ ag2.body\[150\] net1088 vssd1 vssd1 vccd1 vccd1 _05658_ sky130_fd_sc_hd__nand2_1
XFILLER_0_109_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13473_ net250 _07900_ _07901_ net1974 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[529\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__14682__A net1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18000_ net45 _03614_ vssd1 vssd1 vccd1 vccd1 _03615_ sky130_fd_sc_hd__nor2_1
XFILLER_0_63_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15212_ control.body\[810\] net93 _01575_ net2472 vssd1 vssd1 vccd1 vccd1 _00524_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_36_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12424_ _07355_ _07383_ _07385_ _07299_ vssd1 vssd1 vccd1 vccd1 _07386_ sky130_fd_sc_hd__a2bb2o_1
X_16192_ obsg2.obstacleArray\[44\] obsg2.obstacleArray\[45\] net421 vssd1 vssd1 vccd1
+ vccd1 _01871_ sky130_fd_sc_hd__mux2_1
XANTENNA__15497__B net54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_75_2620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14299__A1_N net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15143_ control.body\[877\] net105 _01567_ control.body\[869\] vssd1 vssd1 vccd1
+ vccd1 _00463_ sky130_fd_sc_hd__a22o_1
XANTENNA__13298__A _07480_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12355_ net628 _06506_ vssd1 vssd1 vccd1 vccd1 _07322_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_56_2030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_988 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_56_2041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11591__A3 obsg2.obstacleArray\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11306_ ag2.body\[274\] net1187 vssd1 vssd1 vccd1 vccd1 _06279_ sky130_fd_sc_hd__xor2_1
X_19951_ clknet_leaf_45_clk _00895_ net1382 vssd1 vssd1 vccd1 vccd1 ag2.body\[445\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_121_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12286_ _07255_ vssd1 vssd1 vccd1 vccd1 _07256_ sky130_fd_sc_hd__inv_2
X_15074_ control.body\[943\] net149 _01560_ net2561 vssd1 vssd1 vccd1 vccd1 _00401_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_107_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17059__A2 net877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14025_ net996 ag2.body\[24\] vssd1 vssd1 vccd1 vccd1 _08186_ sky130_fd_sc_hd__xor2_1
X_18902_ clknet_leaf_145_clk img_gen.tracker.next_frame\[340\] net1251 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[340\] sky130_fd_sc_hd__dfrtp_1
X_11237_ ag2.body\[194\] net1177 vssd1 vssd1 vccd1 vccd1 _06210_ sky130_fd_sc_hd__nand2_1
X_19882_ clknet_leaf_83_clk _00826_ net1480 vssd1 vssd1 vccd1 vccd1 ag2.body\[504\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_120_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09941__B1 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11168_ net1049 control.body\[783\] vssd1 vssd1 vccd1 vccd1 _06141_ sky130_fd_sc_hd__nand2_1
X_18833_ clknet_leaf_4_clk img_gen.tracker.next_frame\[271\] net1262 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[271\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_120_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14817__A1 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_2413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10119_ net1098 control.body\[709\] vssd1 vssd1 vccd1 vccd1 _05092_ sky130_fd_sc_hd__nand2_1
X_18764_ clknet_leaf_16_clk img_gen.tracker.next_frame\[202\] net1314 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[202\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_69_2424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11099_ ag2.body\[431\] net1056 vssd1 vssd1 vccd1 vccd1 _06072_ sky130_fd_sc_hd__xor2_1
X_15976_ _08118_ net56 vssd1 vssd1 vccd1 vccd1 _01662_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_69_2435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17715_ obsg2.obstacleArray\[136\] obsg2.obstacleArray\[137\] net427 vssd1 vssd1
+ vccd1 vccd1 _03394_ sky130_fd_sc_hd__mux2_1
XFILLER_0_91_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14927_ net2605 net170 _01543_ control.body\[1061\] vssd1 vssd1 vccd1 vccd1 _00271_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_37_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18695_ clknet_leaf_11_clk img_gen.tracker.next_frame\[133\] net1281 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[133\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__17767__B1 _03187_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17231__A2 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17646_ ag2.body\[34\] net858 vssd1 vssd1 vccd1 vccd1 _03325_ sky130_fd_sc_hd__xnor2_1
X_14858_ _08417_ _08422_ _08413_ vssd1 vssd1 vccd1 vccd1 _01529_ sky130_fd_sc_hd__o21a_1
XANTENNA__10854__A2 _04758_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_1414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12648__Y _07528_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17782__A3 net825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13809_ control.divider.detect.Q\[1\] control.divider.detect.Q\[0\] vssd1 vssd1 vccd1
+ vccd1 _08109_ sky130_fd_sc_hd__and2b_1
X_17577_ _03254_ _03255_ _03253_ vssd1 vssd1 vccd1 vccd1 _03256_ sky130_fd_sc_hd__or3b_1
Xclkbuf_leaf_109_clk clknet_4_10__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_109_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_19_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14789_ net997 ag2.body\[544\] vssd1 vssd1 vccd1 vccd1 _01460_ sky130_fd_sc_hd__xor2_1
XFILLER_0_46_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19316_ clknet_leaf_104_clk _00260_ net1435 vssd1 vssd1 vccd1 vccd1 control.body\[1074\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11281__A net1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16528_ net350 _02206_ vssd1 vssd1 vccd1 vccd1 _02207_ sky130_fd_sc_hd__nand2_1
XFILLER_0_50_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19247_ clknet_leaf_83_clk _00191_ net1482 vssd1 vssd1 vccd1 vccd1 ag2.body\[110\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_27_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16283__S net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16459_ _02057_ _02136_ _02137_ vssd1 vssd1 vccd1 vccd1 _02138_ sky130_fd_sc_hd__and3_1
XANTENNA__15545__A2 net162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18064__A net42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09000_ ag2.body\[101\] vssd1 vssd1 vccd1 vccd1 _04025_ sky130_fd_sc_hd__inv_2
XFILLER_0_61_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_3_7_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_3_7_0_clk sky130_fd_sc_hd__clkbuf_8
X_19178_ clknet_leaf_53_clk _00122_ net1365 vssd1 vssd1 vccd1 vccd1 ag2.body\[41\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_87_1380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18129_ _01691_ _03535_ net39 vssd1 vssd1 vccd1 vccd1 _03701_ sky130_fd_sc_hd__and3b_1
XFILLER_0_83_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11582__A3 _06554_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10344__B net1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11319__B1 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09902_ _04864_ _04872_ _04873_ _04874_ vssd1 vssd1 vccd1 vccd1 _04875_ sky130_fd_sc_hd__or4_1
XFILLER_0_1_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_35_1402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout504 net505 vssd1 vssd1 vccd1 vccd1 net504 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_6_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout515 _06464_ vssd1 vssd1 vccd1 vccd1 net515 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_6_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout526 net527 vssd1 vssd1 vccd1 vccd1 net526 sky130_fd_sc_hd__buf_2
X_20022_ clknet_leaf_58_clk _00966_ net1471 vssd1 vssd1 vccd1 vccd1 ag2.body\[372\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_6_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout537 _01707_ vssd1 vssd1 vccd1 vccd1 net537 sky130_fd_sc_hd__buf_2
X_09833_ net1107 control.body\[925\] vssd1 vssd1 vccd1 vccd1 _04806_ sky130_fd_sc_hd__or2_1
XFILLER_0_22_1559 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout548 net550 vssd1 vssd1 vccd1 vccd1 net548 sky130_fd_sc_hd__clkbuf_4
Xfanout559 net562 vssd1 vssd1 vccd1 vccd1 net559 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout290_A net294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09764_ ag2.body\[213\] net1114 vssd1 vssd1 vccd1 vccd1 _04737_ sky130_fd_sc_hd__xor2_1
XANTENNA__17470__A2 net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1340 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09695_ ag2.body\[71\] net1064 vssd1 vssd1 vccd1 vccd1 _04668_ sky130_fd_sc_hd__or2_1
XANTENNA__14767__A net1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout555_A _06651_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1297_A net1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13671__A net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17222__A2 net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19171__CLK clknet_leaf_53_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18739__CLK clknet_leaf_142_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15784__A2 net210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout722_A net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout343_X net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1464_A net1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1085_X net1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_3310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11191__A net1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_3321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17797__B net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18183__B1 net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout510_X net510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout608_X net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10470_ net1134 control.body\[1012\] vssd1 vssd1 vccd1 vccd1 _05443_ sky130_fd_sc_hd__xor2_1
XFILLER_0_66_1431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09129_ ag2.body\[434\] vssd1 vssd1 vccd1 vccd1 _04154_ sky130_fd_sc_hd__inv_2
XANTENNA__17289__A2 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14007__A net1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10535__A net1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12140_ img_gen.tracker.frame\[519\] net599 vssd1 vssd1 vccd1 vccd1 _07112_ sky130_fd_sc_hd__or2_1
XFILLER_0_102_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_1448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout977_X net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12071_ net1216 net1191 img_gen.tracker.frame\[105\] vssd1 vssd1 vccd1 vccd1 _07043_
+ sky130_fd_sc_hd__and3_1
XANTENNA__12750__A net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold580 control.body\[1116\] vssd1 vssd1 vccd1 vccd1 net2142 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold591 control.body\[908\] vssd1 vssd1 vccd1 vccd1 net2153 sky130_fd_sc_hd__dlygate4sd3_1
X_11022_ ag2.body\[597\] net1098 vssd1 vssd1 vccd1 vccd1 _05995_ sky130_fd_sc_hd__or2_1
XFILLER_0_60_1063 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17997__B1 net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11730__B1 _06649_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13057__S _07720_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11366__A net1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15830_ ag2.body\[256\] net175 net49 ag2.body\[248\] vssd1 vssd1 vccd1 vccd1 _01074_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_99_1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11085__B net1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15761_ ag2.body\[322\] net216 _01636_ ag2.body\[314\] vssd1 vssd1 vccd1 vccd1 _01012_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__13852__Y _08134_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12973_ _07683_ net254 _07681_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[247\]
+ sky130_fd_sc_hd__mux2_1
XANTENNA__14677__A net1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17500_ ag2.body\[237\] net951 vssd1 vssd1 vccd1 vccd1 _03179_ sky130_fd_sc_hd__xor2_1
XFILLER_0_137_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14712_ net1014 ag2.body\[343\] vssd1 vssd1 vccd1 vccd1 _08873_ sky130_fd_sc_hd__xor2_1
X_18480_ net1515 net1509 vssd1 vssd1 vccd1 vccd1 _00011_ sky130_fd_sc_hd__or2_1
X_11924_ img_gen.tracker.frame\[301\] net623 net577 vssd1 vssd1 vccd1 vccd1 _06896_
+ sky130_fd_sc_hd__o21ai_1
X_15692_ ag2.body\[390\] net140 _01616_ ag2.body\[382\] vssd1 vssd1 vccd1 vccd1 _00952_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12468__Y _07423_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17431_ _03104_ _03109_ vssd1 vssd1 vccd1 vccd1 _03110_ sky130_fd_sc_hd__nand2b_4
XTAP_TAPCELL_ROW_16_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14643_ net1002 ag2.body\[512\] vssd1 vssd1 vccd1 vccd1 _08804_ sky130_fd_sc_hd__xor2_1
X_11855_ img_gen.tracker.frame\[217\] net623 net607 img_gen.tracker.frame\[220\] _06826_
+ vssd1 vssd1 vccd1 vccd1 _06827_ sky130_fd_sc_hd__o221a_1
XANTENNA__16892__A ag2.body\[214\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10049__B1 _05021_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17362_ net1044 net1043 _03006_ vssd1 vssd1 vccd1 vccd1 _03041_ sky130_fd_sc_hd__o21a_1
XFILLER_0_55_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10806_ ag2.body\[35\] net1152 vssd1 vssd1 vccd1 vccd1 _05779_ sky130_fd_sc_hd__xor2_1
X_14574_ net973 ag2.body\[491\] vssd1 vssd1 vccd1 vccd1 _08735_ sky130_fd_sc_hd__nand2_1
X_11786_ img_gen.tracker.frame\[347\] net580 net542 img_gen.tracker.frame\[344\] _06757_
+ vssd1 vssd1 vccd1 vccd1 _06758_ sky130_fd_sc_hd__o221a_1
XFILLER_0_27_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11797__B1 net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19101_ clknet_leaf_145_clk img_gen.tracker.next_frame\[539\] net1242 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[539\] sky130_fd_sc_hd__dfrtp_1
X_16313_ obsg2.obstacleArray\[108\] net405 vssd1 vssd1 vccd1 vccd1 _01992_ sky130_fd_sc_hd__or2_1
X_13525_ net2092 net655 _07921_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[561\]
+ sky130_fd_sc_hd__and3_1
XFILLER_0_32_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17293_ ag2.body\[346\] net865 vssd1 vssd1 vccd1 vccd1 _02972_ sky130_fd_sc_hd__xor2_1
XANTENNA__17500__B net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10737_ ag2.body\[251\] net770 _05707_ _05708_ _05709_ vssd1 vssd1 vccd1 vccd1 _05710_
+ sky130_fd_sc_hd__o2111ai_4
XANTENNA__11892__S0 net1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14843__C _08924_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13538__A1 net226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19032_ clknet_leaf_6_clk img_gen.tracker.next_frame\[470\] net1264 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[470\] sky130_fd_sc_hd__dfrtp_1
X_16244_ obsg2.obstacleArray\[44\] obsg2.obstacleArray\[45\] net404 vssd1 vssd1 vccd1
+ vccd1 _01923_ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_2103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13456_ net682 _07894_ vssd1 vssd1 vccd1 vccd1 _07895_ sky130_fd_sc_hd__nor2_1
XFILLER_0_84_1520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10668_ net762 control.body\[884\] control.body\[887\] net746 _05637_ vssd1 vssd1
+ vccd1 vccd1 _05641_ sky130_fd_sc_hd__o221ai_1
XFILLER_0_84_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15020__B net59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12407_ _06477_ _07369_ _07355_ vssd1 vssd1 vccd1 vccd1 _07370_ sky130_fd_sc_hd__a21oi_1
X_16175_ _01728_ _01845_ _01853_ vssd1 vssd1 vccd1 vccd1 _01854_ sky130_fd_sc_hd__or3_1
XFILLER_0_49_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10599_ _05567_ _05570_ _05571_ vssd1 vssd1 vccd1 vccd1 _05572_ sky130_fd_sc_hd__or3_1
XFILLER_0_23_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13387_ _07546_ net304 vssd1 vssd1 vccd1 vccd1 _07868_ sky130_fd_sc_hd__nor2_1
XFILLER_0_112_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15126_ control.body\[894\] net107 _01565_ control.body\[886\] vssd1 vssd1 vccd1
+ vccd1 _00448_ sky130_fd_sc_hd__a22o_1
X_12338_ net628 net467 net563 vssd1 vssd1 vccd1 vccd1 _07305_ sky130_fd_sc_hd__and3_1
XANTENNA__15955__B net60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14161__A1_N net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10164__B net1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19934_ clknet_leaf_47_clk _00878_ net1375 vssd1 vssd1 vccd1 vccd1 ag2.body\[460\]
+ sky130_fd_sc_hd__dfrtp_2
X_15057_ _04759_ _01554_ vssd1 vssd1 vccd1 vccd1 _01559_ sky130_fd_sc_hd__and2b_2
X_12269_ img_gen.updater.commands.count\[8\] img_gen.updater.commands.count\[9\] img_gen.updater.commands.count\[2\]
+ vssd1 vssd1 vccd1 vccd1 _07239_ sky130_fd_sc_hd__nand3_1
X_14008_ net837 ag2.body\[505\] _04185_ net984 vssd1 vssd1 vccd1 vccd1 _08169_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__13710__A1 _04239_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11316__A3 _06277_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19865_ clknet_leaf_94_clk _00809_ net1437 vssd1 vssd1 vccd1 vccd1 ag2.body\[535\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_120_1451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11721__B1 net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17452__A2 net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18816_ clknet_leaf_3_clk img_gen.tracker.next_frame\[254\] net1259 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[254\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_128_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19194__CLK clknet_leaf_53_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19796_ clknet_leaf_127_clk _00740_ net1328 vssd1 vssd1 vccd1 vccd1 ag2.body\[594\]
+ sky130_fd_sc_hd__dfrtp_4
X_15959_ ag2.body\[147\] net198 _01657_ ag2.body\[139\] vssd1 vssd1 vccd1 vccd1 _01189_
+ sky130_fd_sc_hd__a22o_1
X_18747_ clknet_leaf_139_clk img_gen.tracker.next_frame\[185\] net1256 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[185\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_91_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_95_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13491__A net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09480_ _04166_ net1155 net748 ag2.body\[470\] _04452_ vssd1 vssd1 vccd1 vccd1 _04453_
+ sky130_fd_sc_hd__o221a_1
X_18678_ clknet_leaf_27_clk img_gen.tracker.next_frame\[116\] net1339 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[116\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_56_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17629_ ag2.body\[187\] net717 net714 ag2.body\[188\] vssd1 vssd1 vccd1 vccd1 _03308_
+ sky130_fd_sc_hd__o22a_1
XANTENNA__17898__A net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20097__Q ag2.body\[303\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11788__B1 net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17410__B net875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20571_ clknet_leaf_107_clk _01429_ _00035_ vssd1 vssd1 vccd1 vccd1 sound_gen.dac1.dacCount\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_46_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout136_A net139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12835__A _07431_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_1004 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12201__A1 net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout303_A net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1045_A net1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1172 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_498 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15865__B net66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09863__B net1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1212_A net1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout301 _03545_ vssd1 vssd1 vccd1 vccd1 net301 sky130_fd_sc_hd__buf_2
XANTENNA__19537__CLK clknet_leaf_118_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout312 net313 vssd1 vssd1 vccd1 vccd1 net312 sky130_fd_sc_hd__buf_2
Xfanout323 net324 vssd1 vssd1 vccd1 vccd1 net323 sky130_fd_sc_hd__buf_2
Xfanout334 _07423_ vssd1 vssd1 vccd1 vccd1 net334 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09582__C net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout293_X net293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout672_A net674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout345 _03541_ vssd1 vssd1 vccd1 vccd1 net345 sky130_fd_sc_hd__buf_2
X_20005_ clknet_leaf_59_clk _00949_ net1468 vssd1 vssd1 vccd1 vccd1 ag2.body\[387\]
+ sky130_fd_sc_hd__dfrtp_4
Xfanout367 _02067_ vssd1 vssd1 vccd1 vccd1 net367 sky130_fd_sc_hd__clkbuf_2
X_09816_ net1206 control.body\[1049\] vssd1 vssd1 vccd1 vccd1 _04789_ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout1000_X net1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17443__A2 net862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout378 net379 vssd1 vssd1 vccd1 vccd1 net378 sky130_fd_sc_hd__buf_4
XFILLER_0_103_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__20514__CLK clknet_leaf_113_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16651__B1 net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09747_ ag2.body\[353\] net1213 vssd1 vssd1 vccd1 vccd1 _04720_ sky130_fd_sc_hd__xor2_1
XANTENNA_fanout460_X net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18561__CLK clknet_leaf_132_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout937_A net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout558_X net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09678_ ag2.body\[10\] net1175 vssd1 vssd1 vccd1 vccd1 _04651_ sky130_fd_sc_hd__or2_1
XFILLER_0_115_1019 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout49_A _01631_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout725_X net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11640_ obsg2.obstacleArray\[129\] obsg2.obstacleArray\[133\] net513 vssd1 vssd1
+ vccd1 vccd1 _06613_ sky130_fd_sc_hd__mux2_1
XANTENNA__14965__B1 _01547_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_209 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10249__B _05212_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11779__B1 net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_2_0_clk_X clknet_3_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17320__B net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11571_ obsg2.obstacleArray\[90\] obsg2.obstacleArray\[91\] obsg2.obstacleArray\[94\]
+ obsg2.obstacleArray\[95\] net1125 net512 vssd1 vssd1 vccd1 vccd1 _06544_ sky130_fd_sc_hd__mux4_1
XFILLER_0_65_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12745__A net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_30_Left_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13310_ net2114 net647 _07837_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[430\]
+ sky130_fd_sc_hd__and3_1
XFILLER_0_68_1526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10522_ _05476_ _05484_ _05489_ _05494_ vssd1 vssd1 vccd1 vccd1 _05495_ sky130_fd_sc_hd__a22o_1
X_14290_ net811 ag2.body\[476\] ag2.body\[477\] net806 _08449_ vssd1 vssd1 vccd1 vccd1
+ _08451_ sky130_fd_sc_hd__a221o_1
XFILLER_0_24_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10560__A_N net1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10453_ ag2.body\[454\] net1079 vssd1 vssd1 vccd1 vccd1 _05426_ sky130_fd_sc_hd__nand2_1
X_13241_ net283 _07808_ _07809_ net1857 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[389\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__10265__A net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10384_ _05353_ _05354_ _05355_ _05356_ vssd1 vssd1 vccd1 vccd1 _05357_ sky130_fd_sc_hd__or4_1
X_13172_ _07777_ net252 _07775_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[352\]
+ sky130_fd_sc_hd__mux2_1
XANTENNA__10754__A1 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10792__D_N _05685_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16223__Y _01902_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10754__B2 net1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12123_ img_gen.tracker.frame\[546\] net541 net568 vssd1 vssd1 vccd1 vccd1 _07095_
+ sky130_fd_sc_hd__o21a_1
XANTENNA__10415__D _05387_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17980_ net39 _03600_ vssd1 vssd1 vccd1 vccd1 _03601_ sky130_fd_sc_hd__and2_1
XANTENNA__09773__B net1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16931_ _02606_ _02607_ _02609_ vssd1 vssd1 vccd1 vccd1 _02610_ sky130_fd_sc_hd__nand3b_1
X_12054_ net1215 net1190 img_gen.tracker.frame\[81\] vssd1 vssd1 vccd1 vccd1 _07026_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_44_1592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19272__RESET_B net1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18904__CLK clknet_leaf_144_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11005_ net770 control.body\[1083\] control.body\[1084\] net761 vssd1 vssd1 vccd1
+ vccd1 _05978_ sky130_fd_sc_hd__o22a_1
X_16862_ ag2.body\[207\] net933 vssd1 vssd1 vccd1 vccd1 _02541_ sky130_fd_sc_hd__nand2_1
X_19650_ clknet_leaf_119_clk _00594_ net1308 vssd1 vssd1 vccd1 vccd1 control.body\[736\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_74_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19201__RESET_B net1461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15813_ ag2.body\[272\] net206 _01642_ ag2.body\[264\] vssd1 vssd1 vccd1 vccd1 _01058_
+ sky130_fd_sc_hd__a22o_1
Xfanout890 net891 vssd1 vssd1 vccd1 vccd1 net890 sky130_fd_sc_hd__clkbuf_4
X_18601_ clknet_leaf_16_clk img_gen.tracker.next_frame\[39\] net1320 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[39\] sky130_fd_sc_hd__dfrtp_1
X_19581_ clknet_leaf_116_clk _00525_ net1385 vssd1 vssd1 vccd1 vccd1 control.body\[811\]
+ sky130_fd_sc_hd__dfrtp_1
X_16793_ net399 _02469_ _02471_ net363 vssd1 vssd1 vccd1 vccd1 _02472_ sky130_fd_sc_hd__o211a_1
XFILLER_0_137_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18532_ clknet_leaf_137_clk _00058_ net1298 vssd1 vssd1 vccd1 vccd1 img_gen.updater.commands.count\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_15744_ ag2.body\[339\] net215 _01634_ ag2.body\[331\] vssd1 vssd1 vccd1 vccd1 _00997_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_87_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12956_ _07675_ net268 _07673_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[238\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18463_ net883 net871 net861 _03950_ vssd1 vssd1 vccd1 vccd1 _03951_ sky130_fd_sc_hd__a31o_1
X_11907_ img_gen.tracker.frame\[364\] net605 _06877_ _06878_ vssd1 vssd1 vccd1 vccd1
+ _06879_ sky130_fd_sc_hd__o211a_1
X_15675_ ag2.body\[406\] net142 _01626_ ag2.body\[398\] vssd1 vssd1 vccd1 vccd1 _00936_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11482__A2 _06440_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12887_ net678 _07643_ vssd1 vssd1 vccd1 vccd1 _07644_ sky130_fd_sc_hd__nor2_1
X_17414_ ag2.body\[282\] net727 net951 _04096_ _03090_ vssd1 vssd1 vccd1 vccd1 _03093_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_5_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12461__A_N _06644_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14626_ net1008 ag2.body\[471\] vssd1 vssd1 vccd1 vccd1 _08787_ sky130_fd_sc_hd__xor2_1
XFILLER_0_16_1650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18394_ _03812_ _03872_ vssd1 vssd1 vccd1 vccd1 _03884_ sky130_fd_sc_hd__nor2_1
X_11838_ _06803_ _06805_ _06807_ _06809_ net558 net471 vssd1 vssd1 vccd1 vccd1 _06810_
+ sky130_fd_sc_hd__mux4_1
XANTENNA__14956__B1 _01546_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17345_ _03013_ _03017_ _03021_ _03023_ vssd1 vssd1 vccd1 vccd1 _03024_ sky130_fd_sc_hd__or4_1
X_14557_ net990 ag2.body\[65\] vssd1 vssd1 vccd1 vccd1 _08718_ sky130_fd_sc_hd__xor2_1
XFILLER_0_56_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_99_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11769_ net559 _06740_ _06738_ net471 vssd1 vssd1 vccd1 vccd1 _06741_ sky130_fd_sc_hd__a211o_1
XANTENNA__12655__A _06671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_40_clk clknet_4_7__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_40_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_12_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13508_ net250 _07914_ _07915_ net1652 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[550\]
+ sky130_fd_sc_hd__a22o_1
X_17276_ ag2.body\[556\] net962 vssd1 vssd1 vccd1 vccd1 _02955_ sky130_fd_sc_hd__nand2_1
X_14488_ net985 ag2.body\[346\] vssd1 vssd1 vccd1 vccd1 _08649_ sky130_fd_sc_hd__xor2_1
XFILLER_0_82_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_1313 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19015_ clknet_leaf_1_clk img_gen.tracker.next_frame\[453\] net1246 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[453\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_71_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16227_ net496 _01897_ vssd1 vssd1 vccd1 vccd1 _01906_ sky130_fd_sc_hd__nor2_1
XANTENNA__14184__A1 net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_741 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13439_ net282 _07886_ _07887_ net1812 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[509\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_80_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16158_ _01743_ _01823_ _01827_ _01836_ vssd1 vssd1 vccd1 vccd1 _01837_ sky130_fd_sc_hd__a31o_1
XANTENNA__13931__B2 ag2.body\[66\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15109_ net2533 net145 _01564_ control.body\[902\] vssd1 vssd1 vccd1 vccd1 _00432_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__09683__B net1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17673__A2 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10462__X _05435_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08980_ ag2.body\[74\] vssd1 vssd1 vccd1 vccd1 _04005_ sky130_fd_sc_hd__inv_2
X_16089_ obsg2.obstacleArray\[100\] obsg2.obstacleArray\[101\] net425 vssd1 vssd1
+ vccd1 vccd1 _01768_ sky130_fd_sc_hd__mux2_1
XANTENNA__10903__A net1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19917_ clknet_leaf_55_clk _00861_ net1456 vssd1 vssd1 vccd1 vccd1 ag2.body\[475\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_97_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10622__B net1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19848_ clknet_leaf_93_clk _00792_ net1413 vssd1 vssd1 vccd1 vccd1 ag2.body\[550\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_120_1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16633__B1 net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09601_ net640 _04571_ net643 vssd1 vssd1 vccd1 vccd1 _04574_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_78_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19779_ clknet_leaf_127_clk _00723_ net1327 vssd1 vssd1 vccd1 vccd1 ag2.body\[609\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_79_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09532_ net1206 control.body\[1025\] vssd1 vssd1 vccd1 vccd1 _04505_ sky130_fd_sc_hd__and2b_1
XFILLER_0_56_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14110__A net1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09463_ ag2.body\[382\] net1080 vssd1 vssd1 vccd1 vccd1 _04436_ sky130_fd_sc_hd__xor2_1
XANTENNA_fanout253_A net254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09394_ sound_gen.osc1.stayCount\[5\] _04344_ sound_gen.osc1.stayCount\[6\] vssd1
+ vssd1 vccd1 vccd1 _04381_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_93_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17140__B net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20623_ img_gen.updater.update.wr vssd1 vssd1 vccd1 vccd1 net34 sky130_fd_sc_hd__clkbuf_1
XANTENNA__12422__A1 net1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10637__X _05610_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_31_clk clknet_4_4__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_31_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__15579__C net64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1162_A net1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout139_X net139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout518_A net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20554_ clknet_leaf_106_clk _01419_ _00028_ vssd1 vssd1 vccd1 vccd1 sound_gen.osc1.stayCount\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_117_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__20067__CLK clknet_leaf_73_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20485_ clknet_leaf_37_clk _01372_ net1353 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[121\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_85_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10085__A net1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18252__A _03693_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14780__A net1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1048_X net1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09874__A ag2.body\[167\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13922__A1 ag2.body\[66\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13922__B2 ag2.body\[58\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout887_A net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17664__A2 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16321__C1 net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_3671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1215_X net1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_110_3682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_110_3693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1107 net1109 vssd1 vssd1 vccd1 vccd1 net1107 sky130_fd_sc_hd__clkbuf_4
Xfanout120 net128 vssd1 vssd1 vccd1 vccd1 net120 sky130_fd_sc_hd__clkbuf_2
Xfanout1118 net1119 vssd1 vssd1 vccd1 vccd1 net1118 sky130_fd_sc_hd__buf_4
Xfanout131 net132 vssd1 vssd1 vccd1 vccd1 net131 sky130_fd_sc_hd__buf_2
Xfanout1129 ag2.x\[0\] vssd1 vssd1 vccd1 vccd1 net1129 sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout675_X net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_98_clk clknet_4_11__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_98_clk
+ sky130_fd_sc_hd__clkbuf_8
Xfanout142 net143 vssd1 vssd1 vccd1 vccd1 net142 sky130_fd_sc_hd__buf_2
XANTENNA__17416__A2 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout153 net154 vssd1 vssd1 vccd1 vccd1 net153 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_96_1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout164 net165 vssd1 vssd1 vccd1 vccd1 net164 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout175 net176 vssd1 vssd1 vccd1 vccd1 net175 sky130_fd_sc_hd__clkbuf_4
Xfanout186 net187 vssd1 vssd1 vccd1 vccd1 net186 sky130_fd_sc_hd__clkbuf_2
XANTENNA__14939__B _04792_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout197 net200 vssd1 vssd1 vccd1 vccd1 net197 sky130_fd_sc_hd__buf_2
XANTENNA__13843__B net56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout842_X net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_1530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12810_ net286 _07605_ _07606_ net1917 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[161\]
+ sky130_fd_sc_hd__a22o_1
X_13790_ _07195_ _07213_ vssd1 vssd1 vccd1 vccd1 _08097_ sky130_fd_sc_hd__nor2_1
XFILLER_0_39_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12110__B1 net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_3486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_3497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12741_ net258 _07573_ _07574_ net1636 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[124\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_69_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15460_ ag2.body\[599\] net89 _01602_ ag2.body\[591\] vssd1 vssd1 vccd1 vccd1 _00745_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_96_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12672_ net267 _07540_ _07541_ net1625 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[88\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_127_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14411_ net981 _03967_ net1036 _03970_ vssd1 vssd1 vccd1 vccd1 _08572_ sky130_fd_sc_hd__a22o_1
X_11623_ _06588_ _06595_ _06497_ vssd1 vssd1 vccd1 vccd1 _06596_ sky130_fd_sc_hd__or3b_1
XFILLER_0_37_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15391_ net2302 net82 _01596_ net2500 vssd1 vssd1 vccd1 vccd1 _00682_ sky130_fd_sc_hd__a22o_1
XANTENNA__09768__B net1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11847__S0 net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_22_clk clknet_4_6__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_22_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_52_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17130_ _04188_ net874 net853 _04190_ vssd1 vssd1 vccd1 vccd1 _02809_ sky130_fd_sc_hd__o22a_1
XFILLER_0_37_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14342_ net979 ag2.body\[610\] vssd1 vssd1 vccd1 vccd1 _08503_ sky130_fd_sc_hd__xor2_1
XANTENNA__11621__C1 net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11554_ _06509_ _06526_ vssd1 vssd1 vccd1 vccd1 _06527_ sky130_fd_sc_hd__nand2b_1
XANTENNA__10707__B net1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14166__A1 net980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17061_ _04006_ net855 net935 _04010_ vssd1 vssd1 vccd1 vccd1 _02740_ sky130_fd_sc_hd__o22a_1
X_10505_ net769 control.body\[979\] control.body\[981\] net755 _05477_ vssd1 vssd1
+ vccd1 vccd1 _05478_ sky130_fd_sc_hd__a221o_1
X_14273_ _08424_ _08425_ _08426_ _08427_ vssd1 vssd1 vccd1 vccd1 _08434_ sky130_fd_sc_hd__a22o_1
XANTENNA__14166__B2 net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11485_ _05389_ _05839_ _06018_ _06457_ vssd1 vssd1 vccd1 vccd1 _06458_ sky130_fd_sc_hd__or4b_1
XFILLER_0_100_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12177__B1 net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16012_ net858 net848 vssd1 vssd1 vccd1 vccd1 _01691_ sky130_fd_sc_hd__nor2_2
XFILLER_0_85_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13913__A1 ag2.body\[58\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09784__A net1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13224_ net289 _07799_ _07800_ net2088 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[380\]
+ sky130_fd_sc_hd__a22o_1
X_10436_ net1083 control.body\[934\] vssd1 vssd1 vccd1 vccd1 _05409_ sky130_fd_sc_hd__nor2_1
XFILLER_0_0_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11924__B1 net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15115__B1 _01554_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10282__X _05255_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13155_ _07769_ net252 _07767_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[343\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10367_ _05339_ _05337_ _05336_ _05338_ vssd1 vssd1 vccd1 vccd1 _05340_ sky130_fd_sc_hd__or4bb_1
X_12106_ net472 _07077_ _07071_ _06661_ vssd1 vssd1 vccd1 vccd1 _07078_ sky130_fd_sc_hd__a211o_1
XANTENNA__20358__RESET_B net1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10298_ _05239_ _05252_ _05255_ _05270_ vssd1 vssd1 vccd1 vccd1 _05271_ sky130_fd_sc_hd__o22a_2
XFILLER_0_97_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17963_ net318 _03587_ obsg2.obstacleArray\[11\] vssd1 vssd1 vccd1 vccd1 _03588_
+ sky130_fd_sc_hd__a21oi_1
X_13086_ _07736_ net265 _07734_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[307\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_1118 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_89_clk clknet_4_9__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_89_clk
+ sky130_fd_sc_hd__clkbuf_8
X_19702_ clknet_leaf_134_clk net2560 net1307 vssd1 vssd1 vccd1 vccd1 control.body\[692\]
+ sky130_fd_sc_hd__dfrtp_1
X_12037_ img_gen.tracker.frame\[9\] net594 net557 img_gen.tracker.frame\[6\] _07008_
+ vssd1 vssd1 vccd1 vccd1 _07009_ sky130_fd_sc_hd__a221o_1
X_16914_ ag2.body\[560\] net881 vssd1 vssd1 vccd1 vccd1 _02593_ sky130_fd_sc_hd__nand2_1
XANTENNA__17407__A2 net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17894_ obsg2.obstacleCount\[1\] _03531_ _03532_ _03523_ vssd1 vssd1 vccd1 vccd1
+ _01248_ sky130_fd_sc_hd__a22o_1
XANTENNA__16615__B1 net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19633_ clknet_leaf_123_clk _00577_ net1406 vssd1 vssd1 vccd1 vccd1 control.body\[767\]
+ sky130_fd_sc_hd__dfrtp_1
X_16845_ ag2.body\[175\] net691 vssd1 vssd1 vccd1 vccd1 _02524_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_0_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16776_ obsg2.obstacleArray\[28\] net494 _02454_ vssd1 vssd1 vccd1 vccd1 _02455_
+ sky130_fd_sc_hd__a21o_1
X_19564_ clknet_leaf_116_clk _00508_ net1387 vssd1 vssd1 vccd1 vccd1 control.body\[826\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_117_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13988_ ag2.body\[125\] net211 _08159_ ag2.body\[117\] vssd1 vssd1 vccd1 vccd1 _00206_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12101__B1 net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12369__B _07301_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09024__A ag2.body\[160\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15727_ ag2.body\[356\] net197 _01632_ ag2.body\[348\] vssd1 vssd1 vccd1 vccd1 _00982_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11273__B net1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18515_ net1512 net1506 vssd1 vssd1 vccd1 vccd1 _00046_ sky130_fd_sc_hd__or2_1
XANTENNA__19232__CLK clknet_leaf_75_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12652__A1 net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12939_ net294 _07665_ _07666_ net1747 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[230\]
+ sky130_fd_sc_hd__a22o_1
X_19495_ clknet_leaf_113_clk _00439_ net1399 vssd1 vssd1 vccd1 vccd1 control.body\[901\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__17040__B1 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1658 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14929__B1 _01543_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15658_ ag2.body\[423\] net138 _01624_ ag2.body\[415\] vssd1 vssd1 vccd1 vccd1 _00921_
+ sky130_fd_sc_hd__a22o_1
X_18446_ _03828_ _03933_ _03934_ vssd1 vssd1 vccd1 vccd1 _03935_ sky130_fd_sc_hd__or3b_1
XFILLER_0_69_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17591__B2 ag2.body\[62\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14609_ net1003 _04033_ ag2.body\[131\] net822 _08769_ vssd1 vssd1 vccd1 vccd1 _08770_
+ sky130_fd_sc_hd__o221a_1
XANTENNA__09678__B net1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18377_ _08022_ _03867_ vssd1 vssd1 vccd1 vccd1 _03868_ sky130_fd_sc_hd__nand2_1
X_15589_ ag2.body\[472\] net122 _01618_ ag2.body\[464\] vssd1 vssd1 vccd1 vccd1 _00858_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11838__S0 net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_13_clk clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_13_clk
+ sky130_fd_sc_hd__clkbuf_8
X_17328_ ag2.body\[3\] net850 vssd1 vssd1 vccd1 vccd1 _03007_ sky130_fd_sc_hd__xor2_2
XANTENNA__19382__CLK clknet_leaf_102_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16146__A2 net427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_133_4372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_133_4383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14157__A1 net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_133_4394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17259_ _02933_ _02935_ _02936_ _02937_ vssd1 vssd1 vccd1 vccd1 _02938_ sky130_fd_sc_hd__or4_1
XANTENNA__14157__B2 net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16291__S net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17894__A2 _03531_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18072__A net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12168__B1 net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09694__A ag2.body\[71\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20270_ clknet_leaf_36_clk net1576 net1347 vssd1 vssd1 vccd1 vccd1 control.detect1.Q\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_1000 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_wire476_X net476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13928__B net61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19194__RESET_B net1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16304__B net413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14105__A net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08963_ ag2.body\[42\] vssd1 vssd1 vccd1 vccd1 _03988_ sky130_fd_sc_hd__inv_2
XFILLER_0_45_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_1994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20028__RESET_B net1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_127_4187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_4198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09887__A2 net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1008_A net1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17135__B net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11694__A2 net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout468_A _06648_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09205__Y _04230_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16974__B net851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11183__B net1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09515_ net1149 control.body\[835\] vssd1 vssd1 vccd1 vccd1 _04488_ sky130_fd_sc_hd__or2_1
XANTENNA__10779__A2_N _05751_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12643__A1 net242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout256_X net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14775__A net1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1377_A net1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09446_ net891 net898 net901 vssd1 vssd1 vccd1 vccd1 _04419_ sky130_fd_sc_hd__or3_4
XFILLER_0_109_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_1080 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14396__A1 net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout802_A net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14396__B2 net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout423_X net423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09377_ net273 _04360_ _04373_ vssd1 vssd1 vccd1 vccd1 _01415_ sky130_fd_sc_hd__nor3_1
XANTENNA_fanout1165_X net1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20606_ net1538 vssd1 vssd1 vccd1 vccd1 gpio_oeb[18] sky130_fd_sc_hd__buf_2
XANTENNA__11603__C1 net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17300__A2_N net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20537_ clknet_leaf_106_clk _01402_ _00011_ vssd1 vssd1 vccd1 vccd1 sound_gen.osc1.stayCount\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17885__A2 _04239_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_104_Left_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1332_X net1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_3733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_3744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11270_ ag2.body\[127\] net1067 vssd1 vssd1 vccd1 vccd1 _06243_ sky130_fd_sc_hd__or2_1
X_20468_ clknet_leaf_33_clk _01355_ net1346 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[104\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_15_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout792_X net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11906__B1 net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17098__B1 net719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10221_ ag2.body\[562\] net1172 vssd1 vssd1 vccd1 vccd1 _05194_ sky130_fd_sc_hd__nand2_1
X_20399_ clknet_leaf_28_clk _01286_ net1340 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[35\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_63_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10152_ _03997_ net1104 net1057 _03998_ vssd1 vssd1 vccd1 vccd1 _05125_ sky130_fd_sc_hd__a22o_1
XFILLER_0_63_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10083_ net1050 control.body\[799\] vssd1 vssd1 vccd1 vccd1 _05056_ sky130_fd_sc_hd__or2_1
X_14960_ control.body\[1034\] net166 _01547_ net2278 vssd1 vssd1 vccd1 vccd1 _00300_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__08948__A net1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold9 control.button1.Q\[0\] vssd1 vssd1 vccd1 vccd1 net1571 sky130_fd_sc_hd__dlygate4sd3_1
X_13911_ ag2.body\[56\] net120 _08151_ ag2.body\[48\] vssd1 vssd1 vccd1 vccd1 _00137_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__14871__A2 net182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_3548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19255__CLK clknet_leaf_75_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17045__B net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14891_ control.body\[1101\] net180 _01539_ control.body\[1093\] vssd1 vssd1 vccd1
+ vccd1 _00239_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_113_Left_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_106_3559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16630_ obsg2.obstacleArray\[62\] net444 vssd1 vssd1 vccd1 vccd1 _02309_ sky130_fd_sc_hd__or2_1
X_13842_ net686 net223 vssd1 vssd1 vccd1 vccd1 _08132_ sky130_fd_sc_hd__or2_1
XFILLER_0_57_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__20232__CLK clknet_leaf_66_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16561_ net361 _02239_ _02236_ net357 vssd1 vssd1 vccd1 vccd1 _02240_ sky130_fd_sc_hd__o211a_1
XFILLER_0_97_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13773_ img_gen.updater.commands.count\[9\] _08084_ vssd1 vssd1 vccd1 vccd1 _08085_
+ sky130_fd_sc_hd__nand2b_1
XFILLER_0_69_254 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_2880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10985_ net1193 control.body\[753\] vssd1 vssd1 vccd1 vccd1 _05958_ sky130_fd_sc_hd__xor2_1
XANTENNA__18157__A net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17022__B1 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_2891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18300_ net322 _08136_ vssd1 vssd1 vccd1 vccd1 _03796_ sky130_fd_sc_hd__nand2_1
X_15512_ ag2.body\[549\] net155 _01608_ ag2.body\[541\] vssd1 vssd1 vccd1 vccd1 _00791_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_69_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19280_ clknet_leaf_97_clk net2126 net1450 vssd1 vssd1 vccd1 vccd1 control.body\[1118\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10645__B1 _05610_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12724_ net258 _07565_ _07566_ net1867 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[115\]
+ sky130_fd_sc_hd__a22o_1
X_16492_ obsg2.obstacleArray\[26\] obsg2.obstacleArray\[27\] net458 vssd1 vssd1 vccd1
+ vccd1 _02171_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17573__A1 ag2.body\[339\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_2755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17573__B2 ag2.body\[340\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_1534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_80_2766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12476__Y _07431_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18231_ net526 _03754_ vssd1 vssd1 vccd1 vccd1 _01363_ sky130_fd_sc_hd__and2_1
XANTENNA__12917__B net340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14387__A1 net975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_2777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15443_ _05451_ net54 vssd1 vssd1 vccd1 vccd1 _01601_ sky130_fd_sc_hd__nor2_4
XANTENNA__17996__A net46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14387__B2 net1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12655_ _06671_ _07531_ vssd1 vssd1 vccd1 vccd1 _07532_ sky130_fd_sc_hd__or2_2
XANTENNA__09498__B net919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16781__C1 net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_2176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_2187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_983 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_61_2198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09929__D _04901_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11606_ obsg2.obstacleArray\[24\] obsg2.obstacleArray\[25\] obsg2.obstacleArray\[28\]
+ obsg2.obstacleArray\[29\] net1126 net514 vssd1 vssd1 vccd1 vccd1 _06579_ sky130_fd_sc_hd__mux4_1
X_18162_ _03598_ net36 vssd1 vssd1 vccd1 vccd1 _03720_ sky130_fd_sc_hd__nor2_1
XFILLER_0_136_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15374_ net2234 net68 _01594_ net2369 vssd1 vssd1 vccd1 vccd1 _00667_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_122_Left_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12586_ net598 net471 net569 _07312_ vssd1 vssd1 vccd1 vccd1 _07493_ sky130_fd_sc_hd__or4_1
XFILLER_0_26_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14691__Y _08852_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10948__A1 net907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17113_ ag2.body\[537\] net735 net727 ag2.body\[538\] _02791_ vssd1 vssd1 vccd1 vccd1
+ _02792_ sky130_fd_sc_hd__o221a_1
X_14325_ net835 ag2.body\[449\] ag2.body\[450\] net825 vssd1 vssd1 vccd1 vccd1 _08486_
+ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__11070__B1 net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18093_ net38 _03677_ obsg2.obstacleArray\[51\] vssd1 vssd1 vccd1 vccd1 _03678_ sky130_fd_sc_hd__a21oi_1
X_11537_ _06495_ _06508_ vssd1 vssd1 vccd1 vccd1 _06510_ sky130_fd_sc_hd__nand2_1
XFILLER_0_41_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_1164 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20609__1541 vssd1 vssd1 vccd1 vccd1 _20609__1541/HI net1541 sky130_fd_sc_hd__conb_1
XFILLER_0_13_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16405__A net354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17044_ ag2.body\[261\] net951 vssd1 vssd1 vccd1 vccd1 _02723_ sky130_fd_sc_hd__xor2_1
Xhold409 img_gen.tracker.frame\[98\] vssd1 vssd1 vccd1 vccd1 net1971 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14851__C _08683_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_705 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14256_ net977 _04006_ _04009_ net1023 _08414_ vssd1 vssd1 vccd1 vccd1 _08417_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_78_2695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11468_ net920 _04599_ _04982_ _04687_ vssd1 vssd1 vccd1 vccd1 _06441_ sky130_fd_sc_hd__o31a_1
XANTENNA__16124__B net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13207_ net289 _07791_ _07792_ net1959 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[371\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__09566__A1 net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17628__A2 net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10419_ net1183 control.body\[1066\] vssd1 vssd1 vccd1 vccd1 _05392_ sky130_fd_sc_hd__xor2_1
XFILLER_0_46_1473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14187_ net1016 ag2.body\[166\] vssd1 vssd1 vccd1 vccd1 _08348_ sky130_fd_sc_hd__nand2_1
XFILLER_0_42_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11399_ ag2.body\[575\] net1052 vssd1 vssd1 vccd1 vccd1 _06372_ sky130_fd_sc_hd__nand2_1
XANTENNA__11268__B net1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13138_ _07758_ _07760_ _07761_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[334\]
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_104_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18995_ clknet_leaf_0_clk img_gen.tracker.next_frame\[433\] net1244 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[433\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09961__B net1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17946_ net48 net296 _03574_ vssd1 vssd1 vccd1 vccd1 _03575_ sky130_fd_sc_hd__and3_1
X_13069_ _07728_ net268 _07726_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[298\]
+ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_131_Left_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_2_clk clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_2_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__18587__RESET_B net1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_119_Right_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1460 net1461 vssd1 vssd1 vccd1 vccd1 net1460 sky130_fd_sc_hd__clkbuf_4
Xfanout1471 net1473 vssd1 vssd1 vccd1 vccd1 net1471 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_122_4040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1482 net1483 vssd1 vssd1 vccd1 vccd1 net1482 sky130_fd_sc_hd__clkbuf_4
X_17877_ net2130 _03507_ vssd1 vssd1 vccd1 vccd1 _01246_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_122_4051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1493 net1505 vssd1 vssd1 vccd1 vccd1 net1493 sky130_fd_sc_hd__clkbuf_2
XANTENNA__11284__A net1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19616_ clknet_leaf_119_clk _00560_ net1391 vssd1 vssd1 vccd1 vccd1 control.body\[782\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10884__B1 _05856_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16828_ ag2.body\[226\] net726 net943 _04071_ _02506_ vssd1 vssd1 vccd1 vccd1 _02507_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_88_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12625__A1 net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19547_ clknet_leaf_115_clk _00491_ net1397 vssd1 vssd1 vccd1 vccd1 control.body\[841\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__16286__S net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16759_ obsg2.obstacleArray\[16\] net494 net485 obsg2.obstacleArray\[17\] _02437_
+ vssd1 vssd1 vccd1 vccd1 _02438_ sky130_fd_sc_hd__a221o_1
XANTENNA__14595__A net993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18067__A net42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09300_ sound_gen.osc1.count\[1\] sound_gen.osc1.count\[0\] vssd1 vssd1 vccd1 vccd1
+ _04320_ sky130_fd_sc_hd__nand2_1
XFILLER_0_53_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19478_ clknet_leaf_110_clk _00422_ net1418 vssd1 vssd1 vccd1 vccd1 control.body\[916\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_64_909 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_769 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_135_4434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09231_ control.body\[1096\] vssd1 vssd1 vccd1 vccd1 _04256_ sky130_fd_sc_hd__inv_2
XFILLER_0_118_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18429_ _03792_ _03915_ vssd1 vssd1 vccd1 vccd1 _03918_ sky130_fd_sc_hd__nor2_1
XANTENNA__18772__CLK clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_135_4445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10187__X _05160_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10628__A net1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_44_1662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_131_4309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13004__A net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12546__C net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09162_ ag2.body\[511\] vssd1 vssd1 vccd1 vccd1 _04187_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_25_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13050__A1 net246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10347__B net1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_20_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09093_ ag2.body\[336\] vssd1 vssd1 vccd1 vccd1 _04118_ sky130_fd_sc_hd__inv_2
XFILLER_0_128_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20322_ clknet_leaf_43_clk _01218_ net1378 vssd1 vssd1 vccd1 vccd1 obsg2.randCord\[7\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_86_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold910 control.body\[802\] vssd1 vssd1 vccd1 vccd1 net2472 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16034__B net495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold921 _00596_ vssd1 vssd1 vccd1 vccd1 net2483 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12562__B _07480_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold932 control.body\[817\] vssd1 vssd1 vccd1 vccd1 net2494 sky130_fd_sc_hd__dlygate4sd3_1
X_20253_ clknet_leaf_70_clk _01197_ net1499 vssd1 vssd1 vccd1 vccd1 ag2.body\[139\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_90_3062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold943 _00526_ vssd1 vssd1 vccd1 vccd1 net2505 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17619__A2 net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_3073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold954 control.body\[1002\] vssd1 vssd1 vccd1 vccd1 net2516 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_129_4249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1125_A net1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold965 control.body\[882\] vssd1 vssd1 vccd1 vccd1 net2527 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11364__A1 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11364__B2 net1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold976 control.body\[720\] vssd1 vssd1 vccd1 vccd1 net2538 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11903__A3 _06874_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold987 control.body\[760\] vssd1 vssd1 vccd1 vccd1 net2549 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20184_ clknet_leaf_87_clk _01128_ net1460 vssd1 vssd1 vccd1 vccd1 ag2.body\[214\]
+ sky130_fd_sc_hd__dfrtp_4
Xhold998 _00646_ vssd1 vssd1 vccd1 vccd1 net2560 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09995_ _04603_ _04695_ vssd1 vssd1 vccd1 vccd1 _04968_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout585_A net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13674__A _07181_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14302__A1 net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08946_ net1032 vssd1 vssd1 vccd1 vccd1 _03971_ sky130_fd_sc_hd__inv_2
XANTENNA__14302__B2 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16050__A net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1270 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11116__A1 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11116__B2 net1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_4_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout373_X net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout752_A _04233_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11127__A_N net1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1494_A net1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11194__A net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_3401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15802__A1 ag2.body\[295\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_3412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12616__A1 net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16196__S net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout638_X net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09599__A net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10770_ ag2.body\[223\] net1068 vssd1 vssd1 vccd1 vccd1 _05743_ sky130_fd_sc_hd__xor2_1
XFILLER_0_32_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09429_ net1512 net1506 vssd1 vssd1 vccd1 vccd1 ag2.reset sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_118_3920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout805_X net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_118_3931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12440_ _06635_ _06659_ vssd1 vssd1 vccd1 vccd1 _07401_ sky130_fd_sc_hd__nand2_1
XANTENNA__13041__A1 net254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_871 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_114_3806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_1316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10257__B net1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11052__B1 net763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_1349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16515__C1 net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12371_ net263 net289 vssd1 vssd1 vccd1 vccd1 _07337_ sky130_fd_sc_hd__nor2_1
XFILLER_0_30_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14110_ net1035 ag2.body\[572\] vssd1 vssd1 vccd1 vccd1 _08271_ sky130_fd_sc_hd__nand2_1
X_11322_ ag2.body\[558\] net1077 vssd1 vssd1 vccd1 vccd1 _06295_ sky130_fd_sc_hd__xor2_1
X_15090_ control.body\[925\] net148 _01562_ net2196 vssd1 vssd1 vccd1 vccd1 _00415_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_107_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10544__Y _05517_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_1602 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14041_ _08193_ _08194_ _08196_ _08197_ vssd1 vssd1 vccd1 vccd1 _08202_ sky130_fd_sc_hd__a22o_1
XANTENNA__12147__A3 _07118_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1084 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_535 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12001__C1 net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11253_ _06216_ _06223_ _06224_ _06225_ vssd1 vssd1 vccd1 vccd1 _06226_ sky130_fd_sc_hd__or4_1
XANTENNA__17982__C net39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10158__A2 net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16818__B1 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10204_ _05162_ _05170_ _05176_ _05160_ _05151_ vssd1 vssd1 vccd1 vccd1 _05177_ sky130_fd_sc_hd__o32a_2
XANTENNA__16879__B net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11088__B net1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11184_ ag2.body\[181\] net1105 vssd1 vssd1 vccd1 vccd1 _06157_ sky130_fd_sc_hd__xor2_1
XFILLER_0_105_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17800_ _03469_ _03470_ _03471_ vssd1 vssd1 vccd1 vccd1 _01216_ sky130_fd_sc_hd__and3_1
XANTENNA__17491__B1 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10135_ net1075 control.body\[822\] vssd1 vssd1 vccd1 vccd1 _05108_ sky130_fd_sc_hd__nand2_1
X_15992_ _01673_ _01674_ vssd1 vssd1 vccd1 vccd1 _01675_ sky130_fd_sc_hd__xnor2_1
X_18780_ clknet_leaf_13_clk img_gen.tracker.next_frame\[218\] net1284 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[218\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__18645__CLK clknet_leaf_141_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11107__A1 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14844__A2 _08712_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17731_ _01700_ _01818_ vssd1 vssd1 vccd1 vccd1 _03410_ sky130_fd_sc_hd__nor2_1
X_10066_ net1075 control.body\[718\] vssd1 vssd1 vccd1 vccd1 _05039_ sky130_fd_sc_hd__xor2_1
X_14943_ control.body\[1051\] net174 _01545_ net2217 vssd1 vssd1 vccd1 vccd1 _00285_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12855__A1 net239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11816__B net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_86_2931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17662_ ag2.body\[104\] net887 vssd1 vssd1 vccd1 vccd1 _03341_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_86_2953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14874_ net2125 net182 _01537_ control.body\[1110\] vssd1 vssd1 vccd1 vccd1 _00224_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_134_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10330__A2 net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_2352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19401_ clknet_leaf_102_clk _00345_ net1428 vssd1 vssd1 vccd1 vccd1 control.body\[999\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_67_2363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13825_ _08111_ _08112_ vssd1 vssd1 vccd1 vccd1 _08122_ sky130_fd_sc_hd__nor2_1
X_16613_ obsg2.obstacleArray\[91\] net450 net391 vssd1 vssd1 vccd1 vccd1 _02292_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_82_2828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_2374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17593_ _03269_ _03271_ vssd1 vssd1 vccd1 vccd1 _03272_ sky130_fd_sc_hd__nor2_1
XANTENNA__18795__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_2839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_1044 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_2238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16544_ _02220_ _02221_ vssd1 vssd1 vccd1 vccd1 _02223_ sky130_fd_sc_hd__nand2_1
XFILLER_0_74_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19332_ clknet_leaf_103_clk _00276_ net1431 vssd1 vssd1 vccd1 vccd1 control.body\[1058\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_63_2249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13756_ _08065_ _08072_ _08073_ net320 img_gen.updater.commands.count\[3\] vssd1
+ vssd1 vccd1 vccd1 _00060_ sky130_fd_sc_hd__a32o_1
X_10968_ net1157 control.body\[1003\] vssd1 vssd1 vccd1 vccd1 _05941_ sky130_fd_sc_hd__xnor2_1
XANTENNA__13280__A1 net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16119__B net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12707_ net2049 net647 _07556_ _07557_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[107\]
+ sky130_fd_sc_hd__a31o_1
XANTENNA__11551__B net1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19263_ clknet_leaf_74_clk _00207_ net1495 vssd1 vssd1 vccd1 vccd1 ag2.body\[126\]
+ sky130_fd_sc_hd__dfrtp_4
X_16475_ obsg2.obstacleArray\[43\] _02059_ net397 _02153_ vssd1 vssd1 vccd1 vccd1
+ _02154_ sky130_fd_sc_hd__o211a_1
XFILLER_0_2_1415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11830__A2 net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13687_ _04945_ _08029_ vssd1 vssd1 vccd1 vccd1 _08030_ sky130_fd_sc_hd__and2_2
XFILLER_0_57_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10899_ net1168 control.body\[674\] vssd1 vssd1 vccd1 vccd1 _05872_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_14_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18214_ _03656_ net36 vssd1 vssd1 vccd1 vccd1 _03746_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_14_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15426_ ag2.body\[616\] net84 _01599_ ag2.body\[608\] vssd1 vssd1 vccd1 vccd1 _00714_
+ sky130_fd_sc_hd__a22o_1
X_19194_ clknet_leaf_53_clk _00138_ net1455 vssd1 vssd1 vccd1 vccd1 ag2.body\[57\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_5_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12638_ net295 _07520_ _07521_ net1822 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[74\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__10167__B net1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11043__B1 _06015_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18145_ net529 _03711_ vssd1 vssd1 vccd1 vccd1 _01320_ sky130_fd_sc_hd__and2_1
X_15357_ control.body\[682\] net75 _01592_ net2332 vssd1 vssd1 vccd1 vccd1 _00652_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_87_1573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12663__A net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12569_ net679 _07484_ vssd1 vssd1 vccd1 vccd1 _07485_ sky130_fd_sc_hd__nor2_1
XANTENNA__16135__A net737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1161 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14308_ net1007 ag2.body\[55\] vssd1 vssd1 vccd1 vccd1 _08469_ sky130_fd_sc_hd__nand2_1
XFILLER_0_123_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18076_ net43 _03666_ vssd1 vssd1 vccd1 vccd1 _03667_ sky130_fd_sc_hd__nor2_1
XANTENNA__20373__RESET_B net1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold206 img_gen.tracker.frame\[552\] vssd1 vssd1 vccd1 vccd1 net1768 sky130_fd_sc_hd__dlygate4sd3_1
X_15288_ control.body\[749\] net87 _01584_ control.body\[741\] vssd1 vssd1 vccd1 vccd1
+ _00591_ sky130_fd_sc_hd__a22o_1
Xhold217 img_gen.tracker.frame\[127\] vssd1 vssd1 vccd1 vccd1 net1779 sky130_fd_sc_hd__dlygate4sd3_1
Xhold228 img_gen.tracker.frame\[182\] vssd1 vssd1 vccd1 vccd1 net1790 sky130_fd_sc_hd__dlygate4sd3_1
X_17027_ ag2.body\[403\] net720 net706 ag2.body\[405\] _02705_ vssd1 vssd1 vccd1 vccd1
+ _02706_ sky130_fd_sc_hd__a221o_1
X_14239_ net841 ag2.body\[480\] ag2.body\[486\] net799 vssd1 vssd1 vccd1 vccd1 _08400_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__19420__CLK clknet_leaf_111_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold239 img_gen.tracker.frame\[362\] vssd1 vssd1 vccd1 vccd1 net1801 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16809__B1 net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout708 _04267_ vssd1 vssd1 vccd1 vccd1 net708 sky130_fd_sc_hd__buf_4
XFILLER_0_21_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout719 net721 vssd1 vssd1 vccd1 vccd1 net719 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11897__A2 net596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_4102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17482__B1 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_4113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09691__B net1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09780_ net1060 control.body\[951\] vssd1 vssd1 vccd1 vccd1 _04753_ sky130_fd_sc_hd__xor2_1
XPHY_EDGE_ROW_7_Right_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18978_ clknet_leaf_7_clk img_gen.tracker.next_frame\[416\] net1265 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[416\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_33_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19570__CLK clknet_leaf_118_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_1443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_1620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17929_ net463 net495 vssd1 vssd1 vccd1 vccd1 _03561_ sky130_fd_sc_hd__nor2_1
XFILLER_0_94_1511 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11726__B net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17234__B1 net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1290 net1291 vssd1 vssd1 vccd1 vccd1 net1290 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12627__D_N _07515_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20632__1549 vssd1 vssd1 vccd1 vccd1 _20632__1549/HI net1549 sky130_fd_sc_hd__conb_1
XFILLER_0_90_1419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14599__A1 net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14599__B2 net796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_137_4507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_1724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13271__A1 net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12074__A2 net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_1420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16029__B net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12557__B net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11461__B net1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout333_A _07423_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1075_A net1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09214_ net921 vssd1 vssd1 vccd1 vccd1 _04239_ sky130_fd_sc_hd__inv_2
XFILLER_0_130_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16760__A2 net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_96_3260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09145_ ag2.body\[477\] vssd1 vssd1 vccd1 vccd1 _04170_ sky130_fd_sc_hd__inv_2
XANTENNA__14771__A1 net976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13669__A net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout500_A net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10645__X _05618_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16045__A net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_3124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14771__B2 net1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1242_A net1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout219_X net219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_3135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_945 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09076_ ag2.body\[306\] vssd1 vssd1 vccd1 vccd1 _04101_ sky130_fd_sc_hd__inv_2
XFILLER_0_4_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_1360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16512__A2 _02059_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10805__B net1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20305_ clknet_leaf_37_clk net1575 net1349 vssd1 vssd1 vccd1 vccd1 control.divider.detect.Q\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__20043__RESET_B net1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1030_X net1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold740 control.body\[648\] vssd1 vssd1 vccd1 vccd1 net2302 sky130_fd_sc_hd__dlygate4sd3_1
Xhold751 control.body\[1083\] vssd1 vssd1 vccd1 vccd1 net2313 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1128_X net1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold762 _00248_ vssd1 vssd1 vccd1 vccd1 net2324 sky130_fd_sc_hd__dlygate4sd3_1
Xhold773 _00431_ vssd1 vssd1 vccd1 vccd1 net2335 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20236_ clknet_leaf_65_clk _01180_ net1496 vssd1 vssd1 vccd1 vccd1 ag2.body\[154\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA_fanout490_X net490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17699__S1 net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold784 control.body\[780\] vssd1 vssd1 vccd1 vccd1 net2346 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11888__A2 net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold795 _00688_ vssd1 vssd1 vccd1 vccd1 net2357 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout967_A net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16276__A1 net372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1433 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout588_X net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20167_ clknet_leaf_95_clk _01111_ net1441 vssd1 vssd1 vccd1 vccd1 ag2.body\[229\]
+ sky130_fd_sc_hd__dfrtp_4
X_09978_ net1183 control.body\[1114\] vssd1 vssd1 vccd1 vccd1 _04951_ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout79_A net91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20098_ clknet_leaf_79_clk _01042_ net1489 vssd1 vssd1 vccd1 vccd1 ag2.body\[288\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__12837__A1 net239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout755_X net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10540__B net1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17225__B1 net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11940_ img_gen.tracker.frame\[160\] net603 net580 img_gen.tracker.frame\[166\] vssd1
+ vssd1 vccd1 vccd1 _06912_ sky130_fd_sc_hd__o22a_1
X_20608__1540 vssd1 vssd1 vccd1 vccd1 _20608__1540/HI net1540 sky130_fd_sc_hd__conb_1
XANTENNA__16579__A2 net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout922_X net922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11871_ img_gen.tracker.frame\[283\] net548 _06841_ _06842_ vssd1 vssd1 vccd1 vccd1
+ _06843_ sky130_fd_sc_hd__o211a_1
X_13610_ _07957_ net220 _07982_ vssd1 vssd1 vccd1 vccd1 control.divider.next_count\[2\]
+ sky130_fd_sc_hd__and3_1
XANTENNA__11652__A net1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10822_ control.body\[1088\] net1231 vssd1 vssd1 vccd1 vccd1 _05795_ sky130_fd_sc_hd__and2b_1
X_14590_ net815 ag2.body\[84\] _04015_ net1013 vssd1 vssd1 vccd1 vccd1 _08751_ sky130_fd_sc_hd__o22a_1
XANTENNA__13262__A1 net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09466__B1 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12467__B _07306_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11371__B net1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13541_ net1939 net656 _07927_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[571\]
+ sky130_fd_sc_hd__and3_1
XFILLER_0_95_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10753_ net1202 control.body\[889\] vssd1 vssd1 vccd1 vccd1 _05726_ sky130_fd_sc_hd__xor2_1
XFILLER_0_95_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19226__RESET_B net1482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16260_ obsg2.obstacleArray\[54\] obsg2.obstacleArray\[55\] net407 vssd1 vssd1 vccd1
+ vccd1 _01939_ sky130_fd_sc_hd__mux2_1
X_13472_ net230 _07900_ _07901_ net1655 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[528\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_109_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10684_ _04433_ _04695_ _04419_ vssd1 vssd1 vccd1 vccd1 _05657_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_124_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15211_ net2182 net92 _01575_ control.body\[801\] vssd1 vssd1 vccd1 vccd1 _00523_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_35_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12423_ net743 _07384_ vssd1 vssd1 vccd1 vccd1 _07385_ sky130_fd_sc_hd__xnor2_1
X_16191_ _01743_ _01869_ _01862_ _01729_ vssd1 vssd1 vccd1 vccd1 _01870_ sky130_fd_sc_hd__a211o_1
XANTENNA__14762__A1 net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12483__A net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11576__A1 net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_2610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_2621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15142_ control.body\[876\] net106 _01567_ net2254 vssd1 vssd1 vccd1 vccd1 _00462_
+ sky130_fd_sc_hd__a22o_1
X_12354_ img_gen.updater.commands.rR1.rainbowRNG\[0\] net248 vssd1 vssd1 vccd1 vccd1
+ _07321_ sky130_fd_sc_hd__and2_1
XFILLER_0_106_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_56_2020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_2031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10715__B net1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20420__CLK clknet_leaf_37_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_2042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11305_ ag2.body\[279\] net1066 vssd1 vssd1 vccd1 vccd1 _06278_ sky130_fd_sc_hd__xor2_1
X_19950_ clknet_leaf_45_clk _00894_ net1379 vssd1 vssd1 vccd1 vccd1 ag2.body\[444\]
+ sky130_fd_sc_hd__dfrtp_4
X_15073_ control.body\[942\] net149 _01560_ net2409 vssd1 vssd1 vccd1 vccd1 _00400_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_50_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15711__B1 _01629_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12285_ _07251_ _07253_ vssd1 vssd1 vccd1 vccd1 _07255_ sky130_fd_sc_hd__nand2_2
X_14024_ net980 ag2.body\[26\] vssd1 vssd1 vccd1 vccd1 _08185_ sky130_fd_sc_hd__xnor2_1
X_18901_ clknet_leaf_144_clk img_gen.tracker.next_frame\[339\] net1251 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[339\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__13868__A3 _08141_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_1488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11236_ ag2.body\[194\] net1177 vssd1 vssd1 vccd1 vccd1 _06209_ sky130_fd_sc_hd__or2_1
X_19881_ clknet_leaf_82_clk _00825_ net1479 vssd1 vssd1 vccd1 vccd1 ag2.body\[519\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__11879__A2 net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16267__A1 net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18832_ clknet_leaf_4_clk img_gen.tracker.next_frame\[270\] net1260 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[270\] sky130_fd_sc_hd__dfrtp_1
X_11167_ net1130 control.body\[780\] vssd1 vssd1 vccd1 vccd1 _06140_ sky130_fd_sc_hd__nand2_1
XANTENNA__14203__A net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10118_ net1096 control.body\[709\] vssd1 vssd1 vccd1 vccd1 _05091_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_69_2414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18763_ clknet_leaf_16_clk img_gen.tracker.next_frame\[201\] net1314 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[201\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__12568__A_N net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_2425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11098_ ag2.body\[425\] net1199 vssd1 vssd1 vccd1 vccd1 _06071_ sky130_fd_sc_hd__xnor2_1
X_15975_ _08118_ net56 vssd1 vssd1 vccd1 vccd1 _01661_ sky130_fd_sc_hd__nor2_1
XANTENNA__10450__B net1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_2436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17714_ net360 net357 _03392_ _03391_ vssd1 vssd1 vccd1 vccd1 _03393_ sky130_fd_sc_hd__a31o_1
XFILLER_0_89_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10839__B1 _05798_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14926_ control.body\[1068\] net170 _01543_ net2351 vssd1 vssd1 vccd1 vccd1 _00270_
+ sky130_fd_sc_hd__a22o_1
X_10049_ _05008_ _05009_ _05010_ _05021_ vssd1 vssd1 vccd1 vccd1 _05022_ sky130_fd_sc_hd__o31a_1
XFILLER_0_117_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18694_ clknet_leaf_11_clk img_gen.tracker.next_frame\[132\] net1281 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[132\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_72_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17645_ ag2.body\[33\] net868 vssd1 vssd1 vccd1 vccd1 _03324_ sky130_fd_sc_hd__xnor2_1
X_14857_ _08200_ _08204_ _08437_ _08499_ _08722_ vssd1 vssd1 vccd1 vccd1 _01528_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_72_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17782__A4 net974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13808_ _08107_ _08108_ _07410_ vssd1 vssd1 vccd1 vccd1 _00077_ sky130_fd_sc_hd__a21boi_1
X_17576_ ag2.body\[342\] net945 vssd1 vssd1 vccd1 vccd1 _03255_ sky130_fd_sc_hd__xor2_1
XFILLER_0_86_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12056__A2 net555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14788_ _01457_ _01458_ vssd1 vssd1 vccd1 vccd1 _01459_ sky130_fd_sc_hd__nand2_1
XFILLER_0_58_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09457__B1 _04429_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16990__A2 net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19315_ clknet_leaf_104_clk net2294 net1433 vssd1 vssd1 vccd1 vccd1 control.body\[1073\]
+ sky130_fd_sc_hd__dfrtp_1
X_16527_ net433 _02205_ vssd1 vssd1 vccd1 vccd1 _02206_ sky130_fd_sc_hd__nor2_2
XFILLER_0_85_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13739_ _07187_ _07209_ _08057_ _08059_ vssd1 vssd1 vccd1 vccd1 _08060_ sky130_fd_sc_hd__a31o_1
XFILLER_0_86_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_988 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19246_ clknet_leaf_76_clk _00190_ net1482 vssd1 vssd1 vccd1 vccd1 ag2.body\[109\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__13005__A1 net240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16458_ net364 _02123_ _02127_ net363 vssd1 vssd1 vccd1 vccd1 _02137_ sky130_fd_sc_hd__o211ai_1
XANTENNA__16742__A2 net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15409_ net2638 net81 _01597_ control.body\[625\] vssd1 vssd1 vccd1 vccd1 _00699_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_115_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16389_ _02065_ _02066_ vssd1 vssd1 vccd1 vccd1 _02068_ sky130_fd_sc_hd__or2_1
XANTENNA__09686__B net1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19177_ clknet_leaf_20_clk _00121_ net1365 vssd1 vssd1 vccd1 vccd1 ag2.body\[40\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_14_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10906__A net1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_83_clk_A clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11567__A1 net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18128_ obsg2.obstacleArray\[63\] _03700_ net524 vssd1 vssd1 vccd1 vccd1 _01314_
+ sky130_fd_sc_hd__o21a_1
XANTENNA__14505__A1 net981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14505__B2 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18059_ obsg2.obstacleArray\[39\] _03655_ net522 vssd1 vssd1 vccd1 vccd1 _01290_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_112_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09901_ ag2.body\[75\] net1163 vssd1 vssd1 vccd1 vccd1 _04874_ sky130_fd_sc_hd__xor2_1
XFILLER_0_10_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_35_1403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_98_clk_A clknet_4_11__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16258__A1 net417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout505 _06468_ vssd1 vssd1 vccd1 vccd1 net505 sky130_fd_sc_hd__buf_4
X_20021_ clknet_leaf_58_clk _00965_ net1471 vssd1 vssd1 vccd1 vccd1 ag2.body\[371\]
+ sky130_fd_sc_hd__dfrtp_4
Xfanout516 net517 vssd1 vssd1 vccd1 vccd1 net516 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_6_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout527 net528 vssd1 vssd1 vccd1 vccd1 net527 sky130_fd_sc_hd__clkbuf_4
X_09832_ _04801_ _04802_ _04803_ _04804_ vssd1 vssd1 vccd1 vccd1 _04805_ sky130_fd_sc_hd__a22o_1
Xfanout538 _01707_ vssd1 vssd1 vccd1 vccd1 net538 sky130_fd_sc_hd__clkbuf_4
XANTENNA__15209__A _06331_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12531__A3 _07444_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_141_clk_A clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14113__A net1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout549 net550 vssd1 vssd1 vccd1 vccd1 net549 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09207__A net1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09763_ ag2.body\[210\] net1184 vssd1 vssd1 vccd1 vccd1 _04736_ sky130_fd_sc_hd__xor2_1
XANTENNA__11456__B net1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12819__A1 net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout283_A net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_21_clk_A clknet_4_6__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09694_ ag2.body\[71\] net1064 vssd1 vssd1 vccd1 vccd1 _04667_ sky130_fd_sc_hd__nand2_1
XANTENNA__13492__A1 net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17758__A1 net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout450_A net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_29_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1192_A net1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout548_A net550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20558__Q net25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1601 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09213__Y _04238_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12047__A2 net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13244__A1 net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_36_clk_A clknet_4_5__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16981__A2 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_3300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_3311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_98_3322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout715_A net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17797__C net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_385 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1078_X net1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09877__A ag2.body\[165\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16194__B1 net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16733__A2 net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout503_X net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10816__A net1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09128_ ag2.body\[430\] vssd1 vssd1 vccd1 vccd1 _04153_ sky130_fd_sc_hd__inv_2
XANTENNA__16497__A1 net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17694__B1 net963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17158__X _02837_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_855 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09059_ ag2.body\[254\] vssd1 vssd1 vccd1 vccd1 _04084_ sky130_fd_sc_hd__inv_2
X_12070_ img_gen.tracker.frame\[114\] net556 _07041_ net561 vssd1 vssd1 vccd1 vccd1
+ _07042_ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout872_X net872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17318__B net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold570 img_gen.tracker.frame\[574\] vssd1 vssd1 vccd1 vccd1 net2132 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12750__B _07578_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold581 control.body\[1119\] vssd1 vssd1 vccd1 vccd1 net2143 sky130_fd_sc_hd__dlygate4sd3_1
Xhold592 control.body\[907\] vssd1 vssd1 vccd1 vccd1 net2154 sky130_fd_sc_hd__dlygate4sd3_1
X_11021_ ag2.body\[597\] net1098 vssd1 vssd1 vccd1 vccd1 _05994_ sky130_fd_sc_hd__nand2_1
X_20219_ clknet_leaf_60_clk _01163_ net1466 vssd1 vssd1 vccd1 vccd1 ag2.body\[169\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA_clkbuf_leaf_109_clk_A clknet_4_10__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14023__A net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10270__B net1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16649__S net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15760_ ag2.body\[321\] net216 _01636_ ag2.body\[313\] vssd1 vssd1 vccd1 vccd1 _01011_
+ sky130_fd_sc_hd__a22o_1
X_12972_ img_gen.tracker.frame\[247\] net645 vssd1 vssd1 vccd1 vccd1 _07683_ sky130_fd_sc_hd__and2_1
XANTENNA__13483__A1 net250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12749__Y _07578_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14711_ net985 ag2.body\[338\] vssd1 vssd1 vccd1 vccd1 _08872_ sky130_fd_sc_hd__xor2_1
X_11923_ img_gen.tracker.frame\[304\] net606 vssd1 vssd1 vccd1 vccd1 _06895_ sky130_fd_sc_hd__nor2_1
X_15691_ ag2.body\[389\] net140 _01616_ ag2.body\[381\] vssd1 vssd1 vccd1 vccd1 _00951_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__19809__CLK clknet_leaf_124_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11382__A net1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16421__B2 net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17430_ _03106_ _03107_ _03108_ vssd1 vssd1 vccd1 vccd1 _03109_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_16_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12909__C _07315_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14642_ net1021 ag2.body\[518\] vssd1 vssd1 vccd1 vccd1 _08803_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_16_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11854_ img_gen.tracker.frame\[226\] net590 net552 img_gen.tracker.frame\[223\] vssd1
+ vssd1 vccd1 vccd1 _06826_ sky130_fd_sc_hd__o22a_1
XFILLER_0_135_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_16_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16972__A2 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16892__B net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10805_ ag2.body\[33\] net1197 vssd1 vssd1 vccd1 vccd1 _05778_ sky130_fd_sc_hd__xor2_1
X_17361_ _03010_ _03013_ vssd1 vssd1 vccd1 vccd1 _03040_ sky130_fd_sc_hd__nand2_1
X_14573_ net828 ag2.body\[490\] _04178_ net1039 _08733_ vssd1 vssd1 vccd1 vccd1 _08734_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_36_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11785_ img_gen.tracker.frame\[338\] net615 net598 img_gen.tracker.frame\[341\] vssd1
+ vssd1 vccd1 vccd1 _06757_ sky130_fd_sc_hd__o22a_1
XFILLER_0_28_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18165__A net518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11797__A1 net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19100_ clknet_leaf_0_clk img_gen.tracker.next_frame\[538\] net1239 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[538\] sky130_fd_sc_hd__dfrtp_1
X_16312_ obsg2.obstacleArray\[110\] obsg2.obstacleArray\[111\] net405 vssd1 vssd1
+ vccd1 vccd1 _01991_ sky130_fd_sc_hd__mux2_1
XANTENNA__09787__A net1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13524_ _07621_ _07807_ vssd1 vssd1 vccd1 vccd1 _07921_ sky130_fd_sc_hd__or2_1
XFILLER_0_126_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17292_ _02962_ _02963_ _02964_ _02967_ vssd1 vssd1 vccd1 vccd1 _02971_ sky130_fd_sc_hd__or4_1
XANTENNA__18833__CLK clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10736_ ag2.body\[253\] net756 net746 ag2.body\[255\] _05701_ vssd1 vssd1 vccd1 vccd1
+ _05709_ sky130_fd_sc_hd__o221a_1
XFILLER_0_126_936 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11892__S1 net1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16243_ _01920_ _01921_ net415 vssd1 vssd1 vccd1 vccd1 _01922_ sky130_fd_sc_hd__mux2_1
X_19031_ clknet_leaf_6_clk img_gen.tracker.next_frame\[469\] net1265 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[469\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13455_ _07584_ net302 vssd1 vssd1 vccd1 vccd1 _07894_ sky130_fd_sc_hd__nor2_1
X_10667_ net785 control.body\[880\] control.body\[886\] net751 _05638_ vssd1 vssd1
+ vccd1 vccd1 _05640_ sky130_fd_sc_hd__a221o_1
XFILLER_0_24_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_2104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12406_ net1167 net610 vssd1 vssd1 vccd1 vccd1 _07369_ sky130_fd_sc_hd__nand2_1
X_16174_ net348 _01852_ _01849_ _01742_ vssd1 vssd1 vccd1 vccd1 _01853_ sky130_fd_sc_hd__o211a_1
X_13386_ net274 _07866_ _07867_ net2134 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[476\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_84_1554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10598_ _05562_ _05565_ _05566_ _05569_ vssd1 vssd1 vccd1 vccd1 _05571_ sky130_fd_sc_hd__or4_1
X_20631__1548 vssd1 vssd1 vccd1 vccd1 _20631__1548/HI net1548 sky130_fd_sc_hd__conb_1
XANTENNA__16488__A1 net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15125_ control.body\[893\] net104 _01565_ net2328 vssd1 vssd1 vccd1 vccd1 _00447_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_105_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17685__B1 net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12337_ _07301_ _07173_ _06634_ vssd1 vssd1 vccd1 vccd1 _07304_ sky130_fd_sc_hd__or3b_2
XANTENNA__18983__CLK clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12941__A net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19933_ clknet_leaf_47_clk _00877_ net1375 vssd1 vssd1 vccd1 vccd1 ag2.body\[459\]
+ sky130_fd_sc_hd__dfrtp_4
X_15056_ net2220 net163 _01558_ control.body\[951\] vssd1 vssd1 vccd1 vccd1 _00385_
+ sky130_fd_sc_hd__a22o_1
X_12268_ _07234_ _07235_ _07237_ vssd1 vssd1 vccd1 vccd1 _07238_ sky130_fd_sc_hd__a21oi_1
XANTENNA__17437__B1 net693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14007_ net1021 ag2.body\[510\] vssd1 vssd1 vccd1 vccd1 _08168_ sky130_fd_sc_hd__or2_1
XFILLER_0_120_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11219_ _06188_ _06189_ _06190_ _06191_ vssd1 vssd1 vccd1 vccd1 _06192_ sky130_fd_sc_hd__and4_1
X_19864_ clknet_leaf_94_clk _00808_ net1437 vssd1 vssd1 vccd1 vccd1 ag2.body\[534\]
+ sky130_fd_sc_hd__dfrtp_4
X_12199_ net317 _07169_ vssd1 vssd1 vccd1 vccd1 _07171_ sky130_fd_sc_hd__and2_1
XANTENNA__11276__B net1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18815_ clknet_leaf_4_clk img_gen.tracker.next_frame\[253\] net1249 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[253\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__10180__B net1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19795_ clknet_leaf_124_clk _00739_ net1328 vssd1 vssd1 vccd1 vccd1 ag2.body\[593\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__15463__A2 net90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18746_ clknet_leaf_139_clk img_gen.tracker.next_frame\[184\] net1256 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[184\] sky130_fd_sc_hd__dfrtp_1
X_15958_ ag2.body\[146\] net199 _01657_ ag2.body\[138\] vssd1 vssd1 vccd1 vccd1 _01188_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_95_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13474__A1 net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14909_ net2253 net177 _01541_ control.body\[1077\] vssd1 vssd1 vccd1 vccd1 _00255_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_77_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18677_ clknet_leaf_27_clk img_gen.tracker.next_frame\[115\] net1339 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[115\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_76_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15889_ ag2.body\[213\] net184 _01649_ ag2.body\[205\] vssd1 vssd1 vccd1 vccd1 _01127_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_91_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17628_ ag2.body\[188\] net714 net697 ag2.body\[190\] vssd1 vssd1 vccd1 vccd1 _03307_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_56_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17898__B _03531_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10179__Y _05152_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17559_ ag2.body\[354\] net728 net935 _04128_ _03237_ vssd1 vssd1 vccd1 vccd1 _03238_
+ sky130_fd_sc_hd__a221o_1
XANTENNA__16294__S net419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_897 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18075__A net301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20570_ clknet_leaf_107_clk _01428_ _00034_ vssd1 vssd1 vccd1 vccd1 sound_gen.dac1.dacCount\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__16715__A2 net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19229_ clknet_leaf_85_clk _00173_ net1483 vssd1 vssd1 vccd1 vccd1 ag2.body\[92\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__10636__A net1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14108__A net997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout129_A net132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1016 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10355__B net1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1004 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1184 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1038_A net1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17138__B net933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16042__B net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_1396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout498_A net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout302 net303 vssd1 vssd1 vccd1 vccd1 net302 sky130_fd_sc_hd__buf_2
XANTENNA_clkbuf_4_7__f_clk_X clknet_4_7__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17428__B1 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09208__Y _04233_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout313 net314 vssd1 vssd1 vccd1 vccd1 net313 sky130_fd_sc_hd__buf_1
Xfanout324 track.nextHighScore\[4\] vssd1 vssd1 vccd1 vccd1 net324 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_61_1384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1205_A net1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout335 _07423_ vssd1 vssd1 vccd1 vccd1 net335 sky130_fd_sc_hd__clkbuf_2
Xfanout346 _01732_ vssd1 vssd1 vccd1 vccd1 net346 sky130_fd_sc_hd__clkbuf_4
XANTENNA_input3_A gpio_in[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16977__B net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20004_ clknet_leaf_61_clk _00948_ net1468 vssd1 vssd1 vccd1 vccd1 ag2.body\[386\]
+ sky130_fd_sc_hd__dfrtp_4
X_09815_ net1160 _04253_ control.body\[1052\] net761 _04787_ vssd1 vssd1 vccd1 vccd1
+ _04788_ sky130_fd_sc_hd__o221a_1
Xfanout379 _01739_ vssd1 vssd1 vccd1 vccd1 net379 sky130_fd_sc_hd__buf_2
XANTENNA__18706__CLK clknet_leaf_144_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout286_X net286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout665_A net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16651__A1 obsg2.obstacleArray\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09746_ net907 _04718_ vssd1 vssd1 vccd1 vccd1 _04719_ sky130_fd_sc_hd__nor2_2
XFILLER_0_74_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09677_ ag2.body\[10\] net1175 vssd1 vssd1 vccd1 vccd1 _04650_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout453_X net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout832_A net836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1195_X net1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11571__S0 net1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_96_447 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13217__A1 net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__20405__RESET_B net1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout620_X net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1362_X net1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout718_X net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11930__A net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11570_ net506 _06542_ vssd1 vssd1 vccd1 vccd1 _06543_ sky130_fd_sc_hd__or2_1
XFILLER_0_33_1486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16706__A2 net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10521_ _05490_ _05491_ _05492_ _05493_ vssd1 vssd1 vccd1 vccd1 _05494_ sky130_fd_sc_hd__and4_1
XANTENNA__15914__B1 _01652_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13240_ net259 _07808_ _07809_ net1940 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[388\]
+ sky130_fd_sc_hd__a22o_1
X_10452_ ag2.body\[454\] net1079 vssd1 vssd1 vccd1 vccd1 _05425_ sky130_fd_sc_hd__or2_1
XFILLER_0_81_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10265__B net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13171_ img_gen.tracker.frame\[352\] net644 vssd1 vssd1 vccd1 vccd1 _07777_ sky130_fd_sc_hd__and2_1
X_10383_ ag2.body\[108\] net1140 vssd1 vssd1 vccd1 vccd1 _05356_ sky130_fd_sc_hd__xor2_1
XANTENNA__16233__A net460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12122_ img_gen.tracker.frame\[543\] net596 vssd1 vssd1 vccd1 vccd1 _07094_ sky130_fd_sc_hd__or2_1
XFILLER_0_32_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16930_ _04131_ net872 net717 ag2.body\[371\] _02608_ vssd1 vssd1 vccd1 vccd1 _02609_
+ sky130_fd_sc_hd__o221a_1
X_12053_ _06690_ _07024_ vssd1 vssd1 vccd1 vccd1 _07025_ sky130_fd_sc_hd__nor2_1
XANTENNA__20339__CLK clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16520__X _02199_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11004_ net755 control.body\[1085\] control.body\[1087\] net745 _05976_ vssd1 vssd1
+ vccd1 vccd1 _05977_ sky130_fd_sc_hd__o221a_1
XANTENNA__11096__B net1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16861_ _04062_ net886 net943 _04066_ _02539_ vssd1 vssd1 vccd1 vccd1 _02540_ sky130_fd_sc_hd__a221o_1
XANTENNA__10911__C1 _05869_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16642__A1 net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout880 net881 vssd1 vssd1 vccd1 vccd1 net880 sky130_fd_sc_hd__buf_2
X_18600_ clknet_leaf_17_clk img_gen.tracker.next_frame\[38\] net1318 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[38\] sky130_fd_sc_hd__dfrtp_1
Xfanout891 net894 vssd1 vssd1 vccd1 vccd1 net891 sky130_fd_sc_hd__buf_4
X_15812_ _04985_ net66 vssd1 vssd1 vccd1 vccd1 _01642_ sky130_fd_sc_hd__and2_2
X_19580_ clknet_leaf_118_clk _00524_ net1386 vssd1 vssd1 vccd1 vccd1 control.body\[810\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_3_6_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_3_6_0_clk sky130_fd_sc_hd__clkbuf_8
X_16792_ net402 _02470_ vssd1 vssd1 vccd1 vccd1 _02471_ sky130_fd_sc_hd__or2_1
XFILLER_0_88_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18531_ clknet_leaf_137_clk _00057_ net1298 vssd1 vssd1 vccd1 vccd1 img_gen.updater.commands.count\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__20489__CLK clknet_leaf_37_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15743_ ag2.body\[338\] net217 _01634_ ag2.body\[330\] vssd1 vssd1 vccd1 vccd1 _00996_
+ sky130_fd_sc_hd__a22o_1
X_12955_ img_gen.tracker.frame\[238\] net660 vssd1 vssd1 vccd1 vccd1 _07675_ sky130_fd_sc_hd__and2_1
XANTENNA__14804__A1_N net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11906_ img_gen.tracker.frame\[361\] net622 net588 img_gen.tracker.frame\[370\] vssd1
+ vssd1 vccd1 vccd1 _06878_ sky130_fd_sc_hd__o22a_1
XANTENNA__12639__C net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18462_ net717 _01687_ vssd1 vssd1 vccd1 vccd1 _03950_ sky130_fd_sc_hd__or2_1
XFILLER_0_90_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15674_ ag2.body\[405\] net142 _01626_ ag2.body\[397\] vssd1 vssd1 vccd1 vccd1 _00935_
+ sky130_fd_sc_hd__a22o_1
X_12886_ _07439_ _07639_ vssd1 vssd1 vccd1 vccd1 _07643_ sky130_fd_sc_hd__nor2_1
XANTENNA__19781__CLK clknet_leaf_127_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17413_ ag2.body\[282\] net727 net699 ag2.body\[286\] _03089_ vssd1 vssd1 vccd1 vccd1
+ _03092_ sky130_fd_sc_hd__o221ai_1
XFILLER_0_96_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14625_ net972 ag2.body\[467\] vssd1 vssd1 vccd1 vccd1 _08786_ sky130_fd_sc_hd__xor2_1
X_11837_ img_gen.tracker.frame\[563\] net587 net550 img_gen.tracker.frame\[560\] _06808_
+ vssd1 vssd1 vccd1 vccd1 _06809_ sky130_fd_sc_hd__o221a_1
XANTENNA__17511__B net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18393_ _03815_ _03872_ _03880_ _03881_ _03882_ vssd1 vssd1 vccd1 vccd1 _03883_ sky130_fd_sc_hd__o221a_1
XFILLER_0_68_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17344_ _03022_ vssd1 vssd1 vccd1 vccd1 _03023_ sky130_fd_sc_hd__inv_2
X_14556_ _08713_ _08714_ _08716_ vssd1 vssd1 vccd1 vccd1 _08717_ sky130_fd_sc_hd__or3b_1
XFILLER_0_3_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11768_ img_gen.tracker.frame\[59\] net580 net542 img_gen.tracker.frame\[56\] _06739_
+ vssd1 vssd1 vccd1 vccd1 _06740_ sky130_fd_sc_hd__o221a_1
XFILLER_0_56_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_99_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13507_ net230 _07914_ _07915_ net1843 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[549\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__14708__A1 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10719_ _04224_ net1120 net753 ag2.body\[621\] _05687_ vssd1 vssd1 vccd1 vccd1 _05692_
+ sky130_fd_sc_hd__a221o_1
X_14487_ net993 ag2.body\[345\] vssd1 vssd1 vccd1 vccd1 _08648_ sky130_fd_sc_hd__xor2_1
XFILLER_0_83_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14708__B2 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17275_ ag2.body\[552\] net881 vssd1 vssd1 vccd1 vccd1 _02954_ sky130_fd_sc_hd__xor2_1
XFILLER_0_86_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11699_ _06642_ _06670_ vssd1 vssd1 vccd1 vccd1 _06671_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_71_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19014_ clknet_leaf_1_clk img_gen.tracker.next_frame\[452\] net1246 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[452\] sky130_fd_sc_hd__dfrtp_1
X_16226_ net495 _01897_ vssd1 vssd1 vccd1 vccd1 _01905_ sky130_fd_sc_hd__and2_2
X_13438_ net256 _07886_ _07887_ net2021 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[508\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_113_416 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1325 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10175__B net1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16157_ _01742_ _01831_ _01835_ _01729_ vssd1 vssd1 vccd1 vccd1 _01836_ sky130_fd_sc_hd__a31o_1
X_13369_ net1765 _07861_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[465\]
+ sky130_fd_sc_hd__and2_1
XANTENNA__19161__CLK clknet_leaf_52_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15108_ control.body\[909\] net146 _01564_ net2334 vssd1 vssd1 vccd1 vccd1 _00431_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_2_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16088_ net348 _01766_ _01763_ _01743_ vssd1 vssd1 vccd1 vccd1 _01767_ sky130_fd_sc_hd__o211a_1
XANTENNA__13486__B net644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18729__CLK clknet_leaf_142_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11287__A net1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19916_ clknet_leaf_55_clk _00860_ net1456 vssd1 vssd1 vccd1 vccd1 ag2.body\[474\]
+ sky130_fd_sc_hd__dfrtp_4
X_15039_ control.body\[975\] net165 _01557_ control.body\[967\] vssd1 vssd1 vccd1
+ vccd1 _00369_ sky130_fd_sc_hd__a22o_1
XFILLER_0_20_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09899__B1 net1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18083__B1 net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19847_ clknet_leaf_92_clk _00791_ net1412 vssd1 vssd1 vccd1 vccd1 ag2.body\[549\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__16289__S net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16633__A1 net395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09600_ net643 _04571_ vssd1 vssd1 vccd1 vccd1 _04573_ sky130_fd_sc_hd__nand2_4
XANTENNA__13447__A1 net235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19778_ clknet_leaf_19_clk _00722_ net1331 vssd1 vssd1 vccd1 vccd1 ag2.body\[608\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__14644__B1 net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09531_ net1085 control.body\[1030\] vssd1 vssd1 vccd1 vccd1 _04504_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_56_1420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18729_ clknet_leaf_142_clk img_gen.tracker.next_frame\[167\] net1253 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[167\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_64_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17189__A2 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09462_ ag2.body\[383\] net1056 vssd1 vssd1 vccd1 vccd1 _04435_ sky130_fd_sc_hd__xor2_1
XANTENNA__10728__A_N net1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09393_ _04346_ _04380_ vssd1 vssd1 vccd1 vccd1 _01406_ sky130_fd_sc_hd__nor2_1
XANTENNA__18138__A1 net48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12846__A net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout246_A net247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11750__A net1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20622_ img_gen.dcx vssd1 vssd1 vccd1 vccd1 net33 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20553_ clknet_leaf_106_clk _01418_ _00027_ vssd1 vssd1 vccd1 vccd1 sound_gen.osc1.stayCount\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10366__A net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1155_A net1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19504__CLK clknet_leaf_113_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20484_ clknet_leaf_37_clk _01371_ net1353 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[120\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_67_1560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18252__B net35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09874__B net1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12581__A net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17113__A2 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10736__A2 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_110_3672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_41_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_110_3683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1110_X net1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1108 net1109 vssd1 vssd1 vccd1 vccd1 net1108 sky130_fd_sc_hd__buf_4
Xfanout110 net112 vssd1 vssd1 vccd1 vccd1 net110 sky130_fd_sc_hd__clkbuf_2
Xfanout121 net128 vssd1 vssd1 vccd1 vccd1 net121 sky130_fd_sc_hd__buf_2
Xfanout1119 net1121 vssd1 vssd1 vccd1 vccd1 net1119 sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout1208_X net1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout132 net144 vssd1 vssd1 vccd1 vccd1 net132 sky130_fd_sc_hd__clkbuf_2
Xclkbuf_4_1__f_clk clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_1__leaf_clk sky130_fd_sc_hd__clkbuf_16
XANTENNA__09890__A net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout143 net144 vssd1 vssd1 vccd1 vccd1 net143 sky130_fd_sc_hd__buf_2
Xfanout154 net183 vssd1 vssd1 vccd1 vccd1 net154 sky130_fd_sc_hd__buf_2
Xfanout165 net171 vssd1 vssd1 vccd1 vccd1 net165 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout668_X net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout176 net183 vssd1 vssd1 vccd1 vccd1 net176 sky130_fd_sc_hd__clkbuf_2
Xfanout187 net218 vssd1 vssd1 vccd1 vccd1 net187 sky130_fd_sc_hd__clkbuf_2
XANTENNA__11503__A_N net1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14939__C net65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout198 net199 vssd1 vssd1 vccd1 vccd1 net198 sky130_fd_sc_hd__buf_2
XANTENNA__13438__A1 net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout61_A net62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09729_ ag2.body\[92\] net1140 vssd1 vssd1 vccd1 vccd1 _04702_ sky130_fd_sc_hd__or2_1
XFILLER_0_74_1520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout835_X net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12740_ net237 _07573_ _07574_ net1698 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[123\]
+ sky130_fd_sc_hd__a22o_1
X_20630__1547 vssd1 vssd1 vccd1 vccd1 _20630__1547/HI net1547 sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_104_3487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_3498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16927__A2 net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17331__B net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12671_ net242 _07540_ _07541_ net2137 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[87\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12756__A net305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14410_ net1016 net924 vssd1 vssd1 vccd1 vccd1 _08571_ sky130_fd_sc_hd__or2_1
XFILLER_0_93_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11622_ net759 _06593_ _06594_ _06485_ _06591_ vssd1 vssd1 vccd1 vccd1 _06595_ sky130_fd_sc_hd__o311a_1
XFILLER_0_93_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15390_ _05857_ net63 vssd1 vssd1 vccd1 vccd1 _01596_ sky130_fd_sc_hd__and2_2
XANTENNA__12475__B net315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11847__S1 net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10424__A1 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14341_ net987 ag2.body\[609\] vssd1 vssd1 vccd1 vccd1 _08502_ sky130_fd_sc_hd__xor2_1
XANTENNA__10424__B2 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17888__B1 _03521_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11553_ net1174 _06522_ _06504_ vssd1 vssd1 vccd1 vccd1 _06526_ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19184__CLK clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17060_ _04005_ net865 net693 ag2.body\[79\] vssd1 vssd1 vccd1 vccd1 _02739_ sky130_fd_sc_hd__o22a_1
X_10504_ net1181 control.body\[978\] vssd1 vssd1 vccd1 vccd1 _05477_ sky130_fd_sc_hd__xor2_1
X_14272_ net1008 ag2.body\[15\] vssd1 vssd1 vccd1 vccd1 _08433_ sky130_fd_sc_hd__or2_1
XFILLER_0_123_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11484_ _06122_ _06239_ _06343_ _06456_ vssd1 vssd1 vccd1 vccd1 _06457_ sky130_fd_sc_hd__and4b_1
X_16011_ net732 _01685_ vssd1 vssd1 vccd1 vccd1 _01690_ sky130_fd_sc_hd__or2_1
XANTENNA__18162__B net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12177__A1 net317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13223_ _07801_ net263 _07799_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[379\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10435_ net1063 control.body\[935\] vssd1 vssd1 vccd1 vccd1 _05408_ sky130_fd_sc_hd__and2_1
XANTENNA__12491__A _07431_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10188__B1 net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11033__A_N net1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13154_ img_gen.tracker.frame\[343\] net644 vssd1 vssd1 vccd1 vccd1 _07769_ sky130_fd_sc_hd__and2_1
XFILLER_0_46_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10366_ net1052 control.body\[767\] vssd1 vssd1 vccd1 vccd1 _05339_ sky130_fd_sc_hd__xor2_1
XFILLER_0_42_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12105_ net564 _07073_ _07076_ vssd1 vssd1 vccd1 vccd1 _07077_ sky130_fd_sc_hd__o21a_1
X_17962_ net47 net296 _03586_ vssd1 vssd1 vccd1 vccd1 _03587_ sky130_fd_sc_hd__and3_1
X_13085_ img_gen.tracker.frame\[307\] net662 vssd1 vssd1 vccd1 vccd1 _07736_ sky130_fd_sc_hd__and2_1
X_10297_ _05260_ _05265_ _05267_ _05269_ vssd1 vssd1 vccd1 vccd1 _05270_ sky130_fd_sc_hd__or4_2
X_19701_ clknet_leaf_136_clk _00645_ net1300 vssd1 vssd1 vccd1 vccd1 control.body\[691\]
+ sky130_fd_sc_hd__dfrtp_1
X_12036_ img_gen.tracker.frame\[0\] net630 net612 img_gen.tracker.frame\[3\] vssd1
+ vssd1 vccd1 vccd1 _07008_ sky130_fd_sc_hd__a22o_1
X_16913_ ag2.body\[563\] net716 net698 ag2.body\[566\] vssd1 vssd1 vccd1 vccd1 _02592_
+ sky130_fd_sc_hd__a22o_1
X_17893_ _03532_ _03531_ obsg2.obstacleCount\[0\] vssd1 vssd1 vccd1 vccd1 _01247_
+ sky130_fd_sc_hd__mux2_1
XANTENNA__16076__C1 net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17812__B1 net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19632_ clknet_leaf_123_clk net2258 net1409 vssd1 vssd1 vccd1 vccd1 control.body\[766\]
+ sky130_fd_sc_hd__dfrtp_1
X_16844_ ag2.body\[170\] net862 vssd1 vssd1 vccd1 vccd1 _02523_ sky130_fd_sc_hd__or2_1
XANTENNA__14211__A net1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13429__A1 net225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16091__A2 net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19563_ clknet_leaf_116_clk _00507_ net1387 vssd1 vssd1 vccd1 vccd1 control.body\[825\]
+ sky130_fd_sc_hd__dfrtp_1
X_16775_ obsg2.obstacleArray\[31\] net503 net484 obsg2.obstacleArray\[29\] vssd1 vssd1
+ vccd1 vccd1 _02454_ sky130_fd_sc_hd__a22o_1
X_13987_ ag2.body\[124\] net211 _08159_ ag2.body\[116\] vssd1 vssd1 vccd1 vccd1 _00205_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__18368__A1 _07181_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18514_ net1512 net1506 vssd1 vssd1 vccd1 vccd1 _00045_ sky130_fd_sc_hd__or2_1
XANTENNA__09799__X _04772_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15726_ ag2.body\[355\] net200 _01632_ ag2.body\[347\] vssd1 vssd1 vccd1 vccd1 _00981_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_125_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19494_ clknet_leaf_113_clk _00438_ net1399 vssd1 vssd1 vccd1 vccd1 control.body\[900\]
+ sky130_fd_sc_hd__dfrtp_1
X_12938_ net269 _07665_ _07666_ net1819 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[229\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__16918__A2 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18445_ _04642_ _08026_ _03832_ _04645_ vssd1 vssd1 vccd1 vccd1 _03934_ sky130_fd_sc_hd__a211o_1
XANTENNA__17241__B net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15657_ ag2.body\[422\] net143 _01624_ ag2.body\[414\] vssd1 vssd1 vccd1 vccd1 _00920_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__09959__B net1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11860__B1 net607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12869_ net287 _07634_ _07635_ net2115 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[191\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_133_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11570__A net506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14608_ net821 ag2.body\[131\] ag2.body\[134\] net803 vssd1 vssd1 vccd1 vccd1 _08769_
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_51_1361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18376_ _04636_ _03849_ vssd1 vssd1 vccd1 vccd1 _03867_ sky130_fd_sc_hd__xnor2_1
X_15588_ _06351_ net56 vssd1 vssd1 vccd1 vccd1 _01618_ sky130_fd_sc_hd__nor2_2
XANTENNA__11838__S1 net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17327_ ag2.body\[2\] net860 vssd1 vssd1 vccd1 vccd1 _03006_ sky130_fd_sc_hd__xor2_2
XANTENNA__16572__S net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14539_ net1001 ag2.body\[240\] vssd1 vssd1 vccd1 vccd1 _08700_ sky130_fd_sc_hd__nand2_1
XFILLER_0_16_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_133_4373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_133_4384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_42_1590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17258_ _02930_ _02931_ _02932_ _02934_ vssd1 vssd1 vccd1 vccd1 _02937_ sky130_fd_sc_hd__or4_1
XANTENNA__16551__B1 net390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18551__CLK clknet_leaf_132_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16209_ net882 net860 net850 net870 vssd1 vssd1 vccd1 vccd1 _01888_ sky130_fd_sc_hd__and4bb_2
XFILLER_0_124_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09694__B net1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10179__B1 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17189_ ag2.body\[572\] net710 net705 ag2.body\[573\] _02867_ vssd1 vssd1 vccd1 vccd1
+ _02868_ sky130_fd_sc_hd__o221ai_1
XANTENNA__17726__S0 net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1012 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10718__A2 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_1177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09584__A2 _04556_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08962_ ag2.body\[41\] vssd1 vssd1 vccd1 vccd1 _03987_ sky130_fd_sc_hd__inv_2
XFILLER_0_23_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14865__B1 _01535_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_1995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_4188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_4199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout196_A net218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_1504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09887__A3 net923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17803__B1 net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_1564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_1515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14121__A net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14093__A1 net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14093__B2 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09514_ net1149 control.body\[835\] vssd1 vssd1 vccd1 vccd1 _04487_ sky130_fd_sc_hd__nand2_1
XFILLER_0_116_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09445_ net903 _04417_ vssd1 vssd1 vccd1 vccd1 _04418_ sky130_fd_sc_hd__nor2_4
XANTENNA__17151__B net958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09869__B net1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout530_A net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12576__A net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16048__A net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout628_A _06473_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1272_A net1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17582__A2 net741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout249_X net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09376_ sound_gen.osc1.stayCount\[16\] _04358_ vssd1 vssd1 vccd1 vccd1 _04373_ sky130_fd_sc_hd__nor2_1
XFILLER_0_93_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_1423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20605_ net1537 vssd1 vssd1 vccd1 vccd1 gpio_oeb[17] sky130_fd_sc_hd__buf_2
XFILLER_0_90_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11603__B1 net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16482__S net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10096__A net1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1060_X net1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14791__A net980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout416_X net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18263__A net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1158_X net1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20536_ clknet_leaf_107_clk _01401_ _00010_ vssd1 vssd1 vccd1 vccd1 sound_gen.osc1.stayCount\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_116_3870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout997_A net1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12159__B2 net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15896__A2 net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_3734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_112_3745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20467_ clknet_leaf_25_clk _01354_ net1340 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[103\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_63_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_1341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09643__A1_N net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10220_ ag2.body\[562\] net1172 vssd1 vssd1 vccd1 vccd1 _05193_ sky130_fd_sc_hd__or2_1
XFILLER_0_123_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20398_ clknet_leaf_27_clk _01285_ net1340 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[34\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA_fanout785_X net785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10543__B net1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15648__A2 net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10151_ ag2.body\[57\] net1208 vssd1 vssd1 vccd1 vccd1 _05124_ sky130_fd_sc_hd__xor2_1
XANTENNA__14856__B1 _08819_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17326__B net882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10082_ net1050 control.body\[799\] vssd1 vssd1 vccd1 vccd1 _05055_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout952_X net952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11655__A net1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13910_ _05120_ net57 vssd1 vssd1 vccd1 vccd1 _08151_ sky130_fd_sc_hd__nor2_2
XANTENNA__14031__A net977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14890_ control.body\[1100\] net179 _01539_ net2275 vssd1 vssd1 vccd1 vccd1 _00238_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__10342__B1 net745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout64_X net64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_3549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13841_ net686 net223 vssd1 vssd1 vccd1 vccd1 _08131_ sky130_fd_sc_hd__nor2_4
X_16560_ _02237_ _02238_ net395 vssd1 vssd1 vccd1 vccd1 _02239_ sky130_fd_sc_hd__mux2_1
XANTENNA__12095__B1 net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13772_ img_gen.updater.commands.count\[8\] _08082_ _08084_ _08071_ vssd1 vssd1 vccd1
+ vccd1 _00065_ sky130_fd_sc_hd__o211a_1
X_10984_ net1220 control.body\[752\] vssd1 vssd1 vccd1 vccd1 _05957_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_84_2870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_84_2881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_84_2892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15511_ ag2.body\[548\] net155 _01608_ ag2.body\[540\] vssd1 vssd1 vccd1 vccd1 _00790_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_85_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11842__B1 net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12723_ net247 _07565_ _07566_ net1710 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[114\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_112_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16491_ _01817_ _02105_ vssd1 vssd1 vccd1 vccd1 _02170_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_65_2291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17573__A2 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_2756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18230_ net353 _03539_ net37 obsg2.obstacleArray\[112\] vssd1 vssd1 vccd1 vccd1 _03754_
+ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_80_2767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_2778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12654_ net589 net435 net467 net574 vssd1 vssd1 vccd1 vccd1 _07531_ sky130_fd_sc_hd__or4_1
X_15442_ ag2.body\[615\] net90 _01600_ ag2.body\[607\] vssd1 vssd1 vccd1 vccd1 _00729_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_72_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09498__C net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_2177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11605_ net1126 _06574_ _06577_ _06485_ vssd1 vssd1 vccd1 vccd1 _06578_ sky130_fd_sc_hd__o211a_1
XFILLER_0_87_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12398__B2 net1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_2188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18161_ obsg2.obstacleArray\[77\] _03719_ net522 vssd1 vssd1 vccd1 vccd1 _01328_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_37_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12585_ net276 _07491_ _07492_ net1742 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[50\]
+ sky130_fd_sc_hd__a22o_1
X_15373_ net2211 net76 _01594_ net2423 vssd1 vssd1 vccd1 vccd1 _00666_ sky130_fd_sc_hd__a22o_1
XFILLER_0_68_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18173__A net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10948__A2 _04758_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1332 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17112_ ag2.body\[539\] net853 vssd1 vssd1 vccd1 vccd1 _02791_ sky130_fd_sc_hd__xnor2_1
X_14324_ _08480_ _08482_ _08483_ _08484_ vssd1 vssd1 vccd1 vccd1 _08485_ sky130_fd_sc_hd__or4_2
XFILLER_0_108_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11536_ _06479_ _06482_ _06494_ _06508_ vssd1 vssd1 vccd1 vccd1 _06509_ sky130_fd_sc_hd__a211o_1
XANTENNA__09795__A net1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18092_ net345 _03545_ _03557_ vssd1 vssd1 vccd1 vccd1 _03677_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_22_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_1176 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17043_ _02717_ _02718_ _02721_ vssd1 vssd1 vccd1 vccd1 _02722_ sky130_fd_sc_hd__or3b_4
X_14255_ net994 ag2.body\[73\] vssd1 vssd1 vccd1 vccd1 _08416_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_78_2696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11467_ _06435_ _06436_ _06437_ _06439_ vssd1 vssd1 vccd1 vccd1 _06440_ sky130_fd_sc_hd__or4_2
XFILLER_0_106_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13206_ _07793_ net263 _07791_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[370\]
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10418_ net786 control.body\[1064\] control.body\[1065\] net779 _05390_ vssd1 vssd1
+ vccd1 vccd1 _05391_ sky130_fd_sc_hd__o221a_1
XANTENNA__09566__A2 _04446_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14186_ net1017 ag2.body\[166\] vssd1 vssd1 vccd1 vccd1 _08347_ sky130_fd_sc_hd__or2_1
XFILLER_0_21_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11398_ _04236_ _04425_ _05133_ vssd1 vssd1 vccd1 vccd1 _06371_ sky130_fd_sc_hd__o21a_1
XANTENNA__10453__B net1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_1376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12570__A1 net245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13137_ net265 _07758_ vssd1 vssd1 vccd1 vccd1 _07761_ sky130_fd_sc_hd__nand2_1
X_10349_ ag2.body\[291\] net772 net788 ag2.body\[288\] vssd1 vssd1 vccd1 vccd1 _05322_
+ sky130_fd_sc_hd__a2bb2o_1
X_18994_ clknet_leaf_0_clk img_gen.tracker.next_frame\[432\] net1248 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[432\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17945_ _03540_ _03573_ vssd1 vssd1 vccd1 vccd1 _03574_ sky130_fd_sc_hd__and2_2
X_13068_ img_gen.tracker.frame\[298\] net661 vssd1 vssd1 vccd1 vccd1 _07728_ sky130_fd_sc_hd__and2_1
XFILLER_0_20_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1450 net1451 vssd1 vssd1 vccd1 vccd1 net1450 sky130_fd_sc_hd__clkbuf_4
X_12019_ img_gen.tracker.frame\[219\] net611 net556 img_gen.tracker.frame\[222\] _06990_
+ vssd1 vssd1 vccd1 vccd1 _06991_ sky130_fd_sc_hd__a221o_1
XFILLER_0_136_12 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1461 net1465 vssd1 vssd1 vccd1 vccd1 net1461 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_122_4030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1472 net1473 vssd1 vssd1 vccd1 vccd1 net1472 sky130_fd_sc_hd__clkbuf_2
X_17876_ _03507_ _03517_ vssd1 vssd1 vccd1 vccd1 _01245_ sky130_fd_sc_hd__and2_1
XANTENNA__12013__X _06985_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_122_4041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1483 net1484 vssd1 vssd1 vccd1 vccd1 net1483 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_122_4052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1494 net1495 vssd1 vssd1 vccd1 vccd1 net1494 sky130_fd_sc_hd__clkbuf_4
X_19615_ clknet_leaf_120_clk _00559_ net1394 vssd1 vssd1 vccd1 vccd1 control.body\[781\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10884__A1 _04556_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16827_ ag2.body\[224\] net885 vssd1 vssd1 vccd1 vccd1 _02506_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_31_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_1435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19546_ clknet_leaf_115_clk _00490_ net1397 vssd1 vssd1 vccd1 vccd1 control.body\[840\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_117_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16758_ obsg2.obstacleArray\[19\] net503 net489 obsg2.obstacleArray\[18\] vssd1 vssd1
+ vccd1 vccd1 _02437_ sky130_fd_sc_hd__a22o_1
XFILLER_0_88_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16139__Y _01818_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_0_clk_X clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15709_ ag2.body\[373\] net140 _01629_ ag2.body\[365\] vssd1 vssd1 vccd1 vccd1 _00967_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__09689__B net1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19477_ clknet_leaf_110_clk _00421_ net1418 vssd1 vssd1 vccd1 vccd1 control.body\[915\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11833__B1 net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16689_ _02227_ _02282_ _02286_ _02211_ vssd1 vssd1 vccd1 vccd1 _02368_ sky130_fd_sc_hd__a31o_1
XFILLER_0_75_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18917__CLK clknet_leaf_142_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15024__B1 _01555_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09230_ control.body\[1093\] vssd1 vssd1 vccd1 vccd1 _04255_ sky130_fd_sc_hd__inv_2
X_18428_ net321 _03793_ net325 vssd1 vssd1 vccd1 vccd1 _03917_ sky130_fd_sc_hd__o21a_1
XFILLER_0_57_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_135_4435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_4446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16772__B1 net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09161_ ag2.body\[510\] vssd1 vssd1 vccd1 vccd1 _04186_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_44_1663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12546__D net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18359_ _03791_ _03853_ _03851_ vssd1 vssd1 vccd1 vccd1 _03854_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_44_1674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13050__A2 _07718_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11597__C1 net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09092_ ag2.body\[335\] vssd1 vssd1 vccd1 vccd1 _04117_ sky130_fd_sc_hd__inv_2
XFILLER_0_114_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_1265 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20321_ clknet_leaf_43_clk _01217_ net1378 vssd1 vssd1 vccd1 vccd1 obsg2.randCord\[6\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_128_1553 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold900 _00510_ vssd1 vssd1 vccd1 vccd1 net2462 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10644__A _04573_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold911 control.body\[920\] vssd1 vssd1 vccd1 vccd1 net2473 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout209_A net210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold922 control.body\[826\] vssd1 vssd1 vccd1 vccd1 net2484 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13020__A net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20252_ clknet_leaf_70_clk _01196_ net1498 vssd1 vssd1 vccd1 vccd1 ag2.body\[138\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_128_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11459__B net1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold933 control.body\[840\] vssd1 vssd1 vccd1 vccd1 net2495 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_3063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold944 control.body\[952\] vssd1 vssd1 vccd1 vccd1 net2506 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_3074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold955 control.body\[805\] vssd1 vssd1 vccd1 vccd1 net2517 sky130_fd_sc_hd__dlygate4sd3_1
Xhold966 ag2.body\[588\] vssd1 vssd1 vccd1 vccd1 net2528 sky130_fd_sc_hd__dlygate4sd3_1
Xhold977 control.body\[1003\] vssd1 vssd1 vccd1 vccd1 net2539 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_38_1467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1020_A net1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09994_ _04573_ _04964_ _04965_ _04966_ vssd1 vssd1 vccd1 vccd1 _04967_ sky130_fd_sc_hd__or4b_2
Xhold988 _00570_ vssd1 vssd1 vccd1 vccd1 net2550 sky130_fd_sc_hd__dlygate4sd3_1
X_20183_ clknet_leaf_87_clk _01127_ net1460 vssd1 vssd1 vccd1 vccd1 ag2.body\[213\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__14838__B1 _08531_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold999 control.body\[935\] vssd1 vssd1 vccd1 vccd1 net2561 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1118_A net1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_1489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10349__A1_N ag2.body\[291\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08945_ net927 vssd1 vssd1 vccd1 vccd1 _03970_ sky130_fd_sc_hd__inv_2
XANTENNA__17146__B net946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13510__B1 net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout578_A net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16477__S net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout366_X net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout745_A net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_3402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_3413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12077__B1 net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_564 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16049__Y _01728_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12172__S0 net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18597__CLK clknet_leaf_13_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11824__B1 net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout533_X net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17555__A2 net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15015__B1 _01553_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16209__C net850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09428_ obsg2.obsNeeded\[0\] _04399_ _04400_ net2415 vssd1 vssd1 vccd1 vccd1 _00002_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_118_3910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16763__B1 net488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_118_3921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_3932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10538__B net1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout700_X net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09359_ sound_gen.osc1.stayCount\[18\] sound_gen.osc1.stayCount\[17\] _04360_ vssd1
+ vssd1 vccd1 vccd1 _04361_ sky130_fd_sc_hd__and3_1
XANTENNA__09886__Y _04859_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1442_X net1442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_114_3807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_883 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12370_ net293 vssd1 vssd1 vccd1 vccd1 _07336_ sky130_fd_sc_hd__inv_2
XANTENNA__17712__C1 net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10825__Y _05798_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11321_ _04203_ net1203 net1150 _04204_ _06293_ vssd1 vssd1 vccd1 vccd1 _06294_ sky130_fd_sc_hd__a221o_1
X_20519_ clknet_leaf_112_clk track.nextCurrScore\[1\] net1424 vssd1 vssd1 vccd1 vccd1
+ control.body_update.curr_length\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_127_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_1630 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14040_ net1023 ag2.body\[502\] vssd1 vssd1 vccd1 vccd1 _08201_ sky130_fd_sc_hd__xor2_1
XFILLER_0_15_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11252_ _06217_ _06218_ _06221_ _06222_ _06215_ vssd1 vssd1 vccd1 vccd1 _06225_ sky130_fd_sc_hd__a221o_1
XFILLER_0_43_1614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10273__B net1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_1096 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10203_ _05171_ _05172_ _05175_ _05163_ vssd1 vssd1 vccd1 vccd1 _05176_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_73_2560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11986__S0 net471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12552__A1 net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11183_ ag2.body\[179\] net1154 vssd1 vssd1 vccd1 vccd1 _06156_ sky130_fd_sc_hd__and2b_1
XFILLER_0_63_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10134_ net1075 control.body\[822\] vssd1 vssd1 vccd1 vccd1 _05107_ sky130_fd_sc_hd__or2_1
X_15991_ ag2.body\[3\] _08119_ vssd1 vssd1 vccd1 vccd1 _01674_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_98_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17730_ net496 _03408_ net461 vssd1 vssd1 vccd1 vccd1 _03409_ sky130_fd_sc_hd__a21oi_1
X_10065_ net1217 control.body\[712\] vssd1 vssd1 vccd1 vccd1 _05038_ sky130_fd_sc_hd__xor2_1
X_14942_ net2649 net168 _01545_ net2327 vssd1 vssd1 vccd1 vccd1 _00284_ sky130_fd_sc_hd__a22o_1
XANTENNA__19372__CLK clknet_leaf_102_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16895__B net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17661_ ag2.body\[108\] net711 net707 ag2.body\[109\] _03334_ vssd1 vssd1 vccd1 vccd1
+ _03340_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_86_2943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_86_2954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14873_ net2152 net181 _01537_ control.body\[1109\] vssd1 vssd1 vccd1 vccd1 _00223_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__14696__A net1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15254__B1 net50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19400_ clknet_leaf_102_clk _00344_ net1428 vssd1 vssd1 vccd1 vccd1 control.body\[998\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11672__X _06644_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16612_ obsg2.obstacleArray\[90\] net445 vssd1 vssd1 vccd1 vccd1 _02291_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_67_2353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13824_ _08111_ _08112_ _08117_ _08120_ _08116_ vssd1 vssd1 vccd1 vccd1 _08121_ sky130_fd_sc_hd__a41o_1
XTAP_TAPCELL_ROW_82_2818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_2364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_2829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17592_ ag2.body\[57\] net731 net689 ag2.body\[63\] _03270_ vssd1 vssd1 vccd1 vccd1
+ _03271_ sky130_fd_sc_hd__a221o_1
XANTENNA__13804__A1 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_2375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13804__B2 net1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19331_ clknet_leaf_100_clk _00275_ net1443 vssd1 vssd1 vccd1 vccd1 control.body\[1057\]
+ sky130_fd_sc_hd__dfrtp_1
X_16543_ _02220_ _02221_ vssd1 vssd1 vccd1 vccd1 _02222_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_63_2239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13755_ img_gen.updater.commands.count\[3\] _08068_ vssd1 vssd1 vccd1 vccd1 _08073_
+ sky130_fd_sc_hd__nand2_1
X_10967_ net1131 control.body\[1004\] vssd1 vssd1 vccd1 vccd1 _05940_ sky130_fd_sc_hd__and2_1
XANTENNA__15006__B1 _01552_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13280__A2 _07825_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13105__A net344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19262_ clknet_leaf_74_clk _00206_ net1495 vssd1 vssd1 vccd1 vccd1 ag2.body\[125\]
+ sky130_fd_sc_hd__dfrtp_4
X_12706_ net225 _07556_ vssd1 vssd1 vccd1 vccd1 _07557_ sky130_fd_sc_hd__nor2_1
X_16474_ obsg2.obstacleArray\[42\] net453 vssd1 vssd1 vccd1 vccd1 _02153_ sky130_fd_sc_hd__or2_1
XFILLER_0_85_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16754__B1 net486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13686_ net639 _04550_ vssd1 vssd1 vccd1 vccd1 _08029_ sky130_fd_sc_hd__nand2_1
X_10898_ net921 _04603_ _05074_ _05870_ vssd1 vssd1 vccd1 vccd1 _05871_ sky130_fd_sc_hd__o31a_1
XANTENNA__10448__B net1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18213_ obsg2.obstacleArray\[103\] _03745_ net521 vssd1 vssd1 vccd1 vccd1 _01354_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_72_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15425_ _05686_ net52 vssd1 vssd1 vccd1 vccd1 _01599_ sky130_fd_sc_hd__nor2_2
X_19193_ clknet_leaf_53_clk _00137_ net1455 vssd1 vssd1 vccd1 vccd1 ag2.body\[56\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_14_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12637_ net264 _07520_ _07521_ net1676 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[73\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__19855__RESET_B net1415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18144_ net47 _03566_ _03704_ obsg2.obstacleArray\[69\] vssd1 vssd1 vccd1 vccd1 _03711_
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_124_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15356_ control.body\[681\] net68 _01592_ net2453 vssd1 vssd1 vccd1 vccd1 _00651_
+ sky130_fd_sc_hd__a22o_1
X_12568_ net315 _07483_ net343 net335 vssd1 vssd1 vccd1 vccd1 _07484_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_41_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12663__B _07536_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16135__B net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11594__A2 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14307_ net1026 ag2.body\[53\] vssd1 vssd1 vccd1 vccd1 _08468_ sky130_fd_sc_hd__xor2_1
XFILLER_0_53_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11519_ net1222 net1152 vssd1 vssd1 vccd1 vccd1 _06492_ sky130_fd_sc_hd__and2b_1
X_18075_ net301 _03594_ vssd1 vssd1 vccd1 vccd1 _03666_ sky130_fd_sc_hd__nand2_1
X_15287_ control.body\[748\] net87 _01584_ net2450 vssd1 vssd1 vccd1 vccd1 _00590_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__10464__A net1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12499_ net384 net344 vssd1 vssd1 vccd1 vccd1 _07445_ sky130_fd_sc_hd__nand2_1
Xhold207 img_gen.tracker.frame\[43\] vssd1 vssd1 vccd1 vccd1 net1769 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold218 img_gen.tracker.frame\[303\] vssd1 vssd1 vccd1 vccd1 net1780 sky130_fd_sc_hd__dlygate4sd3_1
X_17026_ ag2.body\[404\] net963 vssd1 vssd1 vccd1 vccd1 _02705_ sky130_fd_sc_hd__xor2_1
XFILLER_0_40_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold229 img_gen.tracker.frame\[384\] vssd1 vssd1 vccd1 vccd1 net1791 sky130_fd_sc_hd__dlygate4sd3_1
X_14238_ net819 ag2.body\[483\] ag2.body\[487\] net791 _08398_ vssd1 vssd1 vccd1 vccd1
+ _08399_ sky130_fd_sc_hd__a221o_1
XFILLER_0_1_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10183__B net1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16809__A1 ag2.body\[67\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14169_ net807 ag2.body\[205\] ag2.body\[207\] net791 _08329_ vssd1 vssd1 vccd1 vccd1
+ _08330_ sky130_fd_sc_hd__a221o_1
XFILLER_0_22_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout709 net710 vssd1 vssd1 vccd1 vccd1 net709 sky130_fd_sc_hd__buf_4
XFILLER_0_0_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_52_1910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19715__CLK clknet_leaf_132_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_4103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_4114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20342__RESET_B net1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18977_ clknet_leaf_7_clk img_gen.tracker.next_frame\[415\] net1265 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[415\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_33_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11295__A net1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17928_ net516 _03560_ vssd1 vssd1 vccd1 vccd1 _01254_ sky130_fd_sc_hd__nor2_1
XFILLER_0_56_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_1523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1280 net1287 vssd1 vssd1 vccd1 vccd1 net1280 sky130_fd_sc_hd__buf_2
Xfanout1291 net1293 vssd1 vssd1 vccd1 vccd1 net1291 sky130_fd_sc_hd__clkbuf_2
XANTENNA__14048__A1 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17859_ net2193 _03511_ _03499_ vssd1 vssd1 vccd1 vccd1 _01234_ sky130_fd_sc_hd__o21a_1
XANTENNA__16297__S net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1556 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18078__A net300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14048__B2 net811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12059__B1 net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16993__B1 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_137_4508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_1276 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19529_ clknet_leaf_120_clk _00473_ net1395 vssd1 vssd1 vccd1 vccd1 control.body\[871\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11742__B net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10639__A net1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_1736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout159_A net161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13015__A net668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_27_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10358__B ag2.body\[290\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09213_ net904 vssd1 vssd1 vccd1 vccd1 _04238_ sky130_fd_sc_hd__inv_4
XFILLER_0_107_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1349 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12854__A net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_96_3250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_96_3261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09144_ ag2.body\[475\] vssd1 vssd1 vccd1 vccd1 _04169_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout1068_A net1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11034__A1 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11034__B2 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09778__A2 net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_3114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12573__B _06639_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_3125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19525__RESET_B net1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_3136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19245__CLK clknet_leaf_83_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12782__A1 net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09075_ ag2.body\[302\] vssd1 vssd1 vccd1 vccd1 _04100_ sky130_fd_sc_hd__inv_2
XFILLER_0_60_957 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout114_X net114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1235_A net1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20304_ clknet_leaf_37_clk net1567 net1351 vssd1 vssd1 vccd1 vccd1 control.divider.detect.Q\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_124_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold730 control.body\[671\] vssd1 vssd1 vccd1 vccd1 net2292 sky130_fd_sc_hd__dlygate4sd3_1
Xhold741 control.body\[1045\] vssd1 vssd1 vccd1 vccd1 net2303 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold752 control.body\[736\] vssd1 vssd1 vccd1 vccd1 net2314 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20235_ clknet_leaf_69_clk _01179_ net1499 vssd1 vssd1 vccd1 vccd1 ag2.body\[153\]
+ sky130_fd_sc_hd__dfrtp_4
Xhold763 control.body\[1094\] vssd1 vssd1 vccd1 vccd1 net2325 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_99_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_383 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold774 control.body\[666\] vssd1 vssd1 vccd1 vccd1 net2336 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10661__X _05634_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1023_X net1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold785 control.body\[690\] vssd1 vssd1 vccd1 vccd1 net2347 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1402_A net1403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold796 control.body\[919\] vssd1 vssd1 vccd1 vccd1 net2358 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__19395__CLK clknet_leaf_103_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20166_ clknet_leaf_81_clk _01110_ net1484 vssd1 vssd1 vccd1 vccd1 ag2.body\[228\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA_fanout862_A net867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout483_X net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09977_ net787 control.body\[1112\] control.body\[1115\] net770 _04949_ vssd1 vssd1
+ vccd1 vccd1 _04950_ sky130_fd_sc_hd__o221ai_1
XTAP_TAPCELL_ROW_107_3600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15484__B1 _01605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16681__C1 _02211_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20097_ clknet_leaf_78_clk _01041_ net1490 vssd1 vssd1 vccd1 vccd1 ag2.body\[303\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_99_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout748_X net748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11870_ img_gen.tracker.frame\[277\] net615 net604 img_gen.tracker.frame\[280\] vssd1
+ vssd1 vccd1 vccd1 _06842_ sky130_fd_sc_hd__o22a_1
XANTENNA__16984__B1 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10821_ net1231 control.body\[1088\] vssd1 vssd1 vccd1 vccd1 _05794_ sky130_fd_sc_hd__and2b_1
XANTENNA__11652__B net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout915_X net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13540_ net2108 net655 _07927_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[570\]
+ sky130_fd_sc_hd__and3_1
X_10752_ _05644_ _05669_ _05696_ _05724_ vssd1 vssd1 vccd1 vccd1 _05725_ sky130_fd_sc_hd__nand4_1
XANTENNA__16736__B1 net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10268__B net1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13471_ net666 _07900_ vssd1 vssd1 vccd1 vccd1 _07901_ sky130_fd_sc_hd__nor2_1
X_10683_ _05647_ _05651_ _05654_ _05655_ vssd1 vssd1 vccd1 vccd1 _05656_ sky130_fd_sc_hd__or4_1
XFILLER_0_10_1613 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15210_ control.body\[808\] net95 _01575_ control.body\[800\] vssd1 vssd1 vccd1 vccd1
+ _00522_ sky130_fd_sc_hd__a22o_1
X_12422_ net1094 _06626_ _06643_ vssd1 vssd1 vccd1 vccd1 _07384_ sky130_fd_sc_hd__o21a_1
XFILLER_0_118_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16190_ _01865_ _01868_ net346 vssd1 vssd1 vccd1 vccd1 _01869_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19266__RESET_B net1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_1271 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_2600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_2611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12353_ _07254_ _07285_ vssd1 vssd1 vccd1 vccd1 _07320_ sky130_fd_sc_hd__nor2_1
X_15141_ net2620 net106 _01567_ net2367 vssd1 vssd1 vccd1 vccd1 _00461_ sky130_fd_sc_hd__a22o_1
XFILLER_0_121_801 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_2622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_2021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11304_ _06269_ _06271_ _06274_ _06275_ vssd1 vssd1 vccd1 vccd1 _06277_ sky130_fd_sc_hd__or4_2
X_15072_ net2300 net150 _01560_ net2353 vssd1 vssd1 vccd1 vccd1 _00399_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_56_2032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11099__B net1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12284_ _07248_ _07252_ _04273_ _07241_ vssd1 vssd1 vccd1 vccd1 _07254_ sky130_fd_sc_hd__a2bb2o_2
XTAP_TAPCELL_ROW_56_2043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18170__B _03706_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12525__A1 net227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14023_ net970 ag2.body\[27\] vssd1 vssd1 vccd1 vccd1 _08184_ sky130_fd_sc_hd__xor2_1
XFILLER_0_82_1471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18900_ clknet_leaf_144_clk img_gen.tracker.next_frame\[338\] net1252 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[338\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_120_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11235_ _06201_ _06206_ _06207_ _06193_ vssd1 vssd1 vccd1 vccd1 _06208_ sky130_fd_sc_hd__o31a_1
X_19880_ clknet_leaf_82_clk _00824_ net1479 vssd1 vssd1 vccd1 vccd1 ag2.body\[518\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__09917__A2_N net772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18831_ clknet_leaf_142_clk img_gen.tracker.next_frame\[269\] net1261 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[269\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_101_580 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09941__A2 net1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11166_ net1131 control.body\[780\] vssd1 vssd1 vccd1 vccd1 _06139_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_8_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_8_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10731__B net1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18762__CLK clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10117_ net1121 control.body\[708\] vssd1 vssd1 vccd1 vccd1 _05090_ sky130_fd_sc_hd__nand2_1
X_18762_ clknet_leaf_16_clk img_gen.tracker.next_frame\[200\] net1313 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[200\] sky130_fd_sc_hd__dfrtp_1
X_11097_ ag2.body\[427\] net1154 vssd1 vssd1 vccd1 vccd1 _06070_ sky130_fd_sc_hd__xnor2_1
X_15974_ net223 _08118_ net663 vssd1 vssd1 vccd1 vccd1 _01660_ sky130_fd_sc_hd__o21a_1
XFILLER_0_120_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_2415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_69_2426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_2437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17713_ obsg2.obstacleArray\[136\] obsg2.obstacleArray\[137\] obsg2.obstacleArray\[138\]
+ obsg2.obstacleArray\[139\] net446 net392 vssd1 vssd1 vccd1 vccd1 _03392_ sky130_fd_sc_hd__mux4_1
X_10048_ _04551_ _05015_ _05020_ vssd1 vssd1 vccd1 vccd1 _05021_ sky130_fd_sc_hd__or3_2
X_14925_ control.body\[1067\] net177 _01543_ net2319 vssd1 vssd1 vccd1 vccd1 _00269_
+ sky130_fd_sc_hd__a22o_1
X_18693_ clknet_leaf_28_clk img_gen.tracker.next_frame\[131\] net1336 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[131\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__10839__B2 _05811_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold90 img_gen.tracker.frame\[550\] vssd1 vssd1 vccd1 vccd1 net1652 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_118_1530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17644_ _03316_ _03322_ vssd1 vssd1 vccd1 vccd1 _03323_ sky130_fd_sc_hd__or2_1
XFILLER_0_118_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19118__CLK clknet_leaf_131_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14856_ _08738_ _08743_ _08819_ vssd1 vssd1 vccd1 vccd1 _01527_ sky130_fd_sc_hd__o21a_1
XFILLER_0_89_169 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1128 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13807_ _06557_ _08104_ vssd1 vssd1 vccd1 vccd1 _08108_ sky130_fd_sc_hd__nand2_1
X_17575_ ag2.body\[338\] net866 vssd1 vssd1 vccd1 vccd1 _03254_ sky130_fd_sc_hd__xor2_1
XANTENNA__09457__A1 net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14787_ net837 ag2.body\[545\] _04201_ net974 vssd1 vssd1 vccd1 vccd1 _01458_ sky130_fd_sc_hd__o22a_1
XANTENNA__14450__A1 net846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11999_ img_gen.tracker.frame\[448\] net597 vssd1 vssd1 vccd1 vccd1 _06971_ sky130_fd_sc_hd__or2_1
X_19314_ clknet_leaf_104_clk _00258_ net1435 vssd1 vssd1 vccd1 vccd1 control.body\[1072\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14450__B2 net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16526_ _01709_ net497 _01737_ _02203_ vssd1 vssd1 vccd1 vccd1 _02205_ sky130_fd_sc_hd__a31o_1
XFILLER_0_133_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13738_ _07187_ _07248_ _08058_ _07240_ vssd1 vssd1 vccd1 vccd1 _08059_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_54_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19245_ clknet_leaf_83_clk _00189_ net1482 vssd1 vssd1 vccd1 vccd1 ag2.body\[108\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__09967__B net1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16457_ net365 _02110_ _02114_ _02075_ vssd1 vssd1 vccd1 vccd1 _02136_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_6_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13669_ net480 _06634_ _07171_ vssd1 vssd1 vccd1 vccd1 coll.nextGoodColl sky130_fd_sc_hd__and3_1
XFILLER_0_112_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15408_ control.body\[632\] net83 _01597_ net2491 vssd1 vssd1 vccd1 vccd1 _00698_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_109_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19176_ clknet_leaf_52_clk _00120_ net1366 vssd1 vssd1 vccd1 vccd1 ag2.body\[39\]
+ sky130_fd_sc_hd__dfrtp_2
X_16388_ _02065_ _02066_ vssd1 vssd1 vccd1 vccd1 _02067_ sky130_fd_sc_hd__nor2_1
XFILLER_0_115_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12764__A1 net237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18127_ net38 _03699_ vssd1 vssd1 vccd1 vccd1 _03700_ sky130_fd_sc_hd__and2_1
XFILLER_0_13_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15339_ control.body\[698\] net71 _01590_ net2347 vssd1 vssd1 vccd1 vccd1 _00636_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__16580__S net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_659 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_1523 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09983__A net1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18058_ net43 _03654_ vssd1 vssd1 vccd1 vccd1 _03655_ sky130_fd_sc_hd__nor2_1
XFILLER_0_13_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11319__A2 net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09900_ ag2.body\[73\] net781 net757 ag2.body\[77\] _04867_ vssd1 vssd1 vccd1 vccd1
+ _04873_ sky130_fd_sc_hd__a221o_1
X_17009_ ag2.body\[502\] net942 vssd1 vssd1 vccd1 vccd1 _02688_ sky130_fd_sc_hd__xor2_1
XFILLER_0_61_1522 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_1404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout506 net508 vssd1 vssd1 vccd1 vccd1 net506 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_6_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20020_ clknet_leaf_57_clk _00964_ net1464 vssd1 vssd1 vccd1 vccd1 ag2.body\[370\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_6_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_1566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout517 net518 vssd1 vssd1 vccd1 vccd1 net517 sky130_fd_sc_hd__buf_2
X_09831_ net1229 control.body\[920\] vssd1 vssd1 vccd1 vccd1 _04804_ sky130_fd_sc_hd__or2_1
Xfanout528 net534 vssd1 vssd1 vccd1 vccd1 net528 sky130_fd_sc_hd__buf_2
XANTENNA__15209__B net53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12531__A4 _07460_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout539 _01680_ vssd1 vssd1 vccd1 vccd1 net539 sky130_fd_sc_hd__clkbuf_4
XANTENNA_clkload13_A clknet_leaf_144_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15466__B1 _01603_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09762_ ag2.body\[208\] net1237 vssd1 vssd1 vccd1 vccd1 _04735_ sky130_fd_sc_hd__xor2_1
XFILLER_0_77_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09693_ ag2.body\[65\] net1208 vssd1 vssd1 vccd1 vccd1 _04666_ sky130_fd_sc_hd__nand2_1
XANTENNA__17758__A2 _02211_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16415__C1 net366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout276_A net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16966__B1 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11472__B net1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18095__X _03679_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout443_A _02214_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1185_A net1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_3301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_3312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_3323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17797__D net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09877__B net1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout231_X net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout610_A _06475_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1352_A net1356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout708_A _04267_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18635__CLK clknet_leaf_131_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15941__A1 ag2.body\[163\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11558__A2 net633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09127_ ag2.body\[429\] vssd1 vssd1 vccd1 vccd1 _04152_ sky130_fd_sc_hd__inv_2
XANTENNA__17143__B1 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1140_X net1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09620__A1 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1444 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18271__A net534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09620__B2 net777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1238_X net1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09058_ ag2.body\[253\] vssd1 vssd1 vccd1 vccd1 _04083_ sky130_fd_sc_hd__inv_2
XFILLER_0_103_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout698_X net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold560 sound_gen.dac1.dacCount\[3\] vssd1 vssd1 vccd1 vccd1 net2122 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10518__B1 net1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold571 img_gen.tracker.frame\[69\] vssd1 vssd1 vccd1 vccd1 net2133 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout91_A net219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11020_ ag2.body\[593\] net1196 vssd1 vssd1 vccd1 vccd1 _05993_ sky130_fd_sc_hd__or2_1
Xhold582 _00225_ vssd1 vssd1 vccd1 vccd1 net2144 sky130_fd_sc_hd__dlygate4sd3_1
X_20218_ clknet_leaf_61_clk _01162_ net1469 vssd1 vssd1 vccd1 vccd1 ag2.body\[168\]
+ sky130_fd_sc_hd__dfrtp_4
Xhold593 img_gen.tracker.frame\[21\] vssd1 vssd1 vccd1 vccd1 net2155 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__15119__B net58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11623__C_N _06497_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout865_X net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15457__B1 _01602_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10551__B net1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16654__C1 net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11730__A2 net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20149_ clknet_leaf_98_clk _01093_ net1449 vssd1 vssd1 vccd1 vccd1 ag2.body\[243\]
+ sky130_fd_sc_hd__dfrtp_2
X_12971_ net233 _07681_ _07682_ net1844 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[246\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_137_1438 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14680__A1 net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14680__B2 net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11663__A net1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14710_ _08863_ _08865_ _08869_ _08870_ vssd1 vssd1 vccd1 vccd1 _08871_ sky130_fd_sc_hd__or4_1
X_11922_ _06890_ _06892_ _06893_ net565 vssd1 vssd1 vccd1 vccd1 _06894_ sky130_fd_sc_hd__a22oi_1
X_15690_ ag2.body\[388\] net140 _01616_ ag2.body\[380\] vssd1 vssd1 vccd1 vccd1 _00950_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_99_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16957__B1 net692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14466__A1_N net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14641_ net1031 ag2.body\[517\] vssd1 vssd1 vccd1 vccd1 _08802_ sky130_fd_sc_hd__xor2_1
XFILLER_0_86_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11853_ net384 _06775_ _06801_ _06824_ vssd1 vssd1 vccd1 vccd1 _06825_ sky130_fd_sc_hd__a22o_1
XANTENNA__19410__CLK clknet_leaf_103_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14974__A net637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17360_ net1044 _03008_ vssd1 vssd1 vccd1 vccd1 _03039_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_0_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10804_ ag2.body\[37\] net1103 vssd1 vssd1 vccd1 vccd1 _05777_ sky130_fd_sc_hd__xor2_1
XANTENNA__16709__B1 net483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14572_ net812 ag2.body\[492\] ag2.body\[495\] net791 vssd1 vssd1 vccd1 vccd1 _08733_
+ sky130_fd_sc_hd__a22o_1
X_11784_ img_gen.tracker.frame\[173\] net603 net564 _06755_ vssd1 vssd1 vccd1 vccd1
+ _06756_ sky130_fd_sc_hd__o211a_1
XANTENNA__08972__A ag2.body\[61\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20268__CLK clknet_leaf_37_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16311_ net415 _01989_ _01988_ net369 vssd1 vssd1 vccd1 vccd1 _01990_ sky130_fd_sc_hd__a211o_1
XFILLER_0_113_1471 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13523_ net1980 net657 _07919_ _07920_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[560\]
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_103_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17291_ _02968_ _02969_ vssd1 vssd1 vccd1 vccd1 _02970_ sky130_fd_sc_hd__nand2b_1
X_10735_ ag2.body\[248\] net786 net1111 _04083_ vssd1 vssd1 vccd1 vccd1 _05708_ sky130_fd_sc_hd__o22a_1
XANTENNA__11602__S net514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19030_ clknet_leaf_6_clk img_gen.tracker.next_frame\[468\] net1265 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[468\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14196__B1 ag2.body\[167\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16242_ obsg2.obstacleArray\[42\] obsg2.obstacleArray\[43\] net404 vssd1 vssd1 vccd1
+ vccd1 _01921_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13454_ net281 _07892_ _07893_ net2112 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[518\]
+ sky130_fd_sc_hd__a22o_1
X_10666_ net762 control.body\[884\] _04246_ net1083 _05635_ vssd1 vssd1 vccd1 vccd1
+ _05639_ sky130_fd_sc_hd__a221o_1
XFILLER_0_125_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15932__B2 ag2.body\[162\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_2105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10726__B net1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12746__A1 net237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12405_ img_gen.updater.commands.rR1.rainbowRNG\[4\] net248 net241 vssd1 vssd1 vccd1
+ vccd1 _07368_ sky130_fd_sc_hd__a21o_1
X_16173_ _01850_ _01851_ net374 vssd1 vssd1 vccd1 vccd1 _01852_ sky130_fd_sc_hd__mux2_1
X_13385_ net255 _07866_ _07867_ net2055 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[475\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__18181__A net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10597_ _05560_ _05561_ _05563_ _05564_ _05568_ vssd1 vssd1 vccd1 vccd1 _05570_ sky130_fd_sc_hd__a221o_1
XFILLER_0_134_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11954__C1 net473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15124_ net2657 net103 _01565_ control.body\[884\] vssd1 vssd1 vccd1 vccd1 _00446_
+ sky130_fd_sc_hd__a22o_1
X_12336_ _07173_ _07302_ vssd1 vssd1 vccd1 vccd1 _07303_ sky130_fd_sc_hd__and2b_1
XANTENNA__17509__B net961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_1599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14499__A1 net838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11397__X _06370_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14499__B2 net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19932_ clknet_leaf_47_clk _00876_ net1375 vssd1 vssd1 vccd1 vccd1 ag2.body\[458\]
+ sky130_fd_sc_hd__dfrtp_4
X_12267_ img_gen.updater.commands.count\[16\] img_gen.updater.commands.count\[10\]
+ img_gen.updater.commands.count\[11\] _07236_ vssd1 vssd1 vccd1 vccd1 _07237_ sky130_fd_sc_hd__or4_1
X_15055_ control.body\[958\] net163 _01558_ net2427 vssd1 vssd1 vccd1 vccd1 _00384_
+ sky130_fd_sc_hd__a22o_1
X_14006_ net1021 ag2.body\[510\] vssd1 vssd1 vccd1 vccd1 _08167_ sky130_fd_sc_hd__nand2_1
X_11218_ net1130 control.body\[844\] vssd1 vssd1 vccd1 vccd1 _06191_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_43_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19863_ clknet_leaf_94_clk _00807_ net1436 vssd1 vssd1 vccd1 vccd1 ag2.body\[533\]
+ sky130_fd_sc_hd__dfrtp_4
X_12198_ _07169_ vssd1 vssd1 vccd1 vccd1 _07170_ sky130_fd_sc_hd__inv_2
XFILLER_0_120_1431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_1296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15448__B1 _01601_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11721__A2 net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11149_ _06040_ _06065_ _06091_ _06121_ vssd1 vssd1 vccd1 vccd1 _06122_ sky130_fd_sc_hd__or4b_2
X_18814_ clknet_leaf_2_clk img_gen.tracker.next_frame\[252\] net1249 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[252\] sky130_fd_sc_hd__dfrtp_1
X_19794_ clknet_leaf_127_clk _00738_ net1330 vssd1 vssd1 vccd1 vccd1 ag2.body\[592\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_37_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_113_clk_X clknet_leaf_113_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18745_ clknet_leaf_143_clk img_gen.tracker.next_frame\[183\] net1255 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[183\] sky130_fd_sc_hd__dfrtp_1
X_15957_ ag2.body\[145\] net198 _01657_ ag2.body\[137\] vssd1 vssd1 vccd1 vccd1 _01187_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12669__A net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14671__A1 net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14671__B2 net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14908_ control.body\[1084\] net178 _01541_ control.body\[1076\] vssd1 vssd1 vccd1
+ vccd1 _00254_ sky130_fd_sc_hd__a22o_1
X_18676_ clknet_leaf_27_clk img_gen.tracker.next_frame\[114\] net1339 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[114\] sky130_fd_sc_hd__dfrtp_1
X_15888_ ag2.body\[212\] net184 _01649_ ag2.body\[204\] vssd1 vssd1 vccd1 vccd1 _01126_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_118_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17627_ ag2.body\[186\] net725 net718 ag2.body\[187\] _03305_ vssd1 vssd1 vccd1 vccd1
+ _03306_ sky130_fd_sc_hd__a221o_1
X_14839_ _01463_ _01466_ _08391_ vssd1 vssd1 vccd1 vccd1 _01510_ sky130_fd_sc_hd__o21a_1
XANTENNA__10189__A net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18356__A net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09978__A net1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17558_ ag2.body\[355\] net855 vssd1 vssd1 vccd1 vccd1 _03237_ sky130_fd_sc_hd__xor2_1
XFILLER_0_92_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_824 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19188__RESET_B net1332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16509_ obsg2.obstacleArray\[12\] obsg2.obstacleArray\[13\] net456 vssd1 vssd1 vccd1
+ vccd1 _02188_ sky130_fd_sc_hd__mux2_1
XANTENNA__11788__A2 net615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09697__B net1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17489_ _04129_ net888 net693 ag2.body\[367\] _03167_ vssd1 vssd1 vccd1 vccd1 _03168_
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_131_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09850__A1 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_937 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09850__B2 net1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19228_ clknet_leaf_75_clk _00172_ net1483 vssd1 vssd1 vccd1 vccd1 ag2.body\[91\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_5_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19159_ clknet_leaf_52_clk _00103_ net1367 vssd1 vssd1 vccd1 vccd1 ag2.body\[23\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_6_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11748__A net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14124__A net1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_1461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13162__A1 net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout303 net304 vssd1 vssd1 vccd1 vccd1 net303 sky130_fd_sc_hd__clkbuf_2
Xfanout314 net315 vssd1 vssd1 vccd1 vccd1 net314 sky130_fd_sc_hd__buf_2
Xfanout325 track.nextHighScore\[3\] vssd1 vssd1 vccd1 vccd1 net325 sky130_fd_sc_hd__buf_2
X_20003_ clknet_leaf_59_clk _00947_ net1467 vssd1 vssd1 vccd1 vccd1 ag2.body\[385\]
+ sky130_fd_sc_hd__dfrtp_4
Xfanout336 net337 vssd1 vssd1 vccd1 vccd1 net336 sky130_fd_sc_hd__clkbuf_2
Xfanout347 _01732_ vssd1 vssd1 vccd1 vccd1 net347 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_103_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09814_ net1061 control.body\[1055\] vssd1 vssd1 vccd1 vccd1 _04787_ sky130_fd_sc_hd__xnor2_1
Xfanout369 _01908_ vssd1 vssd1 vccd1 vccd1 net369 sky130_fd_sc_hd__buf_4
XANTENNA_fanout1100_A net1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09745_ net642 _04421_ vssd1 vssd1 vccd1 vccd1 _04718_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout560_A net562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout279_X net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11483__A _06370_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09676_ ag2.body\[13\] net1102 vssd1 vssd1 vccd1 vccd1 _04649_ sky130_fd_sc_hd__nand2_1
XFILLER_0_49_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout825_A net827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1090_X net1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout446_X net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15611__B1 _01620_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1188_X net1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16057__Y _01736_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_610 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18156__A2 _03586_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_695 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11779__A2 net580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout613_X net613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1355_X net1355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10520_ _04421_ net634 _05486_ _05487_ vssd1 vssd1 vccd1 vccd1 _05493_ sky130_fd_sc_hd__o211a_1
XANTENNA__13203__A net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10546__B net1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10451_ _05420_ _05421_ _05422_ _05423_ vssd1 vssd1 vccd1 vccd1 _05424_ sky130_fd_sc_hd__a22o_1
XANTENNA__17116__B1 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13170_ net231 _07775_ _07776_ net1816 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[351\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_21_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10382_ ag2.body\[104\] net1237 vssd1 vssd1 vccd1 vccd1 _05355_ sky130_fd_sc_hd__xor2_1
XANTENNA_fanout982_X net982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17329__B net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15678__B1 _01627_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12121_ net386 _07065_ _07092_ _06723_ vssd1 vssd1 vccd1 vccd1 _07093_ sky130_fd_sc_hd__o31a_1
XFILLER_0_102_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11951__A2 net619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_1415 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14034__A net1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13153__A1 net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12052_ _07017_ _07019_ _07023_ _07021_ net570 net472 vssd1 vssd1 vccd1 vccd1 _07024_
+ sky130_fd_sc_hd__mux4_1
Xhold390 img_gen.tracker.frame\[311\] vssd1 vssd1 vccd1 vccd1 net1952 sky130_fd_sc_hd__dlygate4sd3_1
X_11003_ net786 control.body\[1080\] control.body\[1087\] net745 vssd1 vssd1 vccd1
+ vccd1 _05976_ sky130_fd_sc_hd__a22oi_1
X_16860_ ag2.body\[205\] net706 net700 ag2.body\[206\] vssd1 vssd1 vccd1 vccd1 _02539_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_40_1458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10911__B1 _05855_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout870 net871 vssd1 vssd1 vccd1 vccd1 net870 sky130_fd_sc_hd__buf_4
X_15811_ ag2.body\[287\] net207 _01641_ ag2.body\[279\] vssd1 vssd1 vccd1 vccd1 _01057_
+ sky130_fd_sc_hd__a22o_1
Xfanout881 net889 vssd1 vssd1 vccd1 vccd1 net881 sky130_fd_sc_hd__clkbuf_8
XANTENNA__17064__B net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16791_ obsg2.obstacleArray\[130\] obsg2.obstacleArray\[131\] net457 vssd1 vssd1
+ vccd1 vccd1 _02470_ sky130_fd_sc_hd__mux2_1
Xfanout892 net893 vssd1 vssd1 vccd1 vccd1 net892 sky130_fd_sc_hd__buf_4
XANTENNA__12489__A net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18530_ clknet_leaf_138_clk _00056_ net1292 vssd1 vssd1 vccd1 vccd1 img_gen.updater.commands.cmd_num\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11393__A net1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15742_ ag2.body\[337\] net215 _01634_ ag2.body\[329\] vssd1 vssd1 vccd1 vccd1 _00995_
+ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_82_clk_A clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1212 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12954_ net246 _07673_ _07674_ net1760 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[237\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_137_1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1090 control.body\[840\] vssd1 vssd1 vccd1 vccd1 net2652 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_1354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11044__D_N _05973_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19926__CLK clknet_leaf_51_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_1511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11905_ img_gen.tracker.frame\[367\] net549 net564 vssd1 vssd1 vccd1 vccd1 _06877_
+ sky130_fd_sc_hd__o21a_1
X_18461_ net2078 _08024_ _03932_ _03949_ vssd1 vssd1 vccd1 vccd1 _01398_ sky130_fd_sc_hd__o22a_1
X_15673_ ag2.body\[404\] net142 _01626_ ag2.body\[396\] vssd1 vssd1 vccd1 vccd1 _00934_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12639__D net574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12885_ net292 _07641_ _07642_ net1925 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[200\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_114_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15602__B1 _01619_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17412_ ag2.body\[287\] net692 net740 ag2.body\[280\] vssd1 vssd1 vccd1 vccd1 _03091_
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_16_1630 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14624_ net1027 ag2.body\[469\] vssd1 vssd1 vccd1 vccd1 _08785_ sky130_fd_sc_hd__xor2_1
X_18392_ _08051_ _03810_ _08137_ vssd1 vssd1 vccd1 vccd1 _03882_ sky130_fd_sc_hd__o21ai_1
X_11836_ img_gen.tracker.frame\[554\] net622 net604 img_gen.tracker.frame\[557\] vssd1
+ vssd1 vccd1 vccd1 _06808_ sky130_fd_sc_hd__o22a_1
XFILLER_0_90_1581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19281__RESET_B net1451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16408__B net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12967__A1 net254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_97_clk_A clknet_4_11__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17343_ net925 net948 vssd1 vssd1 vccd1 vccd1 _03022_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_23_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16158__A1 _01743_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14555_ net981 _04000_ ag2.body\[69\] net809 _08715_ vssd1 vssd1 vccd1 vccd1 _08716_
+ sky130_fd_sc_hd__o221a_1
X_11767_ img_gen.tracker.frame\[50\] net613 net596 img_gen.tracker.frame\[53\] vssd1
+ vssd1 vccd1 vccd1 _06739_ sky130_fd_sc_hd__o22a_1
XANTENNA__18950__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14209__A net1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_140_clk_A clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13506_ net664 _07914_ vssd1 vssd1 vccd1 vccd1 _07915_ sky130_fd_sc_hd__nor2_1
XFILLER_0_82_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17274_ ag2.body\[555\] net849 vssd1 vssd1 vccd1 vccd1 _02953_ sky130_fd_sc_hd__xor2_1
X_10718_ ag2.body\[617\] net777 net766 ag2.body\[620\] vssd1 vssd1 vccd1 vccd1 _05691_
+ sky130_fd_sc_hd__a22o_1
X_14486_ net1003 ag2.body\[344\] vssd1 vssd1 vccd1 vccd1 _08647_ sky130_fd_sc_hd__xor2_1
XFILLER_0_99_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11698_ _06631_ _06669_ vssd1 vssd1 vccd1 vccd1 _06670_ sky130_fd_sc_hd__or2_4
XFILLER_0_24_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12719__A1 net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19013_ clknet_leaf_2_clk img_gen.tracker.next_frame\[451\] net1247 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[451\] sky130_fd_sc_hd__dfrtp_1
X_16225_ obsg2.obstacleArray\[37\] net413 _01903_ net418 vssd1 vssd1 vccd1 vccd1 _01904_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_70_337 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13437_ net235 _07886_ _07887_ net2022 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[507\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_20_clk_A clknet_4_6__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17107__B1 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10649_ ag2.body\[280\] net1237 vssd1 vssd1 vccd1 vccd1 _05622_ sky130_fd_sc_hd__nand2_1
XANTENNA__12952__A net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_428 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16156_ net378 _01834_ _01833_ net347 vssd1 vssd1 vccd1 vccd1 _01835_ sky130_fd_sc_hd__a211o_1
XFILLER_0_80_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13368_ net664 _07860_ vssd1 vssd1 vccd1 vccd1 _07861_ sky130_fd_sc_hd__nor2_1
XFILLER_0_126_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_1396 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15107_ net2602 net145 _01564_ control.body\[900\] vssd1 vssd1 vccd1 vccd1 _00430_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_45_1347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12319_ _07243_ _07244_ vssd1 vssd1 vccd1 vccd1 _07286_ sky130_fd_sc_hd__nor2_1
X_16087_ _01764_ _01765_ net377 vssd1 vssd1 vccd1 vccd1 _01766_ sky130_fd_sc_hd__mux2_1
XANTENNA__15133__A2 net114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10472__A net1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13299_ net671 _07833_ vssd1 vssd1 vccd1 vccd1 _07834_ sky130_fd_sc_hd__nor2_1
XANTENNA__13144__A1 net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_35_clk_A clknet_4_5__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19915_ clknet_leaf_52_clk _00859_ net1368 vssd1 vssd1 vccd1 vccd1 ag2.body\[473\]
+ sky130_fd_sc_hd__dfrtp_4
X_15038_ net2204 net166 _01557_ net2471 vssd1 vssd1 vccd1 vccd1 _00368_ sky130_fd_sc_hd__a22o_1
XFILLER_0_23_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10191__B net1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19846_ clknet_leaf_92_clk _00790_ net1412 vssd1 vssd1 vccd1 vccd1 ag2.body\[548\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_48_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_max_cap509_X net509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16989_ _04018_ net863 net712 ag2.body\[92\] vssd1 vssd1 vccd1 vccd1 _02668_ sky130_fd_sc_hd__o22a_1
XANTENNA__20433__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19777_ clknet_leaf_18_clk _00721_ net1322 vssd1 vssd1 vccd1 vccd1 ag2.body\[623\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__15841__B1 _01644_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09530_ _04489_ _04494_ _04501_ _04502_ vssd1 vssd1 vccd1 vccd1 _04503_ sky130_fd_sc_hd__or4_1
XFILLER_0_64_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_1470 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18728_ clknet_leaf_142_clk img_gen.tracker.next_frame\[166\] net1254 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[166\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_56_1454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09461_ net901 _04432_ net642 vssd1 vssd1 vccd1 vccd1 _04434_ sky130_fd_sc_hd__a21o_1
X_18659_ clknet_leaf_5_clk img_gen.tracker.next_frame\[97\] net1268 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[97\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_52_1307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09392_ sound_gen.osc1.stayCount\[7\] _04345_ net270 vssd1 vssd1 vccd1 vccd1 _04380_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_59_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18138__A2 _03554_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12846__B _07535_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20621_ net1546 vssd1 vssd1 vccd1 vccd1 gpio_oeb[33] sky130_fd_sc_hd__buf_2
XFILLER_0_86_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout141_A net144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_108_clk_A clknet_4_10__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout239_A net240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20552_ clknet_leaf_106_clk _01417_ _00026_ vssd1 vssd1 vccd1 vccd1 sound_gen.osc1.stayCount\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_838 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20483_ clknet_leaf_39_clk _01370_ net1352 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[119\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_6_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10934__X _05907_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout406_A net408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1050_A net1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1148_A net1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13677__B net464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17149__B net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12581__B _07490_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16321__A1 net416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1315_A net1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_3673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16988__B net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_110_3684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15892__B net56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11146__B1 net749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout100 net114 vssd1 vssd1 vccd1 vccd1 net100 sky130_fd_sc_hd__buf_2
XFILLER_0_61_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout396_X net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1109 ag2.x\[1\] vssd1 vssd1 vccd1 vccd1 net1109 sky130_fd_sc_hd__buf_2
XANTENNA__14789__A net997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout775_A _04229_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout111 net112 vssd1 vssd1 vccd1 vccd1 net111 sky130_fd_sc_hd__buf_2
Xfanout122 net128 vssd1 vssd1 vccd1 vccd1 net122 sky130_fd_sc_hd__clkbuf_2
Xfanout133 net135 vssd1 vssd1 vccd1 vccd1 net133 sky130_fd_sc_hd__buf_2
Xfanout144 net219 vssd1 vssd1 vccd1 vccd1 net144 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09890__B _04861_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1103_X net1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout155 net162 vssd1 vssd1 vccd1 vccd1 net155 sky130_fd_sc_hd__buf_2
Xfanout166 net169 vssd1 vssd1 vccd1 vccd1 net166 sky130_fd_sc_hd__buf_2
Xfanout177 net180 vssd1 vssd1 vccd1 vccd1 net177 sky130_fd_sc_hd__buf_2
Xfanout188 net192 vssd1 vssd1 vccd1 vccd1 net188 sky130_fd_sc_hd__buf_2
Xfanout199 net200 vssd1 vssd1 vccd1 vccd1 net199 sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout942_A net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_29_Right_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout563_X net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14635__A1 net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14635__B2 net1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09728_ ag2.body\[92\] net1140 vssd1 vssd1 vccd1 vccd1 _04701_ sky130_fd_sc_hd__nand2_1
XANTENNA__12102__A net1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout54_A net55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12110__A2 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_3488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09659_ net899 net902 net906 vssd1 vssd1 vccd1 vccd1 _04632_ sky130_fd_sc_hd__or3_4
XANTENNA__17612__B net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout730_X net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17585__B1 net698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18973__CLK clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_104_3499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout828_X net828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12670_ net680 _07540_ vssd1 vssd1 vccd1 vccd1 _07541_ sky130_fd_sc_hd__nor2_1
XANTENNA__12756__B _07581_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11621_ obsg2.obstacleArray\[55\] net631 net511 obsg2.obstacleArray\[51\] net508
+ vssd1 vssd1 vccd1 vccd1 _06594_ sky130_fd_sc_hd__o221a_1
XFILLER_0_33_1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_963 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19329__CLK clknet_leaf_103_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14340_ net996 ag2.body\[608\] vssd1 vssd1 vccd1 vccd1 _08501_ sky130_fd_sc_hd__xor2_1
XANTENNA__17888__A1 _08141_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11552_ net1167 net767 vssd1 vssd1 vccd1 vccd1 _06525_ sky130_fd_sc_hd__nor2_1
XFILLER_0_92_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10276__B net1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_38_Right_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10503_ _04446_ _04550_ net892 vssd1 vssd1 vccd1 vccd1 _05476_ sky130_fd_sc_hd__a21o_1
X_14271_ net1008 ag2.body\[15\] vssd1 vssd1 vccd1 vccd1 _08432_ sky130_fd_sc_hd__nand2_1
X_11483_ _06370_ _06398_ _06427_ _06455_ vssd1 vssd1 vccd1 vccd1 _06456_ sky130_fd_sc_hd__and4_1
XFILLER_0_135_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16010_ _01683_ _01688_ vssd1 vssd1 vccd1 vccd1 _01689_ sky130_fd_sc_hd__nand2_1
XANTENNA__12177__A2 _07147_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13374__A1 net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10434_ net1058 control.body\[935\] vssd1 vssd1 vccd1 vccd1 _05407_ sky130_fd_sc_hd__nor2_1
X_13222_ img_gen.tracker.frame\[379\] net658 vssd1 vssd1 vccd1 vccd1 _07801_ sky130_fd_sc_hd__and2_1
XFILLER_0_27_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10188__A1 net912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12491__B _07439_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19479__CLK clknet_leaf_111_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11388__A net1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11924__A2 net623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13153_ net231 _07767_ _07768_ net2001 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[342\]
+ sky130_fd_sc_hd__a22o_1
X_10365_ net1201 control.body\[761\] vssd1 vssd1 vccd1 vccd1 _05338_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_81_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12104_ img_gen.tracker.frame\[360\] net628 net575 _07075_ vssd1 vssd1 vccd1 vccd1
+ _07076_ sky130_fd_sc_hd__a211o_1
X_17961_ _03540_ _03585_ vssd1 vssd1 vccd1 vccd1 _03586_ sky130_fd_sc_hd__and2_1
X_13084_ net243 _07734_ _07735_ net1704 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[306\]
+ sky130_fd_sc_hd__a22o_1
X_10296_ ag2.body\[328\] net788 net1142 _04116_ _05268_ vssd1 vssd1 vccd1 vccd1 _05269_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_40_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19700_ clknet_leaf_136_clk _00644_ net1302 vssd1 vssd1 vccd1 vccd1 control.body\[690\]
+ sky130_fd_sc_hd__dfrtp_1
X_12035_ img_gen.tracker.frame\[36\] net630 net566 _07006_ vssd1 vssd1 vccd1 vccd1
+ _07007_ sky130_fd_sc_hd__a211oi_1
X_16912_ ag2.body\[565\] net705 net689 ag2.body\[567\] _02590_ vssd1 vssd1 vccd1 vccd1
+ _02591_ sky130_fd_sc_hd__a221o_1
XFILLER_0_79_1421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17892_ net516 _03530_ vssd1 vssd1 vccd1 vccd1 _03532_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_47_Right_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16843_ ag2.body\[170\] net862 vssd1 vssd1 vccd1 vccd1 _02522_ sky130_fd_sc_hd__nand2_1
XANTENNA__16615__A2 net449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19631_ clknet_leaf_123_clk _00575_ net1406 vssd1 vssd1 vccd1 vccd1 control.body\[765\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__14849__D _01519_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10360__A1 ag2.body\[294\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15823__B1 _01643_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19562_ clknet_leaf_116_clk _00506_ net1387 vssd1 vssd1 vccd1 vccd1 control.body\[824\]
+ sky130_fd_sc_hd__dfrtp_1
X_16774_ obsg2.obstacleArray\[30\] net488 net496 vssd1 vssd1 vccd1 vccd1 _02453_ sky130_fd_sc_hd__a21o_1
XANTENNA__12012__A net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13986_ ag2.body\[123\] net214 _08159_ ag2.body\[115\] vssd1 vssd1 vccd1 vccd1 _00204_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_88_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12101__A2 net610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18513_ net1513 net1506 vssd1 vssd1 vccd1 vccd1 _00044_ sky130_fd_sc_hd__or2_1
X_15725_ ag2.body\[354\] net197 _01632_ ag2.body\[346\] vssd1 vssd1 vccd1 vccd1 _00980_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_92_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19493_ clknet_leaf_113_clk _00437_ net1399 vssd1 vssd1 vccd1 vccd1 control.body\[899\]
+ sky130_fd_sc_hd__dfrtp_1
X_12937_ net246 _07665_ _07666_ net1803 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[228\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12947__A net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11851__A _06724_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17040__A2 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18444_ _04696_ _04791_ _03831_ vssd1 vssd1 vccd1 vccd1 _03933_ sky130_fd_sc_hd__a21oi_1
X_15656_ ag2.body\[421\] net139 _01624_ ag2.body\[413\] vssd1 vssd1 vccd1 vccd1 _00919_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__20586__D net2301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__20367__RESET_B net1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12868_ net261 _07634_ _07635_ net1614 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[190\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_87_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14607_ _08765_ _08766_ _08767_ _08764_ vssd1 vssd1 vccd1 vccd1 _08768_ sky130_fd_sc_hd__a211o_1
X_18375_ track.nextHighScore\[1\] _03818_ vssd1 vssd1 vccd1 vccd1 _03866_ sky130_fd_sc_hd__xor2_1
X_11819_ img_gen.tracker.frame\[386\] net618 net546 img_gen.tracker.frame\[392\] vssd1
+ vssd1 vccd1 vccd1 _06791_ sky130_fd_sc_hd__o22a_1
X_15587_ ag2.body\[487\] net130 _01617_ ag2.body\[479\] vssd1 vssd1 vccd1 vccd1 _00857_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_7_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10467__A net1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12799_ net253 _07601_ _07602_ net2005 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[154\]
+ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_56_Right_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17326_ net1044 net882 vssd1 vssd1 vccd1 vccd1 _03005_ sky130_fd_sc_hd__xor2_1
X_14538_ _08688_ _08693_ _08698_ vssd1 vssd1 vccd1 vccd1 _08699_ sky130_fd_sc_hd__or3b_1
XFILLER_0_71_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10186__B net1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_133_4374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17257_ ag2.body\[545\] net735 net849 _04201_ _02929_ vssd1 vssd1 vccd1 vccd1 _02936_
+ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_133_4385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14469_ net1020 ag2.body\[270\] vssd1 vssd1 vccd1 vccd1 _08630_ sky130_fd_sc_hd__nand2_1
XANTENNA__12682__A net307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16208_ _01813_ _01886_ _01723_ vssd1 vssd1 vccd1 vccd1 _01887_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_12_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13365__A1 net249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12168__A2 net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09569__B1 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10179__A1 _04427_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17188_ ag2.body\[568\] net881 vssd1 vssd1 vccd1 vccd1 _02867_ sky130_fd_sc_hd__xnor2_1
XANTENNA__11376__B1 net1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10914__B net1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17726__S1 net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11915__A2 net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11298__A net1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16139_ _01698_ _01816_ vssd1 vssd1 vccd1 vccd1 _01818_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_80_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_1189 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18846__CLK clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08961_ ag2.body\[39\] vssd1 vssd1 vccd1 vccd1 _03986_ sky130_fd_sc_hd__inv_2
XFILLER_0_23_1431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_65_Right_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14402__A net990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_1996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_127_4189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19829_ clknet_leaf_124_clk _00773_ net1407 vssd1 vssd1 vccd1 vccd1 ag2.body\[563\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_100_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14617__A1 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18996__CLK clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14617__B2 net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout189_A net191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09513_ net1100 control.body\[837\] vssd1 vssd1 vccd1 vccd1 _04486_ sky130_fd_sc_hd__or2_1
XFILLER_0_71_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10103__A1 net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_1430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1098_A net1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09444_ net893 net899 vssd1 vssd1 vccd1 vccd1 _04417_ sky130_fd_sc_hd__or2_4
XFILLER_0_93_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_74_Right_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11480__B net1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09375_ _04367_ _04372_ vssd1 vssd1 vccd1 vccd1 _01416_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout144_X net144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout523_A net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20604_ net1536 vssd1 vssd1 vccd1 vccd1 gpio_oeb[16] sky130_fd_sc_hd__buf_2
XFILLER_0_46_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20535_ clknet_leaf_107_clk _01400_ _00009_ vssd1 vssd1 vccd1 vccd1 sound_gen.osc1.stayCount\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout311_X net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_116_3860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1053_X net1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_116_3871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout409_X net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_3_5_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_3_5_0_clk sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_112_3724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_112_3735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20466_ clknet_leaf_27_clk _01353_ net1340 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[102\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_132_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_112_3746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11906__A2 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17098__A2 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20397_ clknet_leaf_30_clk _01284_ net1338 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[33\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA_fanout1220_X net1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_18_Left_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_83_Right_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10150_ ag2.body\[56\] net1233 vssd1 vssd1 vccd1 vccd1 _05123_ sky130_fd_sc_hd__xor2_1
XFILLER_0_30_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout680_X net680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_987 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout778_X net778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19973__RESET_B net1470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1598 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10081_ net1226 control.body\[792\] vssd1 vssd1 vccd1 vccd1 _05054_ sky130_fd_sc_hd__or2_1
XANTENNA__14312__A net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19902__RESET_B net1464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11655__B net1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout945_X net945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14608__B2 net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15805__B1 _01641_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13840_ net662 net223 vssd1 vssd1 vccd1 vccd1 _08130_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout57_X net57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13771_ img_gen.updater.commands.count\[8\] _07342_ _08061_ _08075_ vssd1 vssd1 vccd1
+ vccd1 _08084_ sky130_fd_sc_hd__nand4_1
X_10983_ net1052 control.body\[759\] vssd1 vssd1 vccd1 vccd1 _05956_ sky130_fd_sc_hd__xor2_1
XANTENNA__10839__X _05812_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12767__A net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_27_Left_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_92_Right_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_84_2871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15510_ ag2.body\[547\] net155 _01608_ ag2.body\[539\] vssd1 vssd1 vccd1 vccd1 _00789_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__17022__A2 net736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_2882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12722_ net683 _07565_ vssd1 vssd1 vccd1 vccd1 _07566_ sky130_fd_sc_hd__nor2_1
XANTENNA__19151__CLK clknet_leaf_51_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16490_ _02075_ _02167_ _02168_ _02166_ vssd1 vssd1 vccd1 vccd1 _02169_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_84_2893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__20460__RESET_B net1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_2292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_2757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_1600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_133_Right_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15441_ ag2.body\[614\] net85 _01600_ ag2.body\[606\] vssd1 vssd1 vccd1 vccd1 _00728_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_80_2768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18719__CLK clknet_leaf_142_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12653_ net289 _07529_ _07530_ net1877 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[80\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__16673__S net392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16781__A1 net380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_2178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11604_ net505 _06575_ _06576_ net760 vssd1 vssd1 vccd1 vccd1 _06577_ sky130_fd_sc_hd__a211o_1
XFILLER_0_108_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18160_ _03595_ net36 vssd1 vssd1 vccd1 vccd1 _03719_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_61_2189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15372_ _05616_ _01581_ vssd1 vssd1 vccd1 vccd1 _01594_ sky130_fd_sc_hd__and2b_2
X_12584_ net250 _07491_ _07492_ net1954 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[49\]
+ sky130_fd_sc_hd__a22o_1
X_17111_ _02784_ _02785_ _02789_ vssd1 vssd1 vccd1 vccd1 _02790_ sky130_fd_sc_hd__or3_4
XFILLER_0_92_281 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14323_ net818 ag2.body\[451\] ag2.body\[452\] net812 vssd1 vssd1 vccd1 vccd1 _08484_
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_25_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18091_ obsg2.obstacleArray\[50\] _03676_ net527 vssd1 vssd1 vccd1 vccd1 _01301_
+ sky130_fd_sc_hd__o21a_1
X_11535_ _06505_ _06507_ _06504_ vssd1 vssd1 vccd1 vccd1 _06508_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_81_977 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_145 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17042_ _02713_ _02715_ _02716_ _02720_ vssd1 vssd1 vccd1 vccd1 _02721_ sky130_fd_sc_hd__and4_1
XFILLER_0_64_1008 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14254_ net1032 ag2.body\[77\] vssd1 vssd1 vccd1 vccd1 _08415_ sky130_fd_sc_hd__xor2_1
X_11466_ _04419_ _06438_ vssd1 vssd1 vccd1 vccd1 _06439_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_2697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_36_Left_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13205_ img_gen.tracker.frame\[370\] net655 vssd1 vssd1 vccd1 vccd1 _07793_ sky130_fd_sc_hd__and2_1
XFILLER_0_110_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10417_ control.body\[1070\] net1087 vssd1 vssd1 vccd1 vccd1 _05390_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_96_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11397_ _06350_ _06351_ _06353_ _06369_ vssd1 vssd1 vccd1 vccd1 _06370_ sky130_fd_sc_hd__o31a_1
X_14185_ _08341_ _08343_ _08345_ _08342_ vssd1 vssd1 vccd1 vccd1 _08346_ sky130_fd_sc_hd__or4b_1
XFILLER_0_21_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10030__B1 net756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13136_ net2202 net653 vssd1 vssd1 vccd1 vccd1 _07760_ sky130_fd_sc_hd__nand2_1
X_10348_ ag2.body\[289\] net1210 vssd1 vssd1 vccd1 vccd1 _05321_ sky130_fd_sc_hd__or2_1
XFILLER_0_81_1388 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18993_ clknet_leaf_8_clk img_gen.tracker.next_frame\[431\] net1272 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[431\] sky130_fd_sc_hd__dfrtp_1
X_10279_ _05246_ _05249_ _05250_ _05251_ vssd1 vssd1 vccd1 vccd1 _05252_ sky130_fd_sc_hd__or4_1
X_17944_ net957 net539 net537 net460 vssd1 vssd1 vccd1 vccd1 _03573_ sky130_fd_sc_hd__and4_1
X_13067_ net246 _07726_ _07727_ net1861 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[297\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_40_1041 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1440 net1442 vssd1 vssd1 vccd1 vccd1 net1440 sky130_fd_sc_hd__clkbuf_4
X_12018_ net1216 net1191 img_gen.tracker.frame\[225\] vssd1 vssd1 vccd1 vccd1 _06990_
+ sky130_fd_sc_hd__and3_1
X_17875_ img_gen.updater.commands.rR1.rainbowRNG\[14\] _03506_ vssd1 vssd1 vccd1 vccd1
+ _03517_ sky130_fd_sc_hd__or2_1
Xfanout1451 net1452 vssd1 vssd1 vccd1 vccd1 net1451 sky130_fd_sc_hd__clkbuf_2
Xfanout1462 net1465 vssd1 vssd1 vccd1 vccd1 net1462 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_136_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_122_4031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1473 net1477 vssd1 vssd1 vccd1 vccd1 net1473 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_75_1104 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_122_4042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1484 net1493 vssd1 vssd1 vccd1 vccd1 net1484 sky130_fd_sc_hd__buf_2
XFILLER_0_136_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_122_4053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1495 net1504 vssd1 vssd1 vccd1 vccd1 net1495 sky130_fd_sc_hd__clkbuf_4
X_19614_ clknet_leaf_120_clk net2104 net1395 vssd1 vssd1 vccd1 vccd1 control.body\[780\]
+ sky130_fd_sc_hd__dfrtp_1
X_16826_ ag2.body\[229\] net951 vssd1 vssd1 vccd1 vccd1 _02505_ sky130_fd_sc_hd__xor2_1
XFILLER_0_88_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17591__A2_N net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_45_Left_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16757_ net460 _02435_ vssd1 vssd1 vccd1 vccd1 _02436_ sky130_fd_sc_hd__or2_1
X_19545_ clknet_leaf_115_clk _00489_ net1389 vssd1 vssd1 vccd1 vccd1 control.body\[855\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__17252__B net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12086__A1 net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17549__B1 net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13969_ ag2.body\[108\] net202 _08157_ ag2.body\[100\] vssd1 vssd1 vccd1 vccd1 _00189_
+ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_139_clk clknet_4_2__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_139_clk
+ sky130_fd_sc_hd__clkbuf_8
X_15708_ ag2.body\[372\] net140 _01629_ ag2.body\[364\] vssd1 vssd1 vccd1 vccd1 _00966_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_88_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16688_ net360 _02289_ _02366_ _02228_ vssd1 vssd1 vccd1 vccd1 _02367_ sky130_fd_sc_hd__o211a_1
XFILLER_0_88_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19476_ clknet_leaf_109_clk _00420_ net1416 vssd1 vssd1 vccd1 vccd1 control.body\[914\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15639_ ag2.body\[438\] net126 _01622_ ag2.body\[430\] vssd1 vssd1 vccd1 vccd1 _00904_
+ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_100_Right_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18427_ _03800_ _03915_ _03799_ vssd1 vssd1 vccd1 vccd1 _03916_ sky130_fd_sc_hd__o21a_1
XFILLER_0_31_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15575__A2 net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20130__RESET_B net1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_135_4436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_135_4447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09160_ ag2.body\[506\] vssd1 vssd1 vccd1 vccd1 _04185_ sky130_fd_sc_hd__inv_2
XFILLER_0_5_1277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_44_1653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18358_ _03795_ _03852_ _03794_ vssd1 vssd1 vccd1 vccd1 _03853_ sky130_fd_sc_hd__o21ba_1
XTAP_TAPCELL_ROW_44_1664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09986__A net1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17309_ ag2.body\[399\] net931 vssd1 vssd1 vccd1 vccd1 _02988_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_20_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_884 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09091_ ag2.body\[332\] vssd1 vssd1 vccd1 vccd1 _04116_ sky130_fd_sc_hd__inv_2
XANTENNA__18525__RESET_B net1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18289_ track.nextHighScore\[6\] _03782_ _03784_ track.nextHighScore\[7\] vssd1 vssd1
+ vccd1 vccd1 _03785_ sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_25_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10925__A net1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09718__A1_N net770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_54_Left_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20320_ clknet_leaf_43_clk _01216_ net1378 vssd1 vssd1 vccd1 vccd1 obsg2.randCord\[5\]
+ sky130_fd_sc_hd__dfstp_2
XFILLER_0_86_1277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19794__CLK clknet_leaf_127_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_1565 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold901 control.body\[915\] vssd1 vssd1 vccd1 vccd1 net2463 sky130_fd_sc_hd__dlygate4sd3_1
Xhold912 control.body\[939\] vssd1 vssd1 vccd1 vccd1 net2474 sky130_fd_sc_hd__dlygate4sd3_1
X_20251_ clknet_leaf_70_clk _01195_ net1497 vssd1 vssd1 vccd1 vccd1 ag2.body\[137\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_114_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13020__B _07532_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold923 control.body\[1082\] vssd1 vssd1 vccd1 vccd1 net2485 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_90_3053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold934 control.body\[679\] vssd1 vssd1 vccd1 vccd1 net2496 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12010__B2 net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_3064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout104_A net114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold945 control.body\[784\] vssd1 vssd1 vccd1 vccd1 net2507 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_90_3075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold956 control.body\[821\] vssd1 vssd1 vccd1 vccd1 net2518 sky130_fd_sc_hd__dlygate4sd3_1
Xhold967 control.body\[879\] vssd1 vssd1 vccd1 vccd1 net2529 sky130_fd_sc_hd__dlygate4sd3_1
X_20182_ clknet_leaf_87_clk _01126_ net1460 vssd1 vssd1 vccd1 vccd1 ag2.body\[212\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_12_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold978 control.body\[1037\] vssd1 vssd1 vccd1 vccd1 net2540 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1131 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold989 control.body\[818\] vssd1 vssd1 vccd1 vccd1 net2551 sky130_fd_sc_hd__dlygate4sd3_1
X_09993_ net1193 _04240_ control.body\[732\] net758 vssd1 vssd1 vccd1 vccd1 _04966_
+ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_38_1468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08944_ net1040 vssd1 vssd1 vccd1 vccd1 _03969_ sky130_fd_sc_hd__inv_2
XFILLER_0_99_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14132__A net1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1013_A net1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09714__B1 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20001__CLK clknet_leaf_66_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11475__B net1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17788__B1 net1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout473_A _06647_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19174__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_3403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17162__B net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_3414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10659__X _05632_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout261_X net261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout738_A _04262_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1382_A net1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout359_X net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11491__A net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12172__S1 net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20151__CLK clknet_leaf_98_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09427_ net1712 _04399_ _04400_ net1726 vssd1 vssd1 vccd1 vccd1 _00003_ sky130_fd_sc_hd__a22o_1
XANTENNA__16209__D net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1170_X net1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout905_A net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_118_3911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_3922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_3933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09358_ sound_gen.osc1.stayCount\[16\] _04358_ vssd1 vssd1 vccd1 vccd1 _04360_ sky130_fd_sc_hd__and2_1
XFILLER_0_81_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_114_3808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11052__A2 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16515__A1 net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09289_ _04309_ vssd1 vssd1 vccd1 vccd1 sound_gen.osc1.freq_nxt\[0\] sky130_fd_sc_hd__inv_2
XFILLER_0_69_1464 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14307__A net1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1435_X net1435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_871 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11320_ ag2.body\[557\] net1101 vssd1 vssd1 vccd1 vccd1 _06293_ sky130_fd_sc_hd__xor2_1
X_20518_ clknet_leaf_112_clk track.nextCurrScore\[0\] net1424 vssd1 vssd1 vccd1 vccd1
+ control.body_update.curr_length\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout895_X net895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18268__A1 net319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11251_ _06211_ _06212_ _06213_ _06214_ vssd1 vssd1 vccd1 vccd1 _06224_ sky130_fd_sc_hd__a22o_1
X_20449_ clknet_leaf_41_clk _01336_ net1371 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[85\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__09548__A3 _04446_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_2550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10202_ _05168_ _05169_ _05173_ _05174_ vssd1 vssd1 vccd1 vccd1 _05175_ sky130_fd_sc_hd__or4_1
XFILLER_0_43_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16818__A2 net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11182_ net1056 ag2.body\[183\] vssd1 vssd1 vccd1 vccd1 _06155_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_73_2561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11986__S1 net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14829__A1 _08650_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11760__B1 net542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10133_ net1049 control.body\[823\] vssd1 vssd1 vccd1 vccd1 _05106_ sky130_fd_sc_hd__nand2_1
XANTENNA__11666__A net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15990_ _01667_ _01668_ _01669_ vssd1 vssd1 vccd1 vccd1 _01673_ sky130_fd_sc_hd__a21o_1
XANTENNA__17491__A2 net718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10570__A net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10064_ net1170 control.body\[714\] vssd1 vssd1 vccd1 vccd1 _05037_ sky130_fd_sc_hd__xor2_1
X_14941_ net2252 net173 _01545_ net2340 vssd1 vssd1 vccd1 vccd1 _00283_ sky130_fd_sc_hd__a22o_1
XANTENNA__17779__B1 net530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17660_ ag2.body\[110\] net944 vssd1 vssd1 vccd1 vccd1 _03339_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_86_2933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14872_ net2142 net181 _01537_ control.body\[1108\] vssd1 vssd1 vccd1 vccd1 _00222_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__08975__A ag2.body\[66\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18168__B net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16611_ obsg2.obstacleArray\[88\] obsg2.obstacleArray\[89\] net445 vssd1 vssd1 vccd1
+ vccd1 _02290_ sky130_fd_sc_hd__mux2_1
X_13823_ _08119_ vssd1 vssd1 vccd1 vccd1 _08120_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_67_2354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17072__B net848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_2819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17591_ ag2.body\[59\] net716 net698 ag2.body\[62\] vssd1 vssd1 vccd1 vccd1 _03270_
+ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_67_2365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12497__A net388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13804__A2 _06505_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_2376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10079__B1 _04587_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16542_ net498 _02219_ vssd1 vssd1 vccd1 vccd1 _02221_ sky130_fd_sc_hd__or2_1
X_19330_ clknet_leaf_100_clk _00274_ net1443 vssd1 vssd1 vccd1 vccd1 control.body\[1056\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_97_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13754_ img_gen.updater.commands.count\[3\] _08068_ vssd1 vssd1 vccd1 vccd1 _08072_
+ sky130_fd_sc_hd__or2_1
XANTENNA__11815__A1 net568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10966_ net1134 control.body\[1004\] vssd1 vssd1 vccd1 vccd1 _05939_ sky130_fd_sc_hd__nor2_1
X_19261_ clknet_leaf_73_clk _00205_ net1500 vssd1 vssd1 vccd1 vccd1 ag2.body\[124\]
+ sky130_fd_sc_hd__dfrtp_4
X_12705_ net2107 net647 _07556_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[106\]
+ sky130_fd_sc_hd__and3_1
X_16473_ _02150_ _02151_ _02148_ vssd1 vssd1 vccd1 vccd1 _02152_ sky130_fd_sc_hd__o21a_1
XANTENNA__13105__B _07575_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15557__A2 net187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13685_ net902 net434 _08027_ _08022_ vssd1 vssd1 vccd1 vccd1 track.nextCurrScore\[5\]
+ sky130_fd_sc_hd__a22o_1
X_10897_ _04237_ net904 _04554_ _05075_ _04573_ vssd1 vssd1 vccd1 vccd1 _05870_ sky130_fd_sc_hd__a41o_1
XFILLER_0_122_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18212_ _03654_ net40 vssd1 vssd1 vccd1 vccd1 _03745_ sky130_fd_sc_hd__nor2_1
XFILLER_0_39_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_14_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15424_ control.body\[631\] net84 _01598_ ag2.body\[623\] vssd1 vssd1 vccd1 vccd1
+ _00713_ sky130_fd_sc_hd__a22o_1
X_19192_ clknet_leaf_53_clk _00136_ net1365 vssd1 vssd1 vccd1 vccd1 ag2.body\[55\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_14_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12636_ net241 _07520_ _07521_ net1804 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[72\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_127_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_130_4300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18143_ net518 _03710_ vssd1 vssd1 vccd1 vccd1 _01319_ sky130_fd_sc_hd__nor2_1
XFILLER_0_5_518 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15355_ control.body\[680\] net75 _01592_ net2542 vssd1 vssd1 vccd1 vccd1 _00650_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11043__A2 net477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12567_ net439 net470 _07452_ vssd1 vssd1 vccd1 vccd1 _07483_ sky130_fd_sc_hd__or3_4
XFILLER_0_48_1515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16135__C _01691_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13121__A net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14306_ _08463_ _08464_ _08466_ vssd1 vssd1 vccd1 vccd1 _08467_ sky130_fd_sc_hd__or3_2
X_18074_ obsg2.obstacleArray\[44\] _03665_ net520 vssd1 vssd1 vccd1 vccd1 _01295_
+ sky130_fd_sc_hd__o21a_1
X_11518_ net1152 net1222 vssd1 vssd1 vccd1 vccd1 _06491_ sky130_fd_sc_hd__and2b_1
XFILLER_0_124_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15286_ control.body\[747\] net87 _01584_ control.body\[739\] vssd1 vssd1 vccd1 vccd1
+ _00589_ sky130_fd_sc_hd__a22o_1
XFILLER_0_125_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12498_ _06724_ net337 vssd1 vssd1 vccd1 vccd1 _07444_ sky130_fd_sc_hd__nor2_4
XANTENNA__19047__CLK clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold208 img_gen.tracker.frame\[121\] vssd1 vssd1 vccd1 vccd1 net1770 sky130_fd_sc_hd__dlygate4sd3_1
X_17025_ ag2.body\[401\] net877 vssd1 vssd1 vccd1 vccd1 _02704_ sky130_fd_sc_hd__xor2_1
Xhold219 img_gen.tracker.frame\[179\] vssd1 vssd1 vccd1 vccd1 net1781 sky130_fd_sc_hd__dlygate4sd3_1
X_14237_ net836 ag2.body\[481\] _04174_ net980 vssd1 vssd1 vccd1 vccd1 _08398_ sky130_fd_sc_hd__a22o_1
X_11449_ net1087 control.body\[958\] vssd1 vssd1 vccd1 vccd1 _06422_ sky130_fd_sc_hd__xor2_1
XFILLER_0_111_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16809__A2 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14168_ net841 ag2.body\[200\] _04067_ net1007 vssd1 vssd1 vccd1 vccd1 _08329_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_128_4240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11751__B1 _06722_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_52_1900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13119_ net265 _07750_ _07751_ net1661 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[325\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__15048__A _06413_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17482__A2 net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_124_4104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19197__CLK clknet_leaf_53_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18976_ clknet_leaf_7_clk img_gen.tracker.next_frame\[414\] net1265 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[414\] sky130_fd_sc_hd__dfrtp_1
X_14099_ net979 ag2.body\[586\] vssd1 vssd1 vccd1 vccd1 _08260_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_124_4115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17927_ net318 _03559_ obsg2.obstacleArray\[3\] vssd1 vssd1 vccd1 vccd1 _03560_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_33_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1270 net1272 vssd1 vssd1 vccd1 vccd1 net1270 sky130_fd_sc_hd__clkbuf_4
XANTENNA__17234__A2 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout1281 net1283 vssd1 vssd1 vccd1 vccd1 net1281 sky130_fd_sc_hd__clkbuf_4
XANTENNA__20382__RESET_B net1374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17858_ net2467 _03509_ _03511_ vssd1 vssd1 vccd1 vccd1 _01233_ sky130_fd_sc_hd__o21ba_1
Xfanout1292 net1293 vssd1 vssd1 vccd1 vccd1 net1292 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_55_1508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_1568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16809_ ag2.body\[67\] net720 net935 _04002_ vssd1 vssd1 vccd1 vccd1 _02488_ sky130_fd_sc_hd__o22a_1
XFILLER_0_117_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17789_ _03463_ _03464_ _03465_ vssd1 vssd1 vccd1 vccd1 _01211_ sky130_fd_sc_hd__and3b_1
XFILLER_0_132_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_137_4509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_1266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19528_ clknet_leaf_120_clk _00472_ net1394 vssd1 vssd1 vccd1 vccd1 control.body\[870\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_49_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12200__A net480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_46_1726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_1411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19459_ clknet_leaf_110_clk _00403_ net1417 vssd1 vssd1 vccd1 vccd1 control.body\[929\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_27_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18094__A net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17942__B1 obsg2.obstacleArray\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_1298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09212_ net900 vssd1 vssd1 vccd1 vccd1 _04237_ sky130_fd_sc_hd__inv_2
XFILLER_0_70_1590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_1552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_96_3240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_62_Left_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16326__B net406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_96_3251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09143_ ag2.body\[473\] vssd1 vssd1 vccd1 vccd1 _04168_ sky130_fd_sc_hd__inv_2
XFILLER_0_16_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_3262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_92_3115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_92_3126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12573__C net440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13031__A net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09074_ ag2.body\[300\] vssd1 vssd1 vccd1 vccd1 _04099_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_92_3137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_1074 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20303_ clknet_leaf_37_clk net1569 net1349 vssd1 vssd1 vccd1 vccd1 control.divider.detect.signal
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_130_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11990__B1 net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_1373 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold720 _00407_ vssd1 vssd1 vccd1 vccd1 net2282 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1130_A net1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout107_X net107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold731 control.body\[1065\] vssd1 vssd1 vccd1 vccd1 net2293 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1228_A net1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold742 _00287_ vssd1 vssd1 vccd1 vccd1 net2304 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20234_ clknet_leaf_69_clk _01178_ net1496 vssd1 vssd1 vccd1 vccd1 ag2.body\[152\]
+ sky130_fd_sc_hd__dfrtp_4
Xhold753 control.body\[645\] vssd1 vssd1 vccd1 vccd1 net2315 sky130_fd_sc_hd__dlygate4sd3_1
Xhold764 control.body\[873\] vssd1 vssd1 vccd1 vccd1 net2326 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout590_A net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold775 _00660_ vssd1 vssd1 vccd1 vccd1 net2337 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout688_A net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold786 sound_gen.osc1.count\[1\] vssd1 vssd1 vccd1 vccd1 net2348 sky130_fd_sc_hd__dlygate4sd3_1
Xhold797 _00417_ vssd1 vssd1 vccd1 vccd1 net2359 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10390__A net1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20165_ clknet_leaf_82_clk _01109_ net1484 vssd1 vssd1 vccd1 vccd1 ag2.body\[227\]
+ sky130_fd_sc_hd__dfrtp_4
X_09976_ net1137 control.body\[1116\] vssd1 vssd1 vccd1 vccd1 _04949_ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout1016_X net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_71_Left_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16996__B net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_3601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_1479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20096_ clknet_leaf_78_clk _01040_ net1490 vssd1 vssd1 vccd1 vccd1 ag2.body\[302\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_77_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout855_A net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18564__CLK clknet_leaf_15_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17225__A2 net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18422__A1 track.nextHighScore\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1012 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16433__B1 net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11933__B net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20052__RESET_B net1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout643_X net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10820_ net751 control.body\[1094\] control.body\[1093\] net755 vssd1 vssd1 vccd1
+ vccd1 _05793_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_95_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10549__B net1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20100__Q ag2.body\[290\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout810_X net810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10751_ _05698_ _05703_ _05710_ _05723_ _04687_ vssd1 vssd1 vccd1 vccd1 _05724_ sky130_fd_sc_hd__o32a_1
XANTENNA__15539__A2 net161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout908_X net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_125 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_968 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13470_ _07592_ net304 vssd1 vssd1 vccd1 vccd1 _07900_ sky130_fd_sc_hd__nor2_1
X_10682_ ag2.body\[347\] net1163 vssd1 vssd1 vccd1 vccd1 _05655_ sky130_fd_sc_hd__xor2_1
XANTENNA__10563__A_N net1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12421_ net549 _07380_ _07381_ _07382_ vssd1 vssd1 vccd1 vccd1 _07383_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_124_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_2601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15140_ net2429 net105 _01567_ control.body\[866\] vssd1 vssd1 vccd1 vccd1 _00460_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_129_1159 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_2612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12352_ net248 _07318_ vssd1 vssd1 vccd1 vccd1 _07319_ sky130_fd_sc_hd__and2_2
XFILLER_0_69_1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10284__B net1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_2623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11303_ _06268_ _06270_ _06272_ _06273_ vssd1 vssd1 vccd1 vccd1 _06276_ sky130_fd_sc_hd__or4_2
XTAP_TAPCELL_ROW_56_2022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15071_ net2354 net150 _01560_ net2536 vssd1 vssd1 vccd1 vccd1 _00398_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_56_2033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14324__X _08485_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12283_ _04273_ _07241_ _07248_ _07252_ vssd1 vssd1 vccd1 vccd1 _07253_ sky130_fd_sc_hd__o2bb2a_2
XANTENNA__12780__A net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_2044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09926__B1 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14022_ net1026 ag2.body\[29\] vssd1 vssd1 vccd1 vccd1 _08183_ sky130_fd_sc_hd__xor2_1
XANTENNA__11667__Y _06639_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11234_ _04695_ _05051_ net636 vssd1 vssd1 vccd1 vccd1 _06207_ sky130_fd_sc_hd__o21ai_2
XANTENNA__17067__B net880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18907__CLK clknet_leaf_144_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11396__A _04573_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18830_ clknet_leaf_141_clk img_gen.tracker.next_frame\[268\] net1262 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[268\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_8_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11165_ net900 net921 _04554_ _05223_ vssd1 vssd1 vccd1 vccd1 _06138_ sky130_fd_sc_hd__a31oi_2
XFILLER_0_101_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_8_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10116_ net1119 control.body\[708\] vssd1 vssd1 vccd1 vccd1 _05089_ sky130_fd_sc_hd__or2_1
X_11096_ ag2.body\[426\] net1176 vssd1 vssd1 vccd1 vccd1 _06069_ sky130_fd_sc_hd__nand2_1
X_15973_ net223 _08118_ net663 vssd1 vssd1 vccd1 vccd1 _01659_ sky130_fd_sc_hd__o21ai_1
X_18761_ clknet_leaf_16_clk img_gen.tracker.next_frame\[199\] net1315 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[199\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__16398__S net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_2416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_2427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17712_ net360 _03390_ _03389_ net358 vssd1 vssd1 vccd1 vccd1 _03391_ sky130_fd_sc_hd__o211a_1
X_10047_ _05016_ _05017_ _05018_ _05019_ vssd1 vssd1 vccd1 vccd1 _05020_ sky130_fd_sc_hd__or4_1
X_14924_ control.body\[1066\] net170 _01543_ control.body\[1058\] vssd1 vssd1 vccd1
+ vccd1 _00268_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_69_2438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18692_ clknet_leaf_28_clk img_gen.tracker.next_frame\[130\] net1336 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[130\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__12498__Y _07444_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold80 img_gen.tracker.frame\[196\] vssd1 vssd1 vccd1 vccd1 net1642 sky130_fd_sc_hd__dlygate4sd3_1
Xhold91 img_gen.tracker.frame\[278\] vssd1 vssd1 vccd1 vccd1 net1653 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17643_ _03317_ _03318_ _03319_ _03321_ vssd1 vssd1 vccd1 vccd1 _03322_ sky130_fd_sc_hd__a211o_1
X_14855_ _08355_ _08358_ _08673_ vssd1 vssd1 vccd1 vccd1 _01526_ sky130_fd_sc_hd__o21a_1
XANTENNA__15778__A2 net210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17811__A net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13116__A _07581_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13806_ net1144 _08105_ vssd1 vssd1 vccd1 vccd1 _08107_ sky130_fd_sc_hd__nand2_1
X_17574_ _04119_ net876 net966 _04120_ _03252_ vssd1 vssd1 vccd1 vccd1 _03253_ sky130_fd_sc_hd__o221a_1
XFILLER_0_19_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14786_ net991 _04200_ ag2.body\[550\] net804 vssd1 vssd1 vccd1 vccd1 _01457_ sky130_fd_sc_hd__o22a_1
XFILLER_0_118_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11998_ net560 _06966_ _06969_ vssd1 vssd1 vccd1 vccd1 _06970_ sky130_fd_sc_hd__a21o_1
XANTENNA__09457__A2 _04238_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10459__B net1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16525_ net956 net536 _02052_ vssd1 vssd1 vccd1 vccd1 _02204_ sky130_fd_sc_hd__or3_1
XFILLER_0_9_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19313_ clknet_leaf_99_clk _00257_ net1445 vssd1 vssd1 vccd1 vccd1 control.body\[1087\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13737_ _04272_ img_gen.updater.commands.cmd_num\[2\] _07225_ _07247_ img_gen.updater.commands.mode\[0\]
+ vssd1 vssd1 vccd1 vccd1 _08058_ sky130_fd_sc_hd__a311oi_1
XFILLER_0_58_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17530__B net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10949_ _05920_ _05921_ vssd1 vssd1 vccd1 vccd1 _05922_ sky130_fd_sc_hd__and2b_1
XFILLER_0_15_1547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_70_clk clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_70_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_133_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16456_ _02057_ _02134_ vssd1 vssd1 vccd1 vccd1 _02135_ sky130_fd_sc_hd__nor2_1
X_19244_ clknet_leaf_76_clk _00188_ net1481 vssd1 vssd1 vccd1 vccd1 ag2.body\[107\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__09600__Y _04573_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13668_ _08016_ _08017_ _08018_ vssd1 vssd1 vccd1 vccd1 obsrand1.next_randY\[3\]
+ sky130_fd_sc_hd__and3_1
XFILLER_0_2_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_22_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12674__B net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_827 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15407_ _04574_ net52 vssd1 vssd1 vccd1 vccd1 _01597_ sky130_fd_sc_hd__nor2_2
X_19175_ clknet_leaf_21_clk _00119_ net1363 vssd1 vssd1 vccd1 vccd1 ag2.body\[38\]
+ sky130_fd_sc_hd__dfrtp_4
X_12619_ _06639_ net440 net569 net554 vssd1 vssd1 vccd1 vccd1 _07511_ sky130_fd_sc_hd__and4_1
X_16387_ net497 _02061_ vssd1 vssd1 vccd1 vccd1 _02066_ sky130_fd_sc_hd__and2_1
XFILLER_0_27_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13599_ _03960_ control.divider.count\[16\] _07972_ _07973_ vssd1 vssd1 vccd1 vccd1
+ _07974_ sky130_fd_sc_hd__a211o_1
XFILLER_0_5_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18126_ _01714_ net345 net300 vssd1 vssd1 vccd1 vccd1 _03699_ sky130_fd_sc_hd__and3_1
X_15338_ control.body\[697\] net71 _01590_ control.body\[689\] vssd1 vssd1 vccd1 vccd1
+ _00635_ sky130_fd_sc_hd__a22o_1
XFILLER_0_112_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10194__B net1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11972__B1 net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18057_ net301 _03574_ vssd1 vssd1 vccd1 vccd1 _03654_ sky130_fd_sc_hd__nand2_1
XFILLER_0_48_1367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15269_ control.body\[764\] net108 _01582_ net2422 vssd1 vssd1 vccd1 vccd1 _00574_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_125_1535 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_846 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17008_ _04180_ net874 net692 ag2.body\[503\] _02686_ vssd1 vssd1 vccd1 vccd1 _02687_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_65_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09917__B1 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_1534 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_1405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11724__B1 net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout507 net508 vssd1 vssd1 vccd1 vccd1 net507 sky130_fd_sc_hd__clkbuf_4
X_09830_ net1229 control.body\[920\] vssd1 vssd1 vccd1 vccd1 _04803_ sky130_fd_sc_hd__nand2_1
XFILLER_0_10_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_6_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout518 net519 vssd1 vssd1 vccd1 vccd1 net518 sky130_fd_sc_hd__clkbuf_2
Xfanout529 net530 vssd1 vssd1 vccd1 vccd1 net529 sky130_fd_sc_hd__clkbuf_2
X_09761_ ag2.body\[209\] net1210 vssd1 vssd1 vccd1 vccd1 _04734_ sky130_fd_sc_hd__xor2_1
X_18959_ clknet_leaf_7_clk img_gen.tracker.next_frame\[397\] net1268 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[397\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__16101__S net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14410__A net1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09692_ ag2.body\[65\] net1208 vssd1 vssd1 vccd1 vccd1 _04665_ sky130_fd_sc_hd__or2_1
XFILLER_0_119_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout171_A net183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13026__A net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12568__C net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1040 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16179__C1 net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_3302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_98_3313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12865__A net383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1080_A net1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_61_clk clknet_4_13__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_61_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_98_3324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout436_A net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1178_A net1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16194__A2 net430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1068 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout603_A net605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13401__B1 net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15941__A2 net195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1345_A net1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09126_ ag2.body\[426\] vssd1 vssd1 vccd1 vccd1 _04151_ sky130_fd_sc_hd__inv_2
XANTENNA__19362__CLK clknet_leaf_102_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11963__B1 net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1456 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17694__A2 net734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09893__B net1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09057_ ag2.body\[251\] vssd1 vssd1 vccd1 vccd1 _04082_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout1133_X net1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold550 img_gen.tracker.frame\[518\] vssd1 vssd1 vccd1 vccd1 net2112 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10391__Y _05364_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout972_A net974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10832__B net1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout593_X net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold561 control.body\[1113\] vssd1 vssd1 vccd1 vccd1 net2123 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1022 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold572 img_gen.tracker.frame\[476\] vssd1 vssd1 vccd1 vccd1 net2134 sky130_fd_sc_hd__dlygate4sd3_1
Xhold583 control.body\[1114\] vssd1 vssd1 vccd1 vccd1 net2145 sky130_fd_sc_hd__dlygate4sd3_1
X_20217_ clknet_leaf_60_clk _01161_ net1466 vssd1 vssd1 vccd1 vccd1 ag2.body\[183\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__09534__A1_N net787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold594 img_gen.tracker.frame\[573\] vssd1 vssd1 vccd1 vccd1 net2156 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16800__A net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20148_ clknet_leaf_98_clk _01092_ net1444 vssd1 vssd1 vccd1 vccd1 ag2.body\[242\]
+ sky130_fd_sc_hd__dfrtp_4
X_09959_ ag2.body\[81\] net1211 vssd1 vssd1 vccd1 vccd1 _04932_ sky130_fd_sc_hd__xor2_1
XANTENNA_fanout760_X net760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17615__B net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout858_X net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15416__A _05685_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20079_ clknet_leaf_76_clk _01023_ net1492 vssd1 vssd1 vccd1 vccd1 ag2.body\[317\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_77_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12970_ net668 _07681_ vssd1 vssd1 vccd1 vccd1 _07682_ sky130_fd_sc_hd__nor2_1
XANTENNA__14320__A net1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11663__B net1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11921_ img_gen.tracker.frame\[313\] img_gen.tracker.frame\[316\] img_gen.tracker.frame\[319\]
+ img_gen.tracker.frame\[322\] net1225 net1191 vssd1 vssd1 vccd1 vccd1 _06893_ sky130_fd_sc_hd__mux4_1
XANTENNA__16957__A1 ag2.body\[294\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12691__A1 net285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16957__B2 ag2.body\[295\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17631__A ag2.body\[165\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14640_ _08797_ _08799_ _08800_ vssd1 vssd1 vccd1 vccd1 _08801_ sky130_fd_sc_hd__or3_1
XANTENNA__15703__X _01629_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14968__B1 net51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11852_ net385 _06820_ net382 _06724_ vssd1 vssd1 vccd1 vccd1 _06824_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_16_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_16_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14974__B net54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10803_ ag2.body\[32\] net1223 vssd1 vssd1 vccd1 vccd1 _05776_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_0_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14571_ _08729_ _08730_ _08731_ vssd1 vssd1 vccd1 vccd1 _08732_ sky130_fd_sc_hd__or3_1
XANTENNA__12443__A1 net625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11783_ img_gen.tracker.frame\[170\] net621 net587 img_gen.tracker.frame\[179\] _06754_
+ vssd1 vssd1 vccd1 vccd1 _06755_ sky130_fd_sc_hd__o221a_1
XFILLER_0_138_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_52_clk clknet_4_6__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_52_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_28_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16310_ obsg2.obstacleArray\[106\] obsg2.obstacleArray\[107\] net405 vssd1 vssd1
+ vccd1 vccd1 _01989_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13522_ net226 _07919_ vssd1 vssd1 vccd1 vccd1 _07920_ sky130_fd_sc_hd__nor2_1
X_17290_ ag2.body\[305\] net736 net729 ag2.body\[306\] vssd1 vssd1 vccd1 vccd1 _02969_
+ sky130_fd_sc_hd__o22a_1
X_10734_ ag2.body\[249\] net780 _05705_ _05706_ _05704_ vssd1 vssd1 vccd1 vccd1 _05707_
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_12_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1483 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14196__A1 net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16241_ obsg2.obstacleArray\[40\] obsg2.obstacleArray\[41\] net404 vssd1 vssd1 vccd1
+ vccd1 _01920_ sky130_fd_sc_hd__mux2_1
XANTENNA__14196__B2 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13453_ net256 _07892_ _07893_ net1657 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[517\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_36_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10665_ net1157 control.body\[883\] vssd1 vssd1 vccd1 vccd1 _05638_ sky130_fd_sc_hd__xor2_1
XANTENNA__18462__A net717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_1610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_2106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_459 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12404_ _07269_ _07274_ _07277_ _07329_ _07347_ vssd1 vssd1 vccd1 vccd1 _07367_ sky130_fd_sc_hd__a2111o_1
X_16172_ obsg2.obstacleArray\[28\] obsg2.obstacleArray\[29\] net428 vssd1 vssd1 vccd1
+ vccd1 _01851_ sky130_fd_sc_hd__mux2_1
XFILLER_0_91_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13384_ net228 _07866_ _07867_ net1637 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[474\]
+ sky130_fd_sc_hd__a22o_1
X_10596_ net1201 control.body\[825\] vssd1 vssd1 vccd1 vccd1 _05569_ sky130_fd_sc_hd__xor2_1
XFILLER_0_2_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15123_ net2634 net104 _01565_ control.body\[883\] vssd1 vssd1 vccd1 vccd1 _00445_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_105_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12335_ _07301_ _06634_ vssd1 vssd1 vccd1 vccd1 _07302_ sky130_fd_sc_hd__and2b_1
XANTENNA__17685__A2 net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19931_ clknet_leaf_47_clk _00875_ net1375 vssd1 vssd1 vccd1 vccd1 ag2.body\[457\]
+ sky130_fd_sc_hd__dfrtp_4
X_15054_ net2375 net164 _01558_ control.body\[949\] vssd1 vssd1 vccd1 vccd1 _00383_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_50_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12266_ img_gen.updater.commands.count\[14\] img_gen.updater.commands.count\[15\]
+ img_gen.updater.commands.count\[13\] img_gen.updater.commands.count\[12\] vssd1
+ vssd1 vccd1 vccd1 _07236_ sky130_fd_sc_hd__or4_1
XFILLER_0_120_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10742__B net1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11706__B1 net551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14005_ net976 ag2.body\[507\] vssd1 vssd1 vccd1 vccd1 _08166_ sky130_fd_sc_hd__xor2_1
XANTENNA__17437__A2 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11217_ net1100 control.body\[845\] vssd1 vssd1 vccd1 vccd1 _06190_ sky130_fd_sc_hd__xnor2_1
X_19862_ clknet_leaf_94_clk _00806_ net1437 vssd1 vssd1 vccd1 vccd1 ag2.body\[532\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_120_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12015__A _06986_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12197_ _07165_ _07168_ vssd1 vssd1 vccd1 vccd1 _07169_ sky130_fd_sc_hd__nor2_2
XFILLER_0_43_1286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_1443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18813_ clknet_leaf_3_clk img_gen.tracker.next_frame\[251\] net1259 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[251\] sky130_fd_sc_hd__dfrtp_1
X_11148_ _06111_ _06113_ _06116_ _06120_ _06109_ vssd1 vssd1 vccd1 vccd1 _06121_ sky130_fd_sc_hd__o41a_1
XANTENNA__17525__B net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1327 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19793_ clknet_leaf_128_clk _00737_ net1329 vssd1 vssd1 vccd1 vccd1 ag2.body\[607\]
+ sky130_fd_sc_hd__dfrtp_4
X_18744_ clknet_leaf_139_clk img_gen.tracker.next_frame\[182\] net1256 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[182\] sky130_fd_sc_hd__dfrtp_1
X_15956_ ag2.body\[144\] net198 _01657_ ag2.body\[136\] vssd1 vssd1 vccd1 vccd1 _01186_
+ sky130_fd_sc_hd__a22o_1
X_11079_ ag2.body\[542\] net751 net1059 _04199_ _06051_ vssd1 vssd1 vccd1 vccd1 _06052_
+ sky130_fd_sc_hd__a221o_1
XANTENNA__12131__B1 net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12669__B _07539_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1614 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11573__B net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14907_ net2615 net178 _01541_ control.body\[1075\] vssd1 vssd1 vccd1 vccd1 _00253_
+ sky130_fd_sc_hd__a22o_1
X_18675_ clknet_leaf_27_clk img_gen.tracker.next_frame\[113\] net1341 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[113\] sky130_fd_sc_hd__dfrtp_1
X_15887_ ag2.body\[211\] net184 _01649_ ag2.body\[203\] vssd1 vssd1 vccd1 vccd1 _01125_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__17070__B1 net688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17626_ ag2.body\[189\] net949 vssd1 vssd1 vccd1 vccd1 _03305_ sky130_fd_sc_hd__xor2_1
XANTENNA__14959__B1 _01547_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14838_ _08383_ _08388_ _08531_ vssd1 vssd1 vccd1 vccd1 _01509_ sky130_fd_sc_hd__o21a_1
XFILLER_0_53_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12434__A1 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17260__B net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17557_ ag2.body\[356\] net963 vssd1 vssd1 vccd1 vccd1 _03236_ sky130_fd_sc_hd__xor2_1
X_14769_ net1020 ag2.body\[102\] vssd1 vssd1 vccd1 vccd1 _08930_ sky130_fd_sc_hd__or2_1
XFILLER_0_114_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_1489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_43_clk clknet_4_7__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_43_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_89_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16508_ obsg2.obstacleArray\[15\] _02059_ net399 _02186_ vssd1 vssd1 vccd1 vccd1
+ _02187_ sky130_fd_sc_hd__o211a_1
XFILLER_0_74_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19385__CLK clknet_leaf_93_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17488_ ag2.body\[366\] net945 vssd1 vssd1 vccd1 vccd1 _03167_ sky130_fd_sc_hd__xnor2_1
XANTENNA__11642__C1 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_9_clk_A clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19227_ clknet_leaf_75_clk _00171_ net1482 vssd1 vssd1 vccd1 vccd1 ag2.body\[90\]
+ sky130_fd_sc_hd__dfrtp_2
X_16439_ net403 _02117_ net366 vssd1 vssd1 vccd1 vccd1 _02118_ sky130_fd_sc_hd__o21a_1
XANTENNA__16581__C1 net361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15923__A2 net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20362__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09994__A _04573_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19158_ clknet_leaf_50_clk _00102_ net1369 vssd1 vssd1 vccd1 vccd1 ag2.body\[22\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_54_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16604__B net447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19157__RESET_B net1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11588__X _06561_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18109_ obsg2.obstacleArray\[56\] _03688_ net525 vssd1 vssd1 vccd1 vccd1 _01307_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_125_993 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16333__C1 _01912_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19089_ clknet_leaf_9_clk img_gen.tracker.next_frame\[527\] net1271 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[527\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_129_1490 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14405__A net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16884__B1 net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10652__B net1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout304 _07814_ vssd1 vssd1 vccd1 vccd1 net304 sky130_fd_sc_hd__clkbuf_4
Xfanout315 net316 vssd1 vssd1 vccd1 vccd1 net315 sky130_fd_sc_hd__buf_2
X_20002_ clknet_leaf_59_clk _00946_ net1467 vssd1 vssd1 vccd1 vccd1 ag2.body\[384\]
+ sky130_fd_sc_hd__dfrtp_4
Xfanout326 track.nextHighScore\[2\] vssd1 vssd1 vccd1 vccd1 net326 sky130_fd_sc_hd__buf_2
Xfanout337 _07309_ vssd1 vssd1 vccd1 vccd1 net337 sky130_fd_sc_hd__clkbuf_4
X_09813_ net786 control.body\[1048\] control.body\[1052\] net761 _04785_ vssd1 vssd1
+ vccd1 vccd1 _04786_ sky130_fd_sc_hd__a221o_1
Xfanout348 _01731_ vssd1 vssd1 vccd1 vccd1 net348 sky130_fd_sc_hd__clkbuf_4
XANTENNA__17435__B net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout359 net360 vssd1 vssd1 vccd1 vccd1 net359 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_96_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11764__A net1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09744_ ag2.body\[358\] net1088 vssd1 vssd1 vccd1 vccd1 _04717_ sky130_fd_sc_hd__xor2_1
X_09675_ ag2.body\[13\] net1102 vssd1 vssd1 vccd1 vccd1 _04648_ sky130_fd_sc_hd__or2_1
XANTENNA__12673__A1 net289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17061__B1 net935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10684__B1 _04419_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_1460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout720_A net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_7_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12595__A _07431_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout341_X net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout818_A net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_34_clk clknet_4_5__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_34_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout1462_A net1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1083_X net1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout439_X net439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09240__Y _04265_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19927__RESET_B net1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10827__B net1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14178__B2 net988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15375__B1 _01594_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_1518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1250_X net1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout606_X net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19580__RESET_B net1386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10450_ ag2.body\[455\] net1055 vssd1 vssd1 vccd1 vccd1 _05423_ sky130_fd_sc_hd__or2_1
XANTENNA__13925__B2 ag2.body\[61\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11936__B1 net603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09109_ ag2.body\[378\] vssd1 vssd1 vccd1 vccd1 _04134_ sky130_fd_sc_hd__inv_2
XFILLER_0_21_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10381_ ag2.body\[105\] net1212 vssd1 vssd1 vccd1 vccd1 _05354_ sky130_fd_sc_hd__xor2_1
XANTENNA__14315__A net1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19108__CLK clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16875__B1 net690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12120_ _07084_ _07091_ net438 _07078_ vssd1 vssd1 vccd1 vccd1 _07092_ sky130_fd_sc_hd__o211a_1
XFILLER_0_62_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11658__B net1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout975_X net975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12051_ img_gen.tracker.frame\[273\] net593 net555 img_gen.tracker.frame\[270\] _07022_
+ vssd1 vssd1 vccd1 vccd1 _07023_ sky130_fd_sc_hd__a221o_1
XFILLER_0_2_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold380 img_gen.tracker.frame\[263\] vssd1 vssd1 vccd1 vccd1 net1942 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16530__A net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold391 img_gen.tracker.frame\[454\] vssd1 vssd1 vccd1 vccd1 net1953 sky130_fd_sc_hd__dlygate4sd3_1
X_11002_ net779 control.body\[1081\] _05974_ vssd1 vssd1 vccd1 vccd1 _05975_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_79_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19258__CLK clknet_leaf_73_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout860 net861 vssd1 vssd1 vccd1 vccd1 net860 sky130_fd_sc_hd__clkbuf_4
Xfanout871 net872 vssd1 vssd1 vccd1 vccd1 net871 sky130_fd_sc_hd__clkbuf_4
X_15810_ ag2.body\[286\] net207 _01641_ ag2.body\[278\] vssd1 vssd1 vccd1 vccd1 _01056_
+ sky130_fd_sc_hd__a22o_1
Xfanout882 net884 vssd1 vssd1 vccd1 vccd1 net882 sky130_fd_sc_hd__buf_2
X_16790_ obsg2.obstacleArray\[128\] obsg2.obstacleArray\[129\] net457 vssd1 vssd1
+ vccd1 vccd1 _02469_ sky130_fd_sc_hd__mux2_1
XANTENNA__09415__Y _04394_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout893 net894 vssd1 vssd1 vccd1 vccd1 net893 sky130_fd_sc_hd__buf_2
XANTENNA__12113__B1 net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15741_ ag2.body\[336\] net217 _01634_ ag2.body\[328\] vssd1 vssd1 vccd1 vccd1 _00994_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12664__A1 net245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12953_ net685 _07673_ vssd1 vssd1 vccd1 vccd1 _07674_ sky130_fd_sc_hd__nor2_1
Xhold1080 control.body\[804\] vssd1 vssd1 vccd1 vccd1 net2642 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_73_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1091 control.body\[841\] vssd1 vssd1 vccd1 vccd1 net2653 sky130_fd_sc_hd__dlygate4sd3_1
X_11904_ _06875_ _06863_ _06850_ _06691_ vssd1 vssd1 vccd1 vccd1 _06876_ sky130_fd_sc_hd__a2bb2o_1
X_15672_ ag2.body\[403\] net142 _01626_ ag2.body\[395\] vssd1 vssd1 vccd1 vccd1 _00933_
+ sky130_fd_sc_hd__a22o_1
X_18460_ _03847_ _03857_ _03948_ net434 vssd1 vssd1 vccd1 vccd1 _03949_ sky130_fd_sc_hd__a31o_1
XFILLER_0_119_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12884_ net267 _07641_ _07642_ net2046 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[199\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__18176__B net41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14623_ net1036 ag2.body\[468\] vssd1 vssd1 vccd1 vccd1 _08784_ sky130_fd_sc_hd__xor2_1
X_17411_ ag2.body\[284\] net965 vssd1 vssd1 vccd1 vccd1 _03090_ sky130_fd_sc_hd__xor2_1
XFILLER_0_114_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17080__B net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18391_ _08051_ _03794_ _03814_ vssd1 vssd1 vccd1 vccd1 _03881_ sky130_fd_sc_hd__a21bo_1
X_11835_ img_gen.tracker.frame\[566\] net622 net549 img_gen.tracker.frame\[572\] _06806_
+ vssd1 vssd1 vccd1 vccd1 _06807_ sky130_fd_sc_hd__o221a_2
XFILLER_0_115_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_25_clk clknet_4_4__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_25_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_16_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__20385__CLK clknet_leaf_43_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17342_ _03019_ _03020_ vssd1 vssd1 vccd1 vccd1 _03021_ sky130_fd_sc_hd__nand2_1
X_14554_ net973 ag2.body\[67\] vssd1 vssd1 vccd1 vccd1 _08715_ sky130_fd_sc_hd__xnor2_1
XANTENNA__17355__A1 net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11766_ img_gen.tracker.frame\[68\] net542 _06737_ net568 vssd1 vssd1 vccd1 vccd1
+ _06738_ sky130_fd_sc_hd__o211a_1
XFILLER_0_55_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14169__A1 net807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13505_ net328 _07515_ _07813_ vssd1 vssd1 vccd1 vccd1 _07914_ sky130_fd_sc_hd__and3_1
XANTENNA__14169__B2 net791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15366__B1 _01593_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17273_ ag2.body\[558\] net938 vssd1 vssd1 vccd1 vccd1 _02952_ sky130_fd_sc_hd__xor2_1
X_10717_ ag2.body\[617\] net777 net753 ag2.body\[621\] vssd1 vssd1 vccd1 vccd1 _05690_
+ sky130_fd_sc_hd__o22ai_1
X_14485_ net1040 ag2.body\[348\] vssd1 vssd1 vccd1 vccd1 _08646_ sky130_fd_sc_hd__xor2_1
XFILLER_0_86_1629 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11697_ net1070 net1045 vssd1 vssd1 vccd1 vccd1 _06669_ sky130_fd_sc_hd__nor2_1
XFILLER_0_130_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16224_ obsg2.obstacleArray\[36\] net405 vssd1 vssd1 vccd1 vccd1 _01903_ sky130_fd_sc_hd__or2_1
XANTENNA__13916__A1 ag2.body\[61\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19012_ clknet_leaf_1_clk img_gen.tracker.next_frame\[450\] net1247 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[450\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13436_ net682 _07886_ vssd1 vssd1 vccd1 vccd1 _07887_ sky130_fd_sc_hd__nor2_1
X_10648_ ag2.body\[287\] net1066 vssd1 vssd1 vccd1 vccd1 _05621_ sky130_fd_sc_hd__nand2_1
XFILLER_0_70_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19250__RESET_B net1492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16155_ obsg2.obstacleArray\[6\] obsg2.obstacleArray\[7\] net426 vssd1 vssd1 vccd1
+ vccd1 _01834_ sky130_fd_sc_hd__mux2_1
XANTENNA__15118__B1 _01554_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16315__C1 net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13367_ net337 net309 _07532_ vssd1 vssd1 vccd1 vccd1 _07860_ sky130_fd_sc_hd__nor3_1
X_10579_ ag2.body\[187\] net1155 vssd1 vssd1 vccd1 vccd1 _05552_ sky130_fd_sc_hd__xor2_1
XANTENNA__10753__A net1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15106_ net2592 net145 _01564_ control.body\[899\] vssd1 vssd1 vccd1 vccd1 _00429_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_11_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12318_ _07246_ _07251_ vssd1 vssd1 vccd1 vccd1 _07285_ sky130_fd_sc_hd__or2_1
X_16086_ obsg2.obstacleArray\[114\] obsg2.obstacleArray\[115\] net423 vssd1 vssd1
+ vccd1 vccd1 _01765_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20155__RESET_B net1442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13298_ _07480_ net302 vssd1 vssd1 vccd1 vccd1 _07833_ sky130_fd_sc_hd__nor2_1
XFILLER_0_107_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19914_ clknet_leaf_55_clk _00858_ net1456 vssd1 vssd1 vccd1 vccd1 ag2.body\[472\]
+ sky130_fd_sc_hd__dfrtp_4
X_15037_ control.body\[973\] net165 _01557_ net2408 vssd1 vssd1 vccd1 vccd1 _00367_
+ sky130_fd_sc_hd__a22o_1
X_12249_ _07196_ _07209_ _07215_ vssd1 vssd1 vccd1 vccd1 _07219_ sky130_fd_sc_hd__and3_1
XANTENNA__09899__A2 net1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19845_ clknet_leaf_92_clk _00789_ net1414 vssd1 vssd1 vccd1 vccd1 ag2.body\[547\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_23_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17255__B net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11584__A net1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19776_ clknet_leaf_19_clk _00720_ net1331 vssd1 vssd1 vccd1 vccd1 ag2.body\[622\]
+ sky130_fd_sc_hd__dfrtp_4
X_16988_ ag2.body\[91\] net853 vssd1 vssd1 vccd1 vccd1 _02667_ sky130_fd_sc_hd__nand2_1
XANTENNA__18625__CLK clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12104__B1 net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18727_ clknet_leaf_144_clk img_gen.tracker.next_frame\[165\] net1253 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[165\] sky130_fd_sc_hd__dfrtp_1
X_15939_ ag2.body\[161\] net195 _01653_ ag2.body\[153\] vssd1 vssd1 vccd1 vccd1 _01171_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_95_1482 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09460_ net894 net899 net907 net903 vssd1 vssd1 vccd1 vccd1 _04433_ sky130_fd_sc_hd__or4b_4
XFILLER_0_17_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18658_ clknet_leaf_14_clk img_gen.tracker.next_frame\[96\] net1276 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[96\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_133_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_1379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17609_ net956 net930 vssd1 vssd1 vccd1 vccd1 _03288_ sky130_fd_sc_hd__nor2_1
XFILLER_0_56_1499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09391_ _04354_ _04379_ vssd1 vssd1 vccd1 vccd1 _01407_ sky130_fd_sc_hd__nor2_1
XANTENNA__18775__CLK clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18589_ clknet_leaf_13_clk img_gen.tracker.next_frame\[27\] net1284 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[27\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_1010 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_16_clk clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_16_clk
+ sky130_fd_sc_hd__clkbuf_8
X_20620_ net1545 vssd1 vssd1 vccd1 vccd1 gpio_oeb[32] sky130_fd_sc_hd__buf_2
XANTENNA__11615__C1 net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13304__A net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09501__B net1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13080__A1 net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_573 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10647__B net1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13023__B net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20551_ clknet_leaf_105_clk _01416_ _00025_ vssd1 vssd1 vccd1 vccd1 sound_gen.osc1.stayCount\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__15357__B1 _01592_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09995__Y _04968_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1106 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout134_A net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20482_ clknet_leaf_39_clk _01369_ net1356 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[118\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_85_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11918__B1 net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16334__B net411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14580__B2 net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10663__A net1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14135__A net972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10382__B net1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14332__A1 net835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_3663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_682 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19400__CLK clknet_leaf_102_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14332__B2 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_3674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_3685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1210_A net1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout101 net104 vssd1 vssd1 vccd1 vccd1 net101 sky130_fd_sc_hd__buf_2
Xfanout112 net113 vssd1 vssd1 vccd1 vccd1 net112 sky130_fd_sc_hd__clkbuf_2
Xfanout123 net124 vssd1 vssd1 vccd1 vccd1 net123 sky130_fd_sc_hd__buf_2
XANTENNA__20258__CLK clknet_leaf_43_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout134 net135 vssd1 vssd1 vccd1 vccd1 net134 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout145 net146 vssd1 vssd1 vccd1 vccd1 net145 sky130_fd_sc_hd__buf_2
XANTENNA_fanout670_A net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout156 net162 vssd1 vssd1 vccd1 vccd1 net156 sky130_fd_sc_hd__clkbuf_2
Xfanout167 net169 vssd1 vssd1 vccd1 vccd1 net167 sky130_fd_sc_hd__buf_2
XANTENNA_fanout768_A _04230_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17733__X _03412_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout178 net180 vssd1 vssd1 vccd1 vccd1 net178 sky130_fd_sc_hd__buf_2
Xfanout189 net191 vssd1 vssd1 vccd1 vccd1 net189 sky130_fd_sc_hd__buf_2
XANTENNA__19550__CLK clknet_leaf_115_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_114_Right_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_1279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09727_ ag2.body\[91\] net772 net757 ag2.body\[93\] _04699_ vssd1 vssd1 vccd1 vccd1
+ _04700_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout935_A net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout556_X net556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12102__B net1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09658_ _04625_ _04627_ _04629_ _04630_ _04618_ vssd1 vssd1 vccd1 vccd1 _04631_ sky130_fd_sc_hd__o41a_1
XANTENNA__17585__A1 ag2.body\[56\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_3489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_2_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout47_A net48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17585__B2 ag2.body\[62\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14399__A1 net821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14399__B2 net1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout723_X net723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16793__C1 net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09589_ net1202 control.body\[905\] vssd1 vssd1 vccd1 vccd1 _04562_ sky130_fd_sc_hd__xor2_1
XANTENNA_fanout1465_X net1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11620_ obsg2.obstacleArray\[49\] net511 net504 _06592_ vssd1 vssd1 vccd1 vccd1 _06593_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_72_1290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13214__A net675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10557__B net1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_1420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_1431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11551_ net1222 net1195 vssd1 vssd1 vccd1 vccd1 _06524_ sky130_fd_sc_hd__nand2_1
XANTENNA__11621__A2 net631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17888__A2 _03519_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16525__A net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10502_ net1205 control.body\[977\] vssd1 vssd1 vccd1 vccd1 _05475_ sky130_fd_sc_hd__xor2_1
X_14270_ net972 _03977_ _03978_ net1036 _08430_ vssd1 vssd1 vccd1 vccd1 _08431_ sky130_fd_sc_hd__a221o_1
Xwire535 _04291_ vssd1 vssd1 vccd1 vccd1 net535 sky130_fd_sc_hd__buf_1
X_11482_ _06433_ _06440_ _06441_ _06454_ vssd1 vssd1 vccd1 vccd1 _06455_ sky130_fd_sc_hd__o22a_1
XANTENNA__11909__B1 net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13221_ net241 _07799_ _07800_ net2019 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[378\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__09578__A1 net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10433_ net1180 control.body\[930\] vssd1 vssd1 vccd1 vccd1 _05406_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_122_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16812__X _02491_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14045__A net1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10188__A2 net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13152_ net667 _07767_ vssd1 vssd1 vccd1 vccd1 _07768_ sky130_fd_sc_hd__nor2_1
X_10364_ net758 control.body\[764\] control.body\[765\] net753 vssd1 vssd1 vccd1 vccd1
+ _05337_ sky130_fd_sc_hd__a22o_1
XFILLER_0_108_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12103_ img_gen.tracker.frame\[363\] net610 net555 img_gen.tracker.frame\[366\] _07074_
+ vssd1 vssd1 vccd1 vccd1 _07075_ sky130_fd_sc_hd__a221o_1
X_17960_ net539 net537 net462 net957 vssd1 vssd1 vccd1 vccd1 _03585_ sky130_fd_sc_hd__and4b_1
XANTENNA__14323__B2 net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13083_ net685 _07734_ vssd1 vssd1 vccd1 vccd1 _07735_ sky130_fd_sc_hd__nor2_1
XANTENNA_clkbuf_leaf_127_clk_X clknet_leaf_127_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10295_ ag2.body\[333\] net1116 vssd1 vssd1 vccd1 vccd1 _05268_ sky130_fd_sc_hd__xor2_1
XANTENNA__12334__B1 _06825_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14874__A2 net182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11675__Y _06647_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12034_ img_gen.tracker.frame\[39\] net612 net557 img_gen.tracker.frame\[42\] _07005_
+ vssd1 vssd1 vccd1 vccd1 _07006_ sky130_fd_sc_hd__a221o_1
X_16911_ _04206_ net869 net710 ag2.body\[564\] vssd1 vssd1 vccd1 vccd1 _02590_ sky130_fd_sc_hd__a22o_1
XANTENNA__17075__B net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17891_ net530 _03530_ vssd1 vssd1 vccd1 vccd1 _03531_ sky130_fd_sc_hd__and2_2
XFILLER_0_40_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12885__A1 net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16076__A1 net375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1571 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19630_ clknet_leaf_123_clk _00574_ net1406 vssd1 vssd1 vccd1 vccd1 control.body\[764\]
+ sky130_fd_sc_hd__dfrtp_1
X_16842_ ag2.body\[169\] net871 vssd1 vssd1 vccd1 vccd1 _02521_ sky130_fd_sc_hd__or2_1
XANTENNA__10360__A2 net752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout690 net691 vssd1 vssd1 vccd1 vccd1 net690 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_137_1011 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19561_ clknet_leaf_115_clk _00505_ net1397 vssd1 vssd1 vccd1 vccd1 control.body\[839\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12637__A1 net264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13985_ ag2.body\[122\] net211 _08159_ ag2.body\[114\] vssd1 vssd1 vccd1 vccd1 _00203_
+ sky130_fd_sc_hd__a22o_1
X_16773_ _02449_ _02451_ net499 vssd1 vssd1 vccd1 vccd1 _02452_ sky130_fd_sc_hd__mux2_1
XANTENNA__18798__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18512_ net1513 net1507 vssd1 vssd1 vccd1 vccd1 _00043_ sky130_fd_sc_hd__or2_1
X_15724_ ag2.body\[353\] net194 _01632_ ag2.body\[345\] vssd1 vssd1 vccd1 vccd1 _00979_
+ sky130_fd_sc_hd__a22o_1
X_12936_ net679 _07665_ vssd1 vssd1 vccd1 vccd1 _07666_ sky130_fd_sc_hd__nor2_1
X_19492_ clknet_leaf_114_clk _00436_ net1399 vssd1 vssd1 vccd1 vccd1 control.body\[898\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_92_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1174 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_4_8__f_clk_A clknet_3_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09602__A net1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18443_ _03929_ _03930_ _03931_ _03851_ vssd1 vssd1 vccd1 vccd1 _03932_ sky130_fd_sc_hd__o22a_1
X_15655_ ag2.body\[420\] net138 _01624_ ag2.body\[412\] vssd1 vssd1 vccd1 vccd1 _00918_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_115_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12867_ net239 _07634_ _07635_ net1659 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[189\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_115_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16784__C1 net352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11860__A2 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14606_ net994 ag2.body\[129\] vssd1 vssd1 vccd1 vccd1 _08767_ sky130_fd_sc_hd__xor2_1
XFILLER_0_28_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11818_ img_gen.tracker.frame\[404\] net545 _06789_ net571 vssd1 vssd1 vccd1 vccd1
+ _06790_ sky130_fd_sc_hd__o211a_1
X_15586_ ag2.body\[486\] net130 _01617_ ag2.body\[478\] vssd1 vssd1 vccd1 vccd1 _00856_
+ sky130_fd_sc_hd__a22o_1
X_18374_ _07181_ track.nextHighScore\[0\] _03865_ vssd1 vssd1 vccd1 vccd1 _01395_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_56_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12798_ net232 _07601_ _07602_ net2090 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[153\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11073__B1 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17325_ _02996_ _02998_ _02999_ _03003_ vssd1 vssd1 vccd1 vccd1 _03004_ sky130_fd_sc_hd__or4_1
XANTENNA__15339__B1 _01590_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14537_ _08695_ _08697_ vssd1 vssd1 vccd1 vccd1 _08698_ sky130_fd_sc_hd__nor2_1
X_11749_ net748 _06630_ vssd1 vssd1 vccd1 vccd1 _06721_ sky130_fd_sc_hd__nand2_1
XANTENNA__12963__A net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_133_4375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14468_ net1020 ag2.body\[270\] vssd1 vssd1 vccd1 vccd1 _08629_ sky130_fd_sc_hd__or2_1
X_17256_ ag2.body\[551\] net688 net723 ag2.body\[546\] vssd1 vssd1 vccd1 vccd1 _02935_
+ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_133_4386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12682__B _07546_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_1592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16207_ _01724_ _01837_ _01854_ _01885_ vssd1 vssd1 vccd1 vccd1 _01886_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_12_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13419_ net282 _07878_ _07879_ net1783 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[497\]
+ sky130_fd_sc_hd__a22o_1
X_17187_ ag2.body\[574\] net938 vssd1 vssd1 vccd1 vccd1 _02866_ sky130_fd_sc_hd__xor2_1
X_14399_ net821 ag2.body\[123\] _04032_ net1014 _08554_ vssd1 vssd1 vccd1 vccd1 _08560_
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_113_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10179__A2 net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16839__B1 net699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16138_ _01698_ _01816_ vssd1 vssd1 vccd1 vccd1 _01817_ sky130_fd_sc_hd__xor2_2
XFILLER_0_110_911 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14314__A1 net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16069_ obsg2.obstacleArray\[122\] obsg2.obstacleArray\[123\] net424 vssd1 vssd1
+ vccd1 vccd1 _01748_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08960_ ag2.body\[31\] vssd1 vssd1 vccd1 vccd1 _03985_ sky130_fd_sc_hd__inv_2
XANTENNA__14314__B2 net980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_5_clk clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_5_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_55_1986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_1997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17264__B1 net873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19828_ clknet_leaf_124_clk _00772_ net1407 vssd1 vssd1 vccd1 vccd1 ag2.body\[562\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__17803__A2 net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14617__A2 ag2.body\[59\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20550__CLK clknet_leaf_105_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19759_ clknet_leaf_130_clk net2488 net1316 vssd1 vssd1 vccd1 vccd1 control.body\[637\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_91_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09512_ net1100 control.body\[837\] vssd1 vssd1 vccd1 vccd1 _04485_ sky130_fd_sc_hd__nand2_1
XFILLER_0_91_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1105 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09512__A net1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09443_ net891 net898 vssd1 vssd1 vccd1 vccd1 _04416_ sky130_fd_sc_hd__nor2_4
XANTENNA_fanout251_A net260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09374_ sound_gen.osc1.stayCount\[17\] _04360_ net270 vssd1 vssd1 vccd1 vccd1 _04372_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_93_249 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10377__B net1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20603_ net1535 vssd1 vssd1 vccd1 vccd1 gpio_oeb[15] sky130_fd_sc_hd__buf_2
XFILLER_0_62_603 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11603__A2 net632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12800__A1 net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1160_A net1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20534_ clknet_leaf_107_clk _01399_ _00008_ vssd1 vssd1 vccd1 vccd1 sound_gen.osc1.stayCount\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_116_3850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_116_3861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11489__A net1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_116_3872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12013__C1 _06724_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_3725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20465_ clknet_leaf_32_clk _01352_ net1345 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[101\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__10393__A net1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout304_X net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_3736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_81_clk_A clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_3747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1046_X net1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20396_ clknet_leaf_30_clk _01283_ net1336 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[32\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA_fanout885_A net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1213_X net1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10080_ net1226 control.body\[792\] vssd1 vssd1 vccd1 vccd1 _05053_ sky130_fd_sc_hd__nand2_1
XANTENNA__12867__A1 net239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_96_clk_A clknet_4_11__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout673_X net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13209__A net676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17904__A net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10342__A2 net780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1331 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout840_X net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17623__B net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout938_X net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13770_ img_gen.updater.commands.count\[7\] _08081_ _08083_ _08071_ vssd1 vssd1 vccd1
+ vccd1 _00064_ sky130_fd_sc_hd__o211a_1
XANTENNA__09496__B1 _04430_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12095__A2 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10982_ net1101 control.body\[757\] vssd1 vssd1 vccd1 vccd1 _05955_ sky130_fd_sc_hd__xor2_1
XANTENNA__13292__A1 net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12767__B _07483_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_84_2872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12721_ net305 _07564_ vssd1 vssd1 vccd1 vccd1 _07565_ sky130_fd_sc_hd__nor2_1
XFILLER_0_116_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_84_2883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11842__A2 net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_2894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15440_ ag2.body\[613\] net82 _01600_ ag2.body\[605\] vssd1 vssd1 vccd1 vccd1 _00727_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_65_2293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_1526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_2758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12652_ net264 _07529_ _07530_ net1693 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[79\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_34_clk_A clknet_4_5__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_2769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11603_ obsg2.obstacleArray\[23\] net632 net514 obsg2.obstacleArray\[19\] net508
+ vssd1 vssd1 vccd1 vccd1 _06576_ sky130_fd_sc_hd__o221a_1
XANTENNA__11055__B1 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15371_ net2606 net68 _01593_ net2292 vssd1 vssd1 vccd1 vccd1 _00665_ sky130_fd_sc_hd__a22o_1
XANTENNA__14792__A1 net974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_2179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16518__C1 _02075_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12583_ net230 _07491_ _07492_ net2064 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[48\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__14792__B2 net1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14322_ net807 ag2.body\[453\] ag2.body\[451\] net818 vssd1 vssd1 vccd1 vccd1 _08483_
+ sky130_fd_sc_hd__a2bb2o_1
X_17110_ _02780_ _02781_ _02787_ _02788_ vssd1 vssd1 vccd1 vccd1 _02789_ sky130_fd_sc_hd__a211o_1
X_18090_ net44 _03675_ vssd1 vssd1 vccd1 vccd1 _03676_ sky130_fd_sc_hd__nor2_1
X_11534_ net777 net1174 net1152 _06491_ vssd1 vssd1 vccd1 vccd1 _06507_ sky130_fd_sc_hd__a31o_1
XFILLER_0_92_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17730__A1 net496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17785__S net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20423__CLK clknet_leaf_37_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17041_ ag2.body\[120\] net740 net944 _04031_ _02719_ vssd1 vssd1 vccd1 vccd1 _02720_
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_81_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_22_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_850 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14253_ net822 ag2.body\[75\] ag2.body\[79\] net797 vssd1 vssd1 vccd1 vccd1 _08414_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_52_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14544__A1 net1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11465_ ag2.body\[257\] net1210 vssd1 vssd1 vccd1 vccd1 _06438_ sky130_fd_sc_hd__xnor2_1
XANTENNA__14544__B2 net1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_2687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_2698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_1312 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13204_ net242 _07791_ _07792_ net1611 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[369\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__19596__CLK clknet_leaf_118_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10416_ _05023_ _05146_ _05272_ _05388_ vssd1 vssd1 vccd1 vccd1 _05389_ sky130_fd_sc_hd__nand4_1
X_14184_ net819 ag2.body\[195\] _08335_ _08336_ _08344_ vssd1 vssd1 vccd1 vccd1 _08345_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_0_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11396_ _04573_ _06358_ _06363_ _06368_ vssd1 vssd1 vccd1 vccd1 _06369_ sky130_fd_sc_hd__or4_2
XFILLER_0_81_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17494__B1 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13135_ net243 _07758_ _07759_ net1784 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[333\]
+ sky130_fd_sc_hd__a22o_1
X_10347_ ag2.body\[289\] net1210 vssd1 vssd1 vccd1 vccd1 _05320_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18992_ clknet_leaf_8_clk img_gen.tracker.next_frame\[430\] net1272 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[430\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__14503__A net1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17943_ net517 _03572_ vssd1 vssd1 vccd1 vccd1 _01257_ sky130_fd_sc_hd__nor2_1
X_13066_ net685 _07726_ vssd1 vssd1 vccd1 vccd1 _07727_ sky130_fd_sc_hd__nor2_1
X_10278_ _05242_ _05243_ _05244_ _05245_ vssd1 vssd1 vccd1 vccd1 _05251_ sky130_fd_sc_hd__or4_1
XFILLER_0_40_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1430 net1435 vssd1 vssd1 vccd1 vccd1 net1430 sky130_fd_sc_hd__buf_2
XANTENNA__17246__B1 net858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12017_ img_gen.tracker.frame\[231\] net612 net594 img_gen.tracker.frame\[237\] _06988_
+ vssd1 vssd1 vccd1 vccd1 _06989_ sky130_fd_sc_hd__a221o_1
XANTENNA_clkbuf_leaf_107_clk_A clknet_4_10__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1441 net1442 vssd1 vssd1 vccd1 vccd1 net1441 sky130_fd_sc_hd__buf_2
X_17874_ _03506_ _03516_ vssd1 vssd1 vccd1 vccd1 _01244_ sky130_fd_sc_hd__nor2_1
XFILLER_0_20_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout1452 net1453 vssd1 vssd1 vccd1 vccd1 net1452 sky130_fd_sc_hd__clkbuf_2
Xfanout1463 net1464 vssd1 vssd1 vccd1 vccd1 net1463 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_79_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout1474 net1475 vssd1 vssd1 vccd1 vccd1 net1474 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_122_4032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19613_ clknet_leaf_120_clk _00557_ net1395 vssd1 vssd1 vccd1 vccd1 control.body\[779\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_50_1850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_122_4043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_50_1861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16825_ ag2.body\[227\] net854 vssd1 vssd1 vccd1 vccd1 _02504_ sky130_fd_sc_hd__xor2_1
Xfanout1485 net1493 vssd1 vssd1 vccd1 vccd1 net1485 sky130_fd_sc_hd__clkbuf_4
Xfanout1496 net1499 vssd1 vssd1 vccd1 vccd1 net1496 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_122_4054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12958__A _07490_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19544_ clknet_leaf_118_clk _00488_ net1389 vssd1 vssd1 vccd1 vccd1 control.body\[854\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_31_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11818__C1 net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16756_ _02427_ _02430_ _02432_ _02434_ net499 net380 vssd1 vssd1 vccd1 vccd1 _02435_
+ sky130_fd_sc_hd__mux4_1
X_13968_ ag2.body\[107\] net202 _08157_ ag2.body\[99\] vssd1 vssd1 vccd1 vccd1 _00188_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__16149__B net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15707_ ag2.body\[371\] net141 _01629_ ag2.body\[363\] vssd1 vssd1 vccd1 vccd1 _00965_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_48_408 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_wire317_A _06459_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11294__B1 _06253_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19475_ clknet_leaf_110_clk net2094 net1416 vssd1 vssd1 vccd1 vccd1 control.body\[913\]
+ sky130_fd_sc_hd__dfrtp_1
X_12919_ net243 _07656_ _07657_ net1694 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[219\]
+ sky130_fd_sc_hd__a22o_1
X_16687_ net395 _02290_ _02291_ _02292_ net361 vssd1 vssd1 vccd1 vccd1 _02366_ sky130_fd_sc_hd__a221o_1
XANTENNA__11833__A2 net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13899_ ag2.body\[46\] net85 _08149_ ag2.body\[38\] vssd1 vssd1 vccd1 vccd1 _00127_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_18_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18426_ _03782_ _03787_ vssd1 vssd1 vccd1 vccd1 _03915_ sky130_fd_sc_hd__nand2b_1
X_15638_ ag2.body\[437\] net125 _01622_ ag2.body\[429\] vssd1 vssd1 vccd1 vccd1 _00903_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_118_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13035__A1 net262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_135_4426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_135_4437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16772__A2 net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_135_4448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18357_ net321 _03787_ _03792_ _03796_ _03784_ vssd1 vssd1 vccd1 vccd1 _03852_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_5_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14783__A1 net975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15569_ _06441_ net61 vssd1 vssd1 vccd1 vccd1 _01615_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_44_1665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14783__B2 net1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11597__A1 net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17308_ ag2.body\[397\] net949 vssd1 vssd1 vccd1 vccd1 _02987_ sky130_fd_sc_hd__or2_1
XFILLER_0_72_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_20_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09090_ ag2.body\[330\] vssd1 vssd1 vccd1 vccd1 _04115_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_20_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18288_ net324 net321 vssd1 vssd1 vccd1 vccd1 _03784_ sky130_fd_sc_hd__or2_1
XFILLER_0_4_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14535__A1 net1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17239_ _04222_ net879 net704 ag2.body\[621\] vssd1 vssd1 vccd1 vccd1 _02918_ sky130_fd_sc_hd__a22o_1
XANTENNA__14535__B2 net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_94_3190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold902 control.body\[725\] vssd1 vssd1 vccd1 vccd1 net2464 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_128_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold913 control.body\[953\] vssd1 vssd1 vccd1 vccd1 net2475 sky130_fd_sc_hd__dlygate4sd3_1
X_20250_ clknet_leaf_68_clk _01194_ net1498 vssd1 vssd1 vccd1 vccd1 ag2.body\[136\]
+ sky130_fd_sc_hd__dfrtp_4
Xhold924 _00244_ vssd1 vssd1 vccd1 vccd1 net2486 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_3054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold935 control.body\[816\] vssd1 vssd1 vccd1 vccd1 net2497 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__16612__B net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_3065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold946 _00546_ vssd1 vssd1 vccd1 vccd1 net2508 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_3076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold957 control.body\[953\] vssd1 vssd1 vccd1 vccd1 net2519 sky130_fd_sc_hd__dlygate4sd3_1
X_20181_ clknet_leaf_87_clk _01125_ net1460 vssd1 vssd1 vccd1 vccd1 ag2.body\[211\]
+ sky130_fd_sc_hd__dfrtp_4
Xhold968 _00465_ vssd1 vssd1 vccd1 vccd1 net2530 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__16104__S net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09992_ net743 control.body\[735\] control.body\[732\] net758 vssd1 vssd1 vccd1 vccd1
+ _04965_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_110_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold979 _00303_ vssd1 vssd1 vccd1 vccd1 net2541 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_86_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_38_1469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_122_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08943_ net977 vssd1 vssd1 vccd1 vccd1 _03968_ sky130_fd_sc_hd__inv_2
XANTENNA__12849__A1 net239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10005__X _04978_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17788__A1 net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_4_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18098__Y _03681_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1006_A net1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_4_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_4_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_105_3540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout466_A _06660_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1537 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_3404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12077__A2 net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_3415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10088__A1 net1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09242__A net947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1009 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10088__B2 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10388__A net1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11824__A2 net584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout254_X net254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16212__A1 net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1375_A net1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09426_ _04402_ vssd1 vssd1 vccd1 vccd1 track.current_collision sky130_fd_sc_hd__inv_2
XFILLER_0_36_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16763__A2 net493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_118_3912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_118_3923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09357_ _04358_ vssd1 vssd1 vccd1 vccd1 _04359_ sky130_fd_sc_hd__inv_2
XFILLER_0_47_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_118_3934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout421_X net421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout800_A net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09896__B net1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1163_X net1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout519_X net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_114_3809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09288_ net2489 _04285_ _04284_ vssd1 vssd1 vccd1 vccd1 _04309_ sky130_fd_sc_hd__o21bai_2
XANTENNA__17712__A1 net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10835__B net1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_1476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20517_ clknet_leaf_114_clk track.nextHighScore\[7\] net1398 vssd1 vssd1 vccd1 vccd1
+ track.highScore\[7\] sky130_fd_sc_hd__dfrtp_2
XANTENNA__18290__A track.nextHighScore\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_1617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11250_ _06209_ _06210_ _06219_ _06220_ vssd1 vssd1 vccd1 vccd1 _06223_ sky130_fd_sc_hd__a22o_1
X_20448_ clknet_leaf_41_clk _01335_ net1371 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[84\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_15_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout790_X net790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout888_X net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10201_ ag2.body\[112\] net1235 vssd1 vssd1 vccd1 vccd1 _05174_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_73_2540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09953__A1 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11181_ ag2.body\[180\] net1127 vssd1 vssd1 vccd1 vccd1 _06154_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_73_2562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1015 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12552__A3 _07444_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20379_ clknet_leaf_25_clk _01266_ net1343 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[15\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_43_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14829__A2 _08654_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10132_ net1049 control.body\[823\] vssd1 vssd1 vccd1 vccd1 _05105_ sky130_fd_sc_hd__or2_1
XFILLER_0_101_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10570__B _04519_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17634__A ag2.body\[164\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14940_ net2406 net173 _01545_ control.body\[1040\] vssd1 vssd1 vccd1 vccd1 _00282_
+ sky130_fd_sc_hd__a22o_1
X_10063_ _04445_ _04519_ _04600_ _04521_ vssd1 vssd1 vccd1 vccd1 _05036_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_86_2934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14871_ net2169 net182 _01537_ control.body\[1107\] vssd1 vssd1 vccd1 vccd1 _00221_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_86_2945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16610_ _02287_ _02288_ net391 vssd1 vssd1 vccd1 vccd1 _02289_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_86_2956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13822_ control.body_update.direction\[0\] _08118_ vssd1 vssd1 vccd1 vccd1 _08119_
+ sky130_fd_sc_hd__nor2_2
XFILLER_0_54_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09469__B1 net1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_2809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17590_ ag2.body\[59\] net716 net947 _03997_ _03268_ vssd1 vssd1 vccd1 vccd1 _03269_
+ sky130_fd_sc_hd__a221o_1
XANTENNA__13265__A1 net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_2355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_2366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10079__A1 _04420_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_2377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16541_ net497 _02219_ vssd1 vssd1 vccd1 vccd1 _02220_ sky130_fd_sc_hd__nand2_4
X_13753_ _08060_ _08069_ _08071_ _08067_ vssd1 vssd1 vccd1 vccd1 _00059_ sky130_fd_sc_hd__o211a_1
XFILLER_0_39_1291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10965_ net1059 control.body\[1007\] vssd1 vssd1 vccd1 vccd1 _05938_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_85_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1521 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12704_ net1968 net647 _07556_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[105\]
+ sky130_fd_sc_hd__and3_1
XFILLER_0_70_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19260_ clknet_leaf_73_clk _00204_ net1500 vssd1 vssd1 vccd1 vccd1 ag2.body\[123\]
+ sky130_fd_sc_hd__dfrtp_4
X_16472_ net364 _02149_ _02075_ vssd1 vssd1 vccd1 vccd1 _02151_ sky130_fd_sc_hd__a21o_1
XANTENNA__18836__CLK clknet_leaf_141_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13684_ _04944_ _05697_ vssd1 vssd1 vccd1 vccd1 _08028_ sky130_fd_sc_hd__nand2_2
X_10896_ _05858_ _05860_ _05868_ _05857_ vssd1 vssd1 vccd1 vccd1 _05869_ sky130_fd_sc_hd__or4b_2
XFILLER_0_39_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18184__B net41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16754__A2 net500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18211_ obsg2.obstacleArray\[102\] _03744_ net521 vssd1 vssd1 vccd1 vccd1 _01353_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_128_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12635_ net676 _07520_ vssd1 vssd1 vccd1 vccd1 _07521_ sky130_fd_sc_hd__nor2_1
X_15423_ control.body\[630\] net81 _01598_ ag2.body\[622\] vssd1 vssd1 vccd1 vccd1
+ _00712_ sky130_fd_sc_hd__a22o_1
XFILLER_0_66_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19191_ clknet_leaf_126_clk _00135_ net1332 vssd1 vssd1 vccd1 vccd1 ag2.body\[54\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_14_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_1464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18142_ _03563_ net37 obsg2.obstacleArray\[68\] vssd1 vssd1 vccd1 vccd1 _03710_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_25_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15354_ _05870_ net53 vssd1 vssd1 vccd1 vccd1 _01592_ sky130_fd_sc_hd__nor2_4
XTAP_TAPCELL_ROW_130_4301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12566_ net292 _07481_ _07482_ net2010 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[41\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__10745__B net1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14305_ _08458_ _08461_ _08462_ _08465_ vssd1 vssd1 vccd1 vccd1 _08466_ sky130_fd_sc_hd__or4b_1
XFILLER_0_41_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18986__CLK clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11517_ net1195 net1174 vssd1 vssd1 vccd1 vccd1 _06490_ sky130_fd_sc_hd__nor2_2
XANTENNA__13121__B _07584_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18073_ net42 _03664_ vssd1 vssd1 vccd1 vccd1 _03665_ sky130_fd_sc_hd__nor2_1
X_15285_ control.body\[746\] net78 _01584_ net2342 vssd1 vssd1 vccd1 vccd1 _00588_
+ sky130_fd_sc_hd__a22o_1
X_12497_ net388 _07442_ vssd1 vssd1 vccd1 vccd1 _07443_ sky130_fd_sc_hd__or2_2
XANTENNA__12018__A net1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17024_ _02697_ _02699_ _02702_ vssd1 vssd1 vccd1 vccd1 _02703_ sky130_fd_sc_hd__or3_2
X_14236_ _08394_ _08395_ _08396_ _08393_ vssd1 vssd1 vccd1 vccd1 _08397_ sky130_fd_sc_hd__a211o_1
XFILLER_0_80_296 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold209 img_gen.tracker.frame\[187\] vssd1 vssd1 vccd1 vccd1 net1771 sky130_fd_sc_hd__dlygate4sd3_1
X_11448_ net1181 control.body\[954\] vssd1 vssd1 vccd1 vccd1 _06421_ sky130_fd_sc_hd__xor2_1
XFILLER_0_1_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17528__B net951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16432__B net453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14167_ net831 ag2.body\[202\] ag2.body\[206\] net799 _08325_ vssd1 vssd1 vccd1 vccd1
+ _08328_ sky130_fd_sc_hd__a221o_1
X_11379_ _04169_ net1155 net1104 _04170_ vssd1 vssd1 vccd1 vccd1 _06352_ sky130_fd_sc_hd__o22a_1
XANTENNA__14233__A net1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_128_4230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_4241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11751__A1 net466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13118_ net243 _07750_ _07751_ net1978 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[324\]
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_52_1901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15048__B net59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18975_ clknet_leaf_8_clk img_gen.tracker.next_frame\[413\] net1270 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[413\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_52_1912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14098_ net1015 ag2.body\[590\] vssd1 vssd1 vccd1 vccd1 _08259_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_124_4105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_4116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17219__B1 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16690__B2 _02368_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17926_ net48 _03552_ _03558_ vssd1 vssd1 vccd1 vccd1 _03559_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_33_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13049_ net680 _07718_ vssd1 vssd1 vccd1 vccd1 _07719_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_0_Left_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_33_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1260 net1263 vssd1 vssd1 vccd1 vccd1 net1260 sky130_fd_sc_hd__clkbuf_2
Xfanout1271 net1272 vssd1 vssd1 vccd1 vccd1 net1271 sky130_fd_sc_hd__clkbuf_4
X_17857_ _07317_ img_gen.updater.commands.rR1.rainbowRNG\[0\] img_gen.updater.commands.rR1.rainbowRNG\[1\]
+ img_gen.updater.commands.rR1.rainbowRNG\[2\] vssd1 vssd1 vccd1 vccd1 _03511_ sky130_fd_sc_hd__and4b_1
Xfanout1282 net1286 vssd1 vssd1 vccd1 vccd1 net1282 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12688__A net673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1293 net1311 vssd1 vssd1 vccd1 vccd1 net1293 sky130_fd_sc_hd__buf_2
X_16808_ _03999_ net877 net693 ag2.body\[71\] vssd1 vssd1 vccd1 vccd1 _02487_ sky130_fd_sc_hd__o22a_1
XANTENNA__12059__A2 net627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13256__A1 net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17788_ net1036 _03460_ net1027 vssd1 vssd1 vccd1 vccd1 _03465_ sky130_fd_sc_hd__a21o_1
Xclkbuf_3_4_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_3_4_0_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__16993__A2 net876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19527_ clknet_leaf_120_clk _00471_ net1393 vssd1 vssd1 vccd1 vccd1 control.body\[869\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__15999__A net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16739_ obsg2.obstacleArray\[48\] net491 net487 obsg2.obstacleArray\[50\] _02417_
+ vssd1 vssd1 vccd1 vccd1 _02418_ sky130_fd_sc_hd__a221o_1
XFILLER_0_88_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16594__S net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18375__A track.nextHighScore\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_46_1727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09997__A net1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19458_ clknet_leaf_110_clk _00402_ net1418 vssd1 vssd1 vccd1 vccd1 control.body\[928\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10001__A net1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_27_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17942__A1 net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09211_ net896 vssd1 vssd1 vccd1 vccd1 _04236_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_27_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18409_ _04639_ _08140_ _03824_ _03898_ vssd1 vssd1 vccd1 vccd1 _03899_ sky130_fd_sc_hd__a22o_1
XFILLER_0_17_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19389_ clknet_leaf_112_clk _00333_ net1425 vssd1 vssd1 vccd1 vccd1 control.body\[1003\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_91_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_96_3241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09142_ ag2.body\[471\] vssd1 vssd1 vccd1 vccd1 _04167_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_96_3252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_96_3263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10655__B net1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_92_3116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15705__B1 _01629_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_3127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09073_ ag2.body\[299\] vssd1 vssd1 vccd1 vccd1 _04098_ sky130_fd_sc_hd__inv_2
XANTENNA__12573__D net559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13031__B _07539_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_1330 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_3138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout214_A net218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20302_ clknet_leaf_37_clk net6 net1349 vssd1 vssd1 vccd1 vccd1 control.divider.synch.Q\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold710 control.body\[686\] vssd1 vssd1 vccd1 vccd1 net2272 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_128_1385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold721 control.body\[691\] vssd1 vssd1 vccd1 vccd1 net2283 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold732 _00259_ vssd1 vssd1 vccd1 vccd1 net2294 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__17458__B1 net703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20233_ clknet_leaf_66_clk _01177_ net1476 vssd1 vssd1 vccd1 vccd1 ag2.body\[167\]
+ sky130_fd_sc_hd__dfrtp_4
Xhold743 control.body\[716\] vssd1 vssd1 vccd1 vccd1 net2305 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold754 control.body\[878\] vssd1 vssd1 vccd1 vccd1 net2316 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14143__A net1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold765 control.body\[1042\] vssd1 vssd1 vccd1 vccd1 net2327 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1123_A net1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold776 control.body\[1063\] vssd1 vssd1 vccd1 vccd1 net2338 sky130_fd_sc_hd__dlygate4sd3_1
Xhold787 control.body\[710\] vssd1 vssd1 vccd1 vccd1 net2349 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09237__A net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09975_ _04421_ _04632_ net892 vssd1 vssd1 vccd1 vccd1 _04948_ sky130_fd_sc_hd__o21ai_2
Xhold798 control.body\[643\] vssd1 vssd1 vccd1 vccd1 net2360 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20164_ clknet_leaf_95_clk _01108_ net1440 vssd1 vssd1 vccd1 vccd1 ag2.body\[226\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA_fanout583_A net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13982__A _06240_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20095_ clknet_leaf_78_clk _01039_ net1492 vssd1 vssd1 vccd1 vccd1 ag2.body\[301\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA_fanout1009_X net1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17173__B net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout371_X net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout750_A net751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19291__CLK clknet_leaf_98_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1492_A net1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout848_A net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09243__Y _04268_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17741__X _03420_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16984__A2 net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1280_X net1280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11007__A _04425_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10750_ _05711_ _05712_ _05717_ _05722_ vssd1 vssd1 vccd1 vccd1 _05723_ sky130_fd_sc_hd__or4_1
XFILLER_0_138_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16736__A2 net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09700__A ag2.body\[67\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09409_ img_gen.updater.commands.mode\[2\] _04387_ vssd1 vssd1 vccd1 vccd1 _04389_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_94_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10681_ _05652_ _05653_ _05645_ vssd1 vssd1 vccd1 vccd1 _05654_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout803_X net803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_137 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12420_ net767 _06477_ net549 vssd1 vssd1 vccd1 vccd1 _07382_ sky130_fd_sc_hd__o21a_1
XFILLER_0_118_660 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xclkbuf_4_7__f_clk clknet_3_3_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_7__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_117_181 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12351_ _07253_ _07285_ vssd1 vssd1 vccd1 vccd1 _07318_ sky130_fd_sc_hd__nor2_1
XFILLER_0_23_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_75_2602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_1484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16533__A _02211_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_2613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_2624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_1295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11302_ net1194 control.body\[681\] vssd1 vssd1 vccd1 vccd1 _06275_ sky130_fd_sc_hd__xor2_1
X_15070_ net2613 net152 _01560_ net2426 vssd1 vssd1 vccd1 vccd1 _00397_ sky130_fd_sc_hd__a22o_1
XFILLER_0_121_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12282_ img_gen.updater.commands.cmd_num\[0\] _07231_ vssd1 vssd1 vccd1 vccd1 _07252_
+ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_56_2023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_1440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_56_2034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_56_2045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14021_ net987 ag2.body\[25\] vssd1 vssd1 vccd1 vccd1 _08182_ sky130_fd_sc_hd__xor2_1
XANTENNA__17449__B1 net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11233_ _06197_ _06198_ _06204_ _06205_ vssd1 vssd1 vccd1 vccd1 _06206_ sky130_fd_sc_hd__or4_1
XFILLER_0_82_1495 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11164_ _06126_ _06127_ _06128_ _06129_ _06136_ vssd1 vssd1 vccd1 vccd1 _06137_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_8_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_1509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10115_ _05052_ _05057_ _05067_ _05087_ vssd1 vssd1 vccd1 vccd1 _05088_ sky130_fd_sc_hd__o31a_1
XANTENNA__13892__A _05813_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18760_ clknet_leaf_16_clk img_gen.tracker.next_frame\[198\] net1315 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[198\] sky130_fd_sc_hd__dfrtp_1
X_15972_ ag2.body\[143\] net212 _01658_ ag2.body\[135\] vssd1 vssd1 vccd1 vccd1 _01201_
+ sky130_fd_sc_hd__a22o_1
X_11095_ ag2.body\[426\] net1176 vssd1 vssd1 vccd1 vccd1 _06068_ sky130_fd_sc_hd__or2_1
XANTENNA__10101__C_N net915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_2417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17711_ obsg2.obstacleArray\[132\] obsg2.obstacleArray\[133\] obsg2.obstacleArray\[134\]
+ obsg2.obstacleArray\[135\] net448 net392 vssd1 vssd1 vccd1 vccd1 _03390_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_69_2428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10046_ net1131 control.body\[900\] vssd1 vssd1 vccd1 vccd1 _05019_ sky130_fd_sc_hd__xor2_1
X_14923_ net2619 net177 _01543_ net2232 vssd1 vssd1 vccd1 vccd1 _00267_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_69_2439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18691_ clknet_leaf_28_clk img_gen.tracker.next_frame\[129\] net1336 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[129\] sky130_fd_sc_hd__dfrtp_1
Xhold70 img_gen.tracker.frame\[332\] vssd1 vssd1 vccd1 vccd1 net1632 sky130_fd_sc_hd__dlygate4sd3_1
Xhold81 img_gen.tracker.frame\[51\] vssd1 vssd1 vccd1 vccd1 net1643 sky130_fd_sc_hd__dlygate4sd3_1
X_17642_ _04049_ net884 net695 ag2.body\[167\] _03320_ vssd1 vssd1 vccd1 vccd1 _03321_
+ sky130_fd_sc_hd__a221o_1
Xhold92 img_gen.tracker.frame\[4\] vssd1 vssd1 vccd1 vccd1 net1654 sky130_fd_sc_hd__dlygate4sd3_1
X_14854_ _08300_ _08301_ _08305_ _08862_ _01521_ vssd1 vssd1 vccd1 vccd1 _01525_ sky130_fd_sc_hd__o311a_1
XFILLER_0_89_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19784__CLK clknet_leaf_127_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1520 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13805_ net1167 _08105_ _08106_ _08104_ vssd1 vssd1 vccd1 vccd1 _00076_ sky130_fd_sc_hd__a22o_1
X_17573_ ag2.body\[339\] net720 net713 ag2.body\[340\] vssd1 vssd1 vccd1 vccd1 _03252_
+ sky130_fd_sc_hd__o22a_1
XANTENNA__13116__B _07639_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11997_ img_gen.tracker.frame\[427\] net545 _06968_ net571 vssd1 vssd1 vccd1 vccd1
+ _06969_ sky130_fd_sc_hd__o211a_1
X_14785_ _01453_ _01454_ _01455_ vssd1 vssd1 vccd1 vccd1 _01456_ sky130_fd_sc_hd__or3_1
XFILLER_0_133_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09457__A3 net640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19312_ clknet_leaf_99_clk _00256_ net1443 vssd1 vssd1 vccd1 vccd1 control.body\[1086\]
+ sky130_fd_sc_hd__dfrtp_1
X_16524_ net536 _02052_ vssd1 vssd1 vccd1 vccd1 _02203_ sky130_fd_sc_hd__or2_1
XFILLER_0_86_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10948_ net907 _04758_ net641 vssd1 vssd1 vccd1 vccd1 _05921_ sky130_fd_sc_hd__a21oi_2
X_13736_ _04272_ img_gen.updater.commands.cmd_num\[0\] _07207_ vssd1 vssd1 vccd1 vccd1
+ _08057_ sky130_fd_sc_hd__or3_1
XFILLER_0_15_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12955__B net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14738__A1 net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19243_ clknet_leaf_75_clk _00187_ net1482 vssd1 vssd1 vccd1 vccd1 ag2.body\[106\]
+ sky130_fd_sc_hd__dfrtp_4
X_16455_ _02120_ _02133_ _02076_ vssd1 vssd1 vccd1 vccd1 _02134_ sky130_fd_sc_hd__mux2_1
XANTENNA__14738__B2 net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_1627 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13667_ _08015_ _08017_ vssd1 vssd1 vccd1 vccd1 obsrand1.next_randY\[2\] sky130_fd_sc_hd__nor2_1
XFILLER_0_112_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10756__A net1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10879_ ag2.body\[535\] net1059 vssd1 vssd1 vccd1 vccd1 _05852_ sky130_fd_sc_hd__xor2_1
XANTENNA__14228__A net980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12674__C _06671_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15406_ net2444 net80 _01581_ control.body\[639\] vssd1 vssd1 vccd1 vccd1 _00697_
+ sky130_fd_sc_hd__a22o_1
X_19174_ clknet_leaf_21_clk _00118_ net1364 vssd1 vssd1 vccd1 vccd1 ag2.body\[37\]
+ sky130_fd_sc_hd__dfrtp_4
X_12618_ net276 _07509_ _07510_ net2000 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[65\]
+ sky130_fd_sc_hd__a22o_1
X_13598_ control.divider.fsm.current_mode\[2\] control.divider.count\[14\] control.divider.count\[15\]
+ _03961_ vssd1 vssd1 vccd1 vccd1 _07973_ sky130_fd_sc_hd__o211a_1
X_16386_ net497 _02061_ vssd1 vssd1 vccd1 vccd1 _02065_ sky130_fd_sc_hd__nor2_4
XFILLER_0_6_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11647__S1 net507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18125_ net526 _03698_ vssd1 vssd1 vccd1 vccd1 _01313_ sky130_fd_sc_hd__and2_1
XFILLER_0_124_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15337_ control.body\[696\] net71 _01590_ net2364 vssd1 vssd1 vccd1 vccd1 _00634_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_5_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12549_ net2073 net652 _07473_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[33\]
+ sky130_fd_sc_hd__and3_1
XFILLER_0_129_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19164__CLK clknet_leaf_52_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_1 _03230_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18056_ obsg2.obstacleArray\[38\] _03653_ net522 vssd1 vssd1 vccd1 vccd1 _01289_
+ sky130_fd_sc_hd__o21a_1
X_15268_ net2557 net109 _01582_ control.body\[755\] vssd1 vssd1 vccd1 vccd1 _00573_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__16162__B net431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_1547 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17007_ ag2.body\[498\] net863 vssd1 vssd1 vccd1 vccd1 _02686_ sky130_fd_sc_hd__xor2_1
XANTENNA__11587__A net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14219_ net819 ag2.body\[395\] ag2.body\[396\] net813 vssd1 vssd1 vccd1 vccd1 _08380_
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_112_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15199_ control.body\[831\] net94 _01573_ net2345 vssd1 vssd1 vccd1 vccd1 _00513_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_46_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout508 _06467_ vssd1 vssd1 vccd1 vccd1 net508 sky130_fd_sc_hd__clkbuf_4
Xfanout519 _04396_ vssd1 vssd1 vccd1 vccd1 net519 sky130_fd_sc_hd__buf_4
XFILLER_0_61_1579 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09760_ _04729_ _04730_ _04731_ _04732_ vssd1 vssd1 vccd1 vccd1 _04733_ sky130_fd_sc_hd__a22o_1
X_18958_ clknet_leaf_7_clk img_gen.tracker.next_frame\[396\] net1266 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[396\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__13477__A1 net230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1300 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17909_ net350 _03533_ vssd1 vssd1 vccd1 vccd1 _03544_ sky130_fd_sc_hd__nor2_1
XANTENNA__20291__CLK clknet_leaf_37_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09691_ ag2.body\[68\] net1139 vssd1 vssd1 vccd1 vccd1 _04664_ sky130_fd_sc_hd__or2_1
XANTENNA__15506__B net65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18889_ clknet_leaf_26_clk img_gen.tracker.next_frame\[327\] net1342 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[327\] sky130_fd_sc_hd__dfrtp_1
Xfanout1090 net1091 vssd1 vssd1 vccd1 vccd1 net1090 sky130_fd_sc_hd__clkbuf_4
XANTENNA__16415__A1 net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13229__A1 net263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10160__B1 net643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16966__A2 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_1388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13026__B _07535_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_98_3303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_98_3314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12865__B net309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_3325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14729__B2 net1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_314 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14138__A net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout429_A _01735_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1073_A net1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11114__X _06087_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19507__CLK clknet_leaf_113_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_1394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09125_ ag2.body\[420\] vssd1 vssd1 vccd1 vccd1 _04150_ sky130_fd_sc_hd__inv_2
XFILLER_0_60_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17679__B1 net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17143__A2 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1240_A net1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1338_A net1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09056_ ag2.body\[250\] vssd1 vssd1 vccd1 vccd1 _04081_ sky130_fd_sc_hd__inv_2
XFILLER_0_66_1468 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout798_A net805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17736__X _03415_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09238__Y _04263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold540 img_gen.tracker.frame\[502\] vssd1 vssd1 vccd1 vccd1 net2102 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold551 control.body\[768\] vssd1 vssd1 vccd1 vccd1 net2113 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1126_X net1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11715__A1 net566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_3_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold562 img_gen.tracker.frame\[286\] vssd1 vssd1 vccd1 vccd1 net2124 sky130_fd_sc_hd__dlygate4sd3_1
X_20216_ clknet_leaf_60_clk _01160_ net1466 vssd1 vssd1 vccd1 vccd1 ag2.body\[182\]
+ sky130_fd_sc_hd__dfrtp_4
Xhold573 control.body\[771\] vssd1 vssd1 vccd1 vccd1 net2135 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_880 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_1300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16103__B1 net374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold584 _00220_ vssd1 vssd1 vccd1 vccd1 net2146 sky130_fd_sc_hd__dlygate4sd3_1
Xhold595 control.body\[1112\] vssd1 vssd1 vccd1 vccd1 net2157 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout965_A net967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout586_X net586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_15__f_clk clknet_3_7_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_15__leaf_clk
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__16654__A1 net362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16800__B net363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20147_ clknet_leaf_100_clk _01091_ net1444 vssd1 vssd1 vccd1 vccd1 ag2.body\[241\]
+ sky130_fd_sc_hd__dfrtp_4
X_09958_ _04922_ _04929_ _04930_ _04916_ _04903_ vssd1 vssd1 vccd1 vccd1 _04931_ sky130_fd_sc_hd__o32a_1
XANTENNA__13468__A1 net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20078_ clknet_leaf_77_clk _01022_ net1491 vssd1 vssd1 vccd1 vccd1 ag2.body\[316\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA_fanout753_X net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15416__B net63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09889_ _04446_ net634 vssd1 vssd1 vccd1 vccd1 _04862_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout1495_X net1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11920_ img_gen.tracker.frame\[328\] net606 net551 img_gen.tracker.frame\[331\] _06891_
+ vssd1 vssd1 vccd1 vccd1 _06892_ sky130_fd_sc_hd__o221a_1
XFILLER_0_87_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16957__A2 net700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11851_ _06724_ net382 vssd1 vssd1 vccd1 vccd1 _06823_ sky130_fd_sc_hd__nand2_1
XANTENNA__17631__B net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout920_X net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16528__A net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10802_ _05771_ _05772_ _05773_ _05774_ _05770_ vssd1 vssd1 vccd1 vccd1 _05775_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_16_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14570_ _08723_ _08724_ _08725_ _08726_ vssd1 vssd1 vccd1 vccd1 _08731_ sky130_fd_sc_hd__or4_1
XFILLER_0_71_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11782_ img_gen.tracker.frame\[176\] net548 vssd1 vssd1 vccd1 vccd1 _06754_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_0_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16709__A2 net492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09430__A net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13521_ net2106 net655 _07919_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[559\]
+ sky130_fd_sc_hd__and3_1
X_10733_ ag2.body\[254\] net1086 vssd1 vssd1 vccd1 vccd1 _05706_ sky130_fd_sc_hd__nor2_1
XANTENNA__15917__B1 _01652_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19187__CLK clknet_leaf_53_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_1495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16240_ _01918_ vssd1 vssd1 vccd1 vccd1 _01919_ sky130_fd_sc_hd__inv_2
X_13452_ net235 _07892_ _07893_ net1860 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[516\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_14_1570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_799 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14196__A2 ag2.body\[161\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10664_ net1202 control.body\[881\] vssd1 vssd1 vccd1 vccd1 _05637_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10295__B net1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12403_ _07300_ _07364_ _07365_ _07366_ vssd1 vssd1 vccd1 vccd1 net28 sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_58_2107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16171_ obsg2.obstacleArray\[30\] obsg2.obstacleArray\[31\] net428 vssd1 vssd1 vccd1
+ vccd1 _01850_ sky130_fd_sc_hd__mux2_1
XANTENNA__10863__X _05836_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13383_ net670 _07866_ vssd1 vssd1 vccd1 vccd1 _07867_ sky130_fd_sc_hd__nor2_1
XANTENNA__12791__A net316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10595_ net1171 control.body\[826\] vssd1 vssd1 vccd1 vccd1 _05568_ sky130_fd_sc_hd__xor2_1
XFILLER_0_134_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_674 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15122_ control.body\[890\] net103 _01565_ net2527 vssd1 vssd1 vccd1 vccd1 _00444_
+ sky130_fd_sc_hd__a22o_1
X_12334_ _06932_ _06985_ _07148_ _06825_ vssd1 vssd1 vccd1 vccd1 _07301_ sky130_fd_sc_hd__o31a_1
XFILLER_0_51_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19930_ clknet_leaf_51_clk _00874_ net1368 vssd1 vssd1 vccd1 vccd1 ag2.body\[456\]
+ sky130_fd_sc_hd__dfrtp_2
X_15053_ control.body\[956\] net150 _01558_ net2279 vssd1 vssd1 vccd1 vccd1 _00382_
+ sky130_fd_sc_hd__a22o_1
X_12265_ img_gen.updater.commands.count\[8\] img_gen.updater.commands.count\[9\] img_gen.updater.commands.count\[7\]
+ vssd1 vssd1 vccd1 vccd1 _07235_ sky130_fd_sc_hd__and3_1
XFILLER_0_32_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_128_Right_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14004_ _08161_ _08163_ _08164_ _08162_ vssd1 vssd1 vccd1 vccd1 _08165_ sky130_fd_sc_hd__or4b_1
XFILLER_0_120_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11216_ net1149 control.body\[843\] vssd1 vssd1 vccd1 vccd1 _06189_ sky130_fd_sc_hd__xnor2_1
X_19861_ clknet_leaf_94_clk _00805_ net1436 vssd1 vssd1 vccd1 vccd1 ag2.body\[531\]
+ sky130_fd_sc_hd__dfrtp_4
X_12196_ _07151_ _07152_ _07166_ _07167_ vssd1 vssd1 vccd1 vccd1 _07168_ sky130_fd_sc_hd__or4_1
XFILLER_0_128_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18812_ clknet_leaf_3_clk img_gen.tracker.next_frame\[250\] net1259 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[250\] sky130_fd_sc_hd__dfrtp_1
X_11147_ _06112_ _06115_ _06118_ _06119_ vssd1 vssd1 vccd1 vccd1 _06120_ sky130_fd_sc_hd__or4_1
XANTENNA__16202__S net376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19792_ clknet_leaf_127_clk _00736_ net1328 vssd1 vssd1 vccd1 vccd1 ag2.body\[606\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__13459__A1 net281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1339 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18743_ clknet_leaf_139_clk img_gen.tracker.next_frame\[181\] net1256 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[181\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09605__A net1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15955_ _05237_ net60 vssd1 vssd1 vccd1 vccd1 _01657_ sky130_fd_sc_hd__nor2_2
X_11078_ ag2.body\[539\] net1158 vssd1 vssd1 vccd1 vccd1 _06051_ sky130_fd_sc_hd__xor2_1
X_10029_ ag2.body\[509\] net756 net746 ag2.body\[511\] vssd1 vssd1 vccd1 vccd1 _05002_
+ sky130_fd_sc_hd__a22o_1
X_14906_ net2577 net178 _01541_ control.body\[1074\] vssd1 vssd1 vccd1 vccd1 _00252_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__13127__A net343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18674_ clknet_leaf_27_clk img_gen.tracker.next_frame\[112\] net1340 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[112\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_56_1626 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15886_ ag2.body\[210\] net184 _01649_ ag2.body\[202\] vssd1 vssd1 vccd1 vccd1 _01124_
+ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_90_Left_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17625_ _03302_ _03303_ _03301_ vssd1 vssd1 vccd1 vccd1 _03304_ sky130_fd_sc_hd__or3b_1
XFILLER_0_91_1539 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14837_ _08475_ _08479_ _08852_ _08904_ _08346_ vssd1 vssd1 vccd1 vccd1 _01508_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_99_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15620__A2 net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17556_ ag2.body\[358\] net945 vssd1 vssd1 vccd1 vccd1 _03235_ sky130_fd_sc_hd__xor2_1
X_14768_ net1011 ag2.body\[103\] vssd1 vssd1 vccd1 vccd1 _08929_ sky130_fd_sc_hd__xor2_1
X_16507_ obsg2.obstacleArray\[14\] net456 vssd1 vssd1 vccd1 vccd1 _02186_ sky130_fd_sc_hd__or2_1
XFILLER_0_89_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13719_ track.current_collision _08036_ track.highScore\[7\] vssd1 vssd1 vccd1 vccd1
+ _08053_ sky130_fd_sc_hd__a21oi_4
X_17487_ ag2.body\[361\] net734 net693 ag2.body\[367\] vssd1 vssd1 vccd1 vccd1 _03166_
+ sky130_fd_sc_hd__a22o_1
X_14699_ net830 ag2.body\[322\] _04112_ net1012 _08859_ vssd1 vssd1 vccd1 vccd1 _08860_
+ sky130_fd_sc_hd__o221a_1
X_19226_ clknet_leaf_75_clk _00170_ net1482 vssd1 vssd1 vccd1 vccd1 ag2.body\[89\]
+ sky130_fd_sc_hd__dfrtp_4
X_16438_ obsg2.obstacleArray\[90\] obsg2.obstacleArray\[91\] net459 vssd1 vssd1 vccd1
+ vccd1 _02117_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18554__CLK clknet_leaf_37_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19157_ clknet_leaf_50_clk _00101_ net1369 vssd1 vssd1 vccd1 vccd1 ag2.body\[21\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_5_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16369_ _01912_ _02042_ _02046_ _01919_ _02038_ vssd1 vssd1 vccd1 vccd1 _02048_ sky130_fd_sc_hd__a311o_1
X_18108_ net44 _03687_ vssd1 vssd1 vccd1 vccd1 _03688_ sky130_fd_sc_hd__nor2_1
XFILLER_0_81_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19088_ clknet_leaf_9_clk img_gen.tracker.next_frame\[526\] net1272 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[526\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_44_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18039_ obsg2.obstacleArray\[32\] _03642_ net521 vssd1 vssd1 vccd1 vccd1 _01283_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_83_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_688 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19197__RESET_B net1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout305 _07445_ vssd1 vssd1 vccd1 vccd1 net305 sky130_fd_sc_hd__clkbuf_4
Xfanout316 _07428_ vssd1 vssd1 vccd1 vccd1 net316 sky130_fd_sc_hd__buf_4
X_20001_ clknet_leaf_66_clk _00945_ net1471 vssd1 vssd1 vccd1 vccd1 ag2.body\[399\]
+ sky130_fd_sc_hd__dfrtp_2
Xfanout327 net328 vssd1 vssd1 vccd1 vccd1 net327 sky130_fd_sc_hd__clkbuf_2
X_09812_ net786 control.body\[1048\] net895 vssd1 vssd1 vccd1 vccd1 _04785_ sky130_fd_sc_hd__o21ai_1
Xfanout338 net340 vssd1 vssd1 vccd1 vccd1 net338 sky130_fd_sc_hd__buf_2
Xfanout349 _01731_ vssd1 vssd1 vccd1 vccd1 net349 sky130_fd_sc_hd__clkbuf_2
XANTENNA__16112__S net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09515__A net1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11679__A_N net1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09743_ ag2.body\[352\] net788 net763 ag2.body\[356\] _04715_ vssd1 vssd1 vccd1 vccd1
+ _04716_ sky130_fd_sc_hd__a221o_1
XANTENNA__11764__B net1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15236__B net63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_129_Left_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout281_A net282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13037__A net342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09674_ net894 _04646_ vssd1 vssd1 vccd1 vccd1 _04647_ sky130_fd_sc_hd__nor2_2
XFILLER_0_90_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_1185 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1190_A net1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12876__A net339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout546_A net547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09521__Y _04494_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1592 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10396__A net1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout713_A net714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1076_X net1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1455_A net1465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20187__CLK clknet_leaf_88_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_138_Left_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19967__RESET_B net1470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout501_X net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1243_X net1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09108_ ag2.body\[376\] vssd1 vssd1 vccd1 vccd1 _04133_ sky130_fd_sc_hd__inv_2
XANTENNA__13500__A _07607_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10380_ ag2.body\[109\] net1115 vssd1 vssd1 vccd1 vccd1 _05353_ sky130_fd_sc_hd__xor2_1
XFILLER_0_102_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09039_ ag2.body\[202\] vssd1 vssd1 vccd1 vccd1 _04064_ sky130_fd_sc_hd__inv_2
XFILLER_0_66_1298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13689__A1 net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12050_ img_gen.tracker.frame\[264\] net628 net609 img_gen.tracker.frame\[267\] vssd1
+ vssd1 vccd1 vccd1 _07022_ sky130_fd_sc_hd__a22o_1
Xhold370 img_gen.tracker.frame\[138\] vssd1 vssd1 vccd1 vccd1 net1932 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout870_X net870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17626__B net949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold381 img_gen.tracker.frame\[434\] vssd1 vssd1 vccd1 vccd1 net1943 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout968_X net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16088__C1 _01743_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold392 img_gen.tracker.frame\[49\] vssd1 vssd1 vccd1 vccd1 net1954 sky130_fd_sc_hd__dlygate4sd3_1
X_11001_ net779 control.body\[1081\] control.body\[1083\] net769 vssd1 vssd1 vccd1
+ vccd1 _05974_ sky130_fd_sc_hd__a22o_1
XANTENNA__14331__A net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20454__RESET_B net1356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout850 net852 vssd1 vssd1 vccd1 vccd1 net850 sky130_fd_sc_hd__buf_4
XANTENNA__10911__A2 _05883_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout861 net862 vssd1 vssd1 vccd1 vccd1 net861 sky130_fd_sc_hd__buf_4
XANTENNA__11674__B _06644_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout872 obsg2.randCord\[1\] vssd1 vssd1 vccd1 vccd1 net872 sky130_fd_sc_hd__buf_4
Xfanout883 net884 vssd1 vssd1 vccd1 vccd1 net883 sky130_fd_sc_hd__buf_4
XFILLER_0_99_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout894 control.body_update.curr_length\[7\] vssd1 vssd1 vccd1 vccd1 net894 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12489__C net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15740_ _05253_ net60 vssd1 vssd1 vccd1 vccd1 _01634_ sky130_fd_sc_hd__nor2_2
X_12952_ net339 _07487_ vssd1 vssd1 vccd1 vccd1 _07673_ sky130_fd_sc_hd__and2_1
XANTENNA__12664__A2 _07536_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1070 control.body\[821\] vssd1 vssd1 vccd1 vccd1 net2632 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1081 control.body\[1009\] vssd1 vssd1 vccd1 vccd1 net2643 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11903_ net438 _06867_ _06874_ _06691_ vssd1 vssd1 vccd1 vccd1 _06875_ sky130_fd_sc_hd__a31o_1
Xhold1092 control.body\[624\] vssd1 vssd1 vccd1 vccd1 net2654 sky130_fd_sc_hd__dlygate4sd3_1
X_15671_ ag2.body\[402\] net142 _01626_ ag2.body\[394\] vssd1 vssd1 vccd1 vccd1 _00932_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12786__A net669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12883_ net245 _07641_ _07642_ net2099 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[198\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_119_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17410_ ag2.body\[281\] net875 vssd1 vssd1 vccd1 vccd1 _03089_ sky130_fd_sc_hd__xnor2_1
X_14622_ _08779_ _08780_ _08782_ vssd1 vssd1 vccd1 vccd1 _08783_ sky130_fd_sc_hd__nand3b_2
XFILLER_0_115_1546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18390_ _03808_ _03872_ _03879_ _03794_ vssd1 vssd1 vccd1 vccd1 _03880_ sky130_fd_sc_hd__a211oi_1
X_11834_ img_gen.tracker.frame\[569\] net605 net588 img_gen.tracker.frame\[575\] vssd1
+ vssd1 vccd1 vccd1 _06806_ sky130_fd_sc_hd__o22a_1
XFILLER_0_23_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18001__B1 net533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17341_ _03970_ net960 vssd1 vssd1 vccd1 vccd1 _03020_ sky130_fd_sc_hd__nand2_1
XFILLER_0_16_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__18577__CLK clknet_leaf_15_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14553_ net1000 ag2.body\[64\] vssd1 vssd1 vccd1 vccd1 _08714_ sky130_fd_sc_hd__xor2_1
X_11765_ img_gen.tracker.frame\[65\] net596 net579 img_gen.tracker.frame\[71\] _06736_
+ vssd1 vssd1 vccd1 vccd1 _06737_ sky130_fd_sc_hd__o221a_1
XFILLER_0_126_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13504_ net276 _07912_ _07913_ net1872 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[548\]
+ sky130_fd_sc_hd__a22o_1
X_10716_ ag2.body\[622\] net1078 vssd1 vssd1 vccd1 vccd1 _05689_ sky130_fd_sc_hd__xor2_1
X_17272_ ag2.body\[557\] net947 vssd1 vssd1 vccd1 vccd1 _02951_ sky130_fd_sc_hd__xor2_1
X_14484_ _08642_ _08643_ _08644_ vssd1 vssd1 vccd1 vccd1 _08645_ sky130_fd_sc_hd__or3_2
X_11696_ net469 _06657_ _06661_ _06667_ vssd1 vssd1 vccd1 vccd1 _06668_ sky130_fd_sc_hd__o211a_1
XANTENNA__18192__B net41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19011_ clknet_leaf_1_clk img_gen.tracker.next_frame\[449\] net1244 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[449\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16223_ _01725_ _01888_ _01900_ vssd1 vssd1 vccd1 vccd1 _01902_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_82_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10647_ ag2.body\[287\] net1066 vssd1 vssd1 vccd1 vccd1 _05620_ sky130_fd_sc_hd__or2_1
X_13435_ _07572_ net302 vssd1 vssd1 vccd1 vccd1 _07886_ sky130_fd_sc_hd__nor2_1
XFILLER_0_67_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14506__A net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17107__A2 net732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_617 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13410__A _07558_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16154_ obsg2.obstacleArray\[4\] net427 net374 _01832_ vssd1 vssd1 vccd1 vccd1 _01833_
+ sky130_fd_sc_hd__o211a_1
X_13366_ net274 _07858_ _07859_ net2149 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[464\]
+ sky130_fd_sc_hd__a22o_1
X_10578_ _05547_ _05548_ _05549_ _05550_ vssd1 vssd1 vccd1 vccd1 _05551_ sky130_fd_sc_hd__a22o_1
XFILLER_0_84_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15105_ net2565 net145 _01564_ control.body\[898\] vssd1 vssd1 vccd1 vccd1 _00428_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_126_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12317_ _04389_ _07232_ vssd1 vssd1 vccd1 vccd1 _07284_ sky130_fd_sc_hd__nand2_1
X_16085_ obsg2.obstacleArray\[112\] obsg2.obstacleArray\[113\] net423 vssd1 vssd1
+ vccd1 vccd1 _01764_ sky130_fd_sc_hd__mux2_1
X_13297_ net280 _07831_ _07832_ net1717 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[422\]
+ sky130_fd_sc_hd__a22o_1
X_19913_ clknet_leaf_54_clk _00857_ net1457 vssd1 vssd1 vccd1 vccd1 ag2.body\[487\]
+ sky130_fd_sc_hd__dfrtp_4
X_12248_ img_gen.updater.commands.cmd_num\[1\] _07217_ _07187_ vssd1 vssd1 vccd1 vccd1
+ _07218_ sky130_fd_sc_hd__mux2_2
X_15036_ net2239 net152 _01557_ net2296 vssd1 vssd1 vccd1 vccd1 _00366_ sky130_fd_sc_hd__a22o_1
XFILLER_0_23_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19202__CLK clknet_leaf_88_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19844_ clknet_leaf_92_clk _00788_ net1412 vssd1 vssd1 vccd1 vccd1 ag2.body\[546\]
+ sky130_fd_sc_hd__dfrtp_4
X_12179_ net1128 ag2.apple_cord\[4\] vssd1 vssd1 vccd1 vccd1 _07151_ sky130_fd_sc_hd__xor2_1
XFILLER_0_120_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11584__B net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19775_ clknet_leaf_19_clk _00719_ net1321 vssd1 vssd1 vccd1 vccd1 ag2.body\[621\]
+ sky130_fd_sc_hd__dfrtp_4
X_16987_ ag2.body\[91\] net853 vssd1 vssd1 vccd1 vccd1 _02666_ sky130_fd_sc_hd__or2_1
X_18726_ clknet_leaf_142_clk img_gen.tracker.next_frame\[164\] net1257 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[164\] sky130_fd_sc_hd__dfrtp_1
X_15938_ ag2.body\[160\] net196 _01653_ ag2.body\[152\] vssd1 vssd1 vccd1 vccd1 _01170_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_3_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10115__B1 _05087_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10666__A1 net762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10666__B2 net1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18657_ clknet_leaf_131_clk img_gen.tracker.next_frame\[95\] net1312 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[95\] sky130_fd_sc_hd__dfrtp_1
X_15869_ ag2.body\[227\] net201 _01647_ ag2.body\[219\] vssd1 vssd1 vccd1 vccd1 _01109_
+ sky130_fd_sc_hd__a22o_1
X_17608_ _04260_ obsg2.obsNeeded\[2\] vssd1 vssd1 vccd1 vccd1 _03287_ sky130_fd_sc_hd__nor2_1
X_09390_ sound_gen.osc1.stayCount\[8\] _04346_ net270 vssd1 vssd1 vccd1 vccd1 _04379_
+ sky130_fd_sc_hd__o21ai_1
X_18588_ clknet_leaf_14_clk img_gen.tracker.next_frame\[26\] net1276 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[26\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_133_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10418__A1 net786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10418__B2 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1022 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17539_ _03213_ _03215_ _03217_ vssd1 vssd1 vccd1 vccd1 _03218_ sky130_fd_sc_hd__or3b_2
XFILLER_0_80_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_703 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12421__A1_N net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_585 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20550_ clknet_leaf_105_clk _01415_ _00024_ vssd1 vssd1 vccd1 vccd1 sound_gen.osc1.stayCount\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_104_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19209_ clknet_leaf_58_clk _00153_ net1473 vssd1 vssd1 vccd1 vccd1 ag2.body\[72\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_105_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_89_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20481_ clknet_leaf_39_clk _01368_ net1352 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[117\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__16107__S net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout127_A net128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_408 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13722__A_N net26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12040__B1 net594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12591__A1 net250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1438 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout1036_A net1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_110_3664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17446__B net940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_3675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11146__A2 net768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_3686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout102 net104 vssd1 vssd1 vccd1 vccd1 net102 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_11_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout113 net114 vssd1 vssd1 vccd1 vccd1 net113 sky130_fd_sc_hd__clkbuf_4
Xfanout124 net128 vssd1 vssd1 vccd1 vccd1 net124 sky130_fd_sc_hd__buf_2
Xfanout135 net144 vssd1 vssd1 vccd1 vccd1 net135 sky130_fd_sc_hd__buf_2
XFILLER_0_61_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1203_A net1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1214 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout146 net183 vssd1 vssd1 vccd1 vccd1 net146 sky130_fd_sc_hd__buf_2
XANTENNA_input1_A en vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout157 net159 vssd1 vssd1 vccd1 vccd1 net157 sky130_fd_sc_hd__buf_2
Xfanout168 net169 vssd1 vssd1 vccd1 vccd1 net168 sky130_fd_sc_hd__clkbuf_2
XANTENNA__14096__A1 net820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout179 net180 vssd1 vssd1 vccd1 vccd1 net179 sky130_fd_sc_hd__buf_2
XFILLER_0_138_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13828__D1 _08114_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout663_A _04394_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout284_X net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14096__B2 net816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09726_ _04018_ net1184 net747 ag2.body\[95\] vssd1 vssd1 vccd1 vccd1 _04699_ sky130_fd_sc_hd__a22o_1
XANTENNA__16468__S0 net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17181__B net948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout830_A net831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout451_X net451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09657_ _04621_ _04624_ _04626_ _04628_ vssd1 vssd1 vccd1 vccd1 _04630_ sky130_fd_sc_hd__or4_1
XANTENNA__11854__B1 net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17585__A2 net738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout928_A net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout549_X net549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1193_X net1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09588_ net1227 control.body\[904\] vssd1 vssd1 vccd1 vccd1 _04561_ sky130_fd_sc_hd__nand2_1
XFILLER_0_96_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout716_X net716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11550_ net1217 net1192 vssd1 vssd1 vccd1 vccd1 _06523_ sky130_fd_sc_hd__and2_1
XFILLER_0_33_1297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10501_ net1060 control.body\[983\] vssd1 vssd1 vccd1 vccd1 _05474_ sky130_fd_sc_hd__xnor2_1
XANTENNA__15899__A2 net133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11481_ _06446_ _06451_ _06452_ _06453_ vssd1 vssd1 vccd1 vccd1 _06454_ sky130_fd_sc_hd__or4_1
XFILLER_0_123_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_1573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13220_ net676 _07799_ vssd1 vssd1 vccd1 vccd1 _07800_ sky130_fd_sc_hd__nor2_1
X_10432_ _05400_ _05401_ _05404_ vssd1 vssd1 vccd1 vccd1 _05405_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09578__A2 net902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12031__B1 net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17908__Y _03543_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10573__B net1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19225__CLK clknet_leaf_75_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10188__A3 net916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13151_ _07497_ net327 net336 vssd1 vssd1 vccd1 vccd1 _07767_ sky130_fd_sc_hd__and3b_1
XFILLER_0_60_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10363_ net773 control.body\[762\] control.body\[765\] net753 vssd1 vssd1 vccd1 vccd1
+ _05336_ sky130_fd_sc_hd__o22a_1
XANTENNA__16541__A net497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12102_ net1215 net1190 img_gen.tracker.frame\[369\] vssd1 vssd1 vccd1 vccd1 _07074_
+ sky130_fd_sc_hd__and3_1
X_13082_ net343 _07564_ vssd1 vssd1 vccd1 vccd1 _07734_ sky130_fd_sc_hd__nor2_1
X_10294_ _04113_ net1236 net764 ag2.body\[332\] _05266_ vssd1 vssd1 vccd1 vccd1 _05267_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_104_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_1371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16910_ _02585_ _02586_ _02588_ vssd1 vssd1 vccd1 vccd1 _02589_ sky130_fd_sc_hd__or3_1
X_12033_ net1216 net1191 img_gen.tracker.frame\[45\] vssd1 vssd1 vccd1 vccd1 _07005_
+ sky130_fd_sc_hd__and3_1
X_17890_ _04398_ _03457_ _03529_ vssd1 vssd1 vccd1 vccd1 _03530_ sky130_fd_sc_hd__nand3_1
XANTENNA__12133__X _07105_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19375__CLK clknet_leaf_93_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_1583 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16841_ ag2.body\[169\] net870 vssd1 vssd1 vccd1 vccd1 _02520_ sky130_fd_sc_hd__nand2_1
XANTENNA_clkbuf_leaf_8_clk_A clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout680 net681 vssd1 vssd1 vccd1 vccd1 net680 sky130_fd_sc_hd__clkbuf_4
XANTENNA__17372__A net927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout691 net695 vssd1 vssd1 vccd1 vccd1 net691 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12098__B1 net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19560_ clknet_leaf_116_clk _00504_ net1389 vssd1 vssd1 vccd1 vccd1 control.body\[838\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16772_ obsg2.obstacleArray\[12\] net492 net483 obsg2.obstacleArray\[13\] _02450_
+ vssd1 vssd1 vccd1 vccd1 _02451_ sky130_fd_sc_hd__a221o_1
X_13984_ ag2.body\[121\] net214 _08159_ ag2.body\[113\] vssd1 vssd1 vccd1 vccd1 _00202_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_92_1623 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18511_ net1513 net1507 vssd1 vssd1 vccd1 vccd1 _00042_ sky130_fd_sc_hd__or2_1
X_15723_ ag2.body\[352\] net197 _01632_ ag2.body\[344\] vssd1 vssd1 vccd1 vccd1 _00978_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_125_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11845__B1 net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19491_ clknet_leaf_113_clk _00435_ net1399 vssd1 vssd1 vccd1 vccd1 control.body\[897\]
+ sky130_fd_sc_hd__dfrtp_1
X_12935_ _07476_ _07639_ vssd1 vssd1 vccd1 vccd1 _07665_ sky130_fd_sc_hd__nor2_1
XFILLER_0_115_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18442_ net464 _03915_ vssd1 vssd1 vccd1 vccd1 _03931_ sky130_fd_sc_hd__nor2_1
XANTENNA__13405__A net313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15654_ ag2.body\[419\] net138 _01624_ ag2.body\[411\] vssd1 vssd1 vccd1 vccd1 _00917_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_92_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_1574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12866_ net675 _07634_ vssd1 vssd1 vccd1 vccd1 _07635_ sky130_fd_sc_hd__nor2_1
XFILLER_0_96_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10748__B net1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14605_ net1012 ag2.body\[135\] vssd1 vssd1 vccd1 vccd1 _08766_ sky130_fd_sc_hd__or2_1
XFILLER_0_69_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19889__RESET_B net1480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13124__B net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18373_ toggle1.bcd_ones\[0\] track.current_collision net464 _08020_ vssd1 vssd1
+ vccd1 vccd1 _03865_ sky130_fd_sc_hd__o211a_1
XFILLER_0_29_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11817_ img_gen.tracker.frame\[398\] net617 net600 img_gen.tracker.frame\[401\] _06788_
+ vssd1 vssd1 vccd1 vccd1 _06789_ sky130_fd_sc_hd__o221a_1
X_15585_ ag2.body\[485\] net130 _01617_ ag2.body\[477\] vssd1 vssd1 vccd1 vccd1 _00855_
+ sky130_fd_sc_hd__a22o_1
X_12797_ net667 _07601_ vssd1 vssd1 vccd1 vccd1 _07602_ sky130_fd_sc_hd__nor2_1
X_17324_ ag2.body\[221\] net952 vssd1 vssd1 vccd1 vccd1 _03003_ sky130_fd_sc_hd__xor2_1
X_14536_ net975 _04082_ _04084_ net1020 _08696_ vssd1 vssd1 vccd1 vccd1 _08697_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_137_4490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11748_ net466 _06673_ vssd1 vssd1 vccd1 vccd1 _06720_ sky130_fd_sc_hd__nand2_1
XFILLER_0_44_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17255_ ag2.body\[550\] net938 vssd1 vssd1 vccd1 vccd1 _02934_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_133_4365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14467_ net1030 ag2.body\[269\] vssd1 vssd1 vccd1 vccd1 _08628_ sky130_fd_sc_hd__xor2_1
XANTENNA__10820__B2 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_133_4376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11679_ net1225 net1199 vssd1 vssd1 vccd1 vccd1 _06651_ sky130_fd_sc_hd__and2b_2
XTAP_TAPCELL_ROW_133_4387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16206_ _01724_ _01870_ _01884_ vssd1 vssd1 vccd1 vccd1 _01885_ sky130_fd_sc_hd__and3b_1
XANTENNA__13140__A _07592_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_1593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_12_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12022__B1 net595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13418_ net257 _07878_ _07879_ net1705 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[496\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__09569__A2 net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17186_ ag2.body\[571\] net849 vssd1 vssd1 vccd1 vccd1 _02865_ sky130_fd_sc_hd__xor2_1
X_14398_ net815 ag2.body\[124\] ag2.body\[127\] net796 _08558_ vssd1 vssd1 vccd1 vccd1
+ _08559_ sky130_fd_sc_hd__o221a_1
XFILLER_0_12_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10483__B net1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11376__A2 net1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16137_ net850 _01815_ _01814_ vssd1 vssd1 vccd1 vccd1 _01816_ sky130_fd_sc_hd__a21oi_2
X_13349_ net228 _07852_ _07853_ net1740 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[453\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_11_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16068_ net377 _01746_ _01745_ net346 vssd1 vssd1 vccd1 vccd1 _01747_ sky130_fd_sc_hd__a211o_1
X_15019_ control.body\[991\] net166 _01553_ control.body\[983\] vssd1 vssd1 vccd1
+ vccd1 _00353_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_55_1987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_1477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_55_1998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19827_ clknet_leaf_124_clk _00771_ net1408 vssd1 vssd1 vccd1 vccd1 ag2.body\[561\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__17803__A3 net939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16597__S _02214_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12089__B1 net557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10004__A net1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19758_ clknet_leaf_129_clk _00702_ net1326 vssd1 vssd1 vccd1 vccd1 control.body\[636\]
+ sky130_fd_sc_hd__dfrtp_1
X_09511_ _04480_ _04482_ _04483_ _04472_ vssd1 vssd1 vccd1 vccd1 _04484_ sky130_fd_sc_hd__or4b_4
XANTENNA__18213__B1 net521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18709_ clknet_leaf_143_clk img_gen.tracker.next_frame\[147\] net1255 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[147\] sky130_fd_sc_hd__dfrtp_1
X_19689_ clknet_leaf_136_clk net2455 net1300 vssd1 vssd1 vccd1 vccd1 control.body\[711\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_91_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15027__B1 _01555_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09442_ _04406_ _04413_ _04414_ vssd1 vssd1 vccd1 vccd1 _04415_ sky130_fd_sc_hd__nor3_1
XFILLER_0_17_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_1117 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16775__B1 net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09373_ sound_gen.osc1.stayCount\[18\] _04367_ _04362_ net271 vssd1 vssd1 vccd1 vccd1
+ _01417_ sky130_fd_sc_hd__o211a_1
XANTENNA__10010__Y _04983_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkload132_A clknet_leaf_73_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14250__A1 net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout244_A net247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14250__B2 net1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20602_ net1534 vssd1 vssd1 vccd1 vccd1 gpio_oeb[14] sky130_fd_sc_hd__buf_2
XFILLER_0_47_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20533_ clknet_leaf_114_clk _01398_ net1398 vssd1 vssd1 vccd1 vccd1 toggle1.bcd_ones\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout411_A net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14146__A net970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_116_3851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1153_A net1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_116_3862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_116_3873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11489__B net1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20464_ clknet_leaf_25_clk _01351_ net1340 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[100\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_112_3726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_112_3737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12564__A1 net245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_3748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20395_ clknet_leaf_42_clk _01282_ net1371 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[31\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_105_1501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1320_A net1324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19398__CLK clknet_leaf_103_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1039_X net1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17176__B net930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout780_A net781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout878_A obsg2.randCord\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout499_X net499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_1582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11709__S net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout1206_X net1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_2490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout666_X net666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09703__A ag2.body\[66\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09709_ ag2.body\[242\] net1183 vssd1 vssd1 vccd1 vccd1 _04682_ sky130_fd_sc_hd__nand2_1
X_10981_ net1150 control.body\[755\] vssd1 vssd1 vccd1 vccd1 _05954_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout833_X net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15018__B1 _01553_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_1353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12720_ net335 _07453_ vssd1 vssd1 vccd1 vccd1 _07564_ sky130_fd_sc_hd__or2_2
XTAP_TAPCELL_ROW_84_2873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16766__B1 net484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_2884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_84_2895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_2748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_2294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_792 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12651_ net242 _07529_ _07530_ net1722 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[78\]
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_80_2759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_4_0__f_clk_X clknet_4_0__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16536__A net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11602_ obsg2.obstacleArray\[17\] obsg2.obstacleArray\[21\] net514 vssd1 vssd1 vccd1
+ vccd1 _06575_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11055__A1 _04427_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_2169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12582_ net666 _07491_ vssd1 vssd1 vccd1 vccd1 _07492_ sky130_fd_sc_hd__nor2_1
X_15370_ control.body\[678\] net69 _01593_ net2241 vssd1 vssd1 vccd1 vccd1 _00664_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__09799__A2 _04519_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14321_ net812 ag2.body\[452\] ag2.body\[454\] net800 vssd1 vssd1 vccd1 vccd1 _08482_
+ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__19229__RESET_B net1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11533_ net1167 net1144 vssd1 vssd1 vccd1 vccd1 _06506_ sky130_fd_sc_hd__nand2_1
XFILLER_0_108_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14056__A net1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17040_ ag2.body\[126\] net701 net694 ag2.body\[127\] vssd1 vssd1 vccd1 vccd1 _02719_
+ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_22_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11464_ ag2.body\[260\] net764 net770 ag2.body\[259\] vssd1 vssd1 vccd1 vccd1 _06437_
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_34_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11399__B net1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14252_ _08410_ _08411_ _08412_ vssd1 vssd1 vccd1 vccd1 _08413_ sky130_fd_sc_hd__or3_2
XFILLER_0_20_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_78_2688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11358__A2 _04238_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_2699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13203_ net676 _07791_ vssd1 vssd1 vccd1 vccd1 _07792_ sky130_fd_sc_hd__nor2_1
X_10415_ _05301_ _05335_ _05359_ _05387_ vssd1 vssd1 vccd1 vccd1 _05388_ sky130_fd_sc_hd__and4_1
X_14183_ net806 ag2.body\[197\] ag2.body\[196\] net811 vssd1 vssd1 vccd1 vccd1 _08344_
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_81_1324 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11395_ _06364_ _06365_ _06366_ _06367_ vssd1 vssd1 vccd1 vccd1 _06368_ sky130_fd_sc_hd__or4_1
XFILLER_0_81_1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10346_ _05314_ _05315_ _05316_ _05318_ vssd1 vssd1 vccd1 vccd1 _05319_ sky130_fd_sc_hd__or4_1
X_13134_ net684 _07758_ vssd1 vssd1 vccd1 vccd1 _07759_ sky130_fd_sc_hd__nor2_1
XANTENNA__10030__A2 net771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17086__B net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18991_ clknet_leaf_7_clk img_gen.tracker.next_frame\[429\] net1265 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[429\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_131_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18765__CLK clknet_leaf_16_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17654__X _03333_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17942_ net318 _03571_ obsg2.obstacleArray\[6\] vssd1 vssd1 vccd1 vccd1 _03572_ sky130_fd_sc_hd__a21oi_1
X_13065_ net340 net330 _07438_ vssd1 vssd1 vccd1 vccd1 _07726_ sky130_fd_sc_hd__and3_2
X_10277_ _05240_ _05241_ _05247_ _05248_ vssd1 vssd1 vccd1 vccd1 _05250_ sky130_fd_sc_hd__a22o_1
XANTENNA__11515__C1 net759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1420 net1423 vssd1 vssd1 vccd1 vccd1 net1420 sky130_fd_sc_hd__clkbuf_4
X_12016_ img_gen.tracker.frame\[228\] net630 net557 img_gen.tracker.frame\[234\] vssd1
+ vssd1 vccd1 vccd1 _06988_ sky130_fd_sc_hd__a22o_1
Xfanout1431 net1432 vssd1 vssd1 vccd1 vccd1 net1431 sky130_fd_sc_hd__clkbuf_4
X_17873_ net2198 _03505_ vssd1 vssd1 vccd1 vccd1 _03516_ sky130_fd_sc_hd__nor2_1
Xfanout1442 net1453 vssd1 vssd1 vccd1 vccd1 net1442 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_126_4180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18198__A _03543_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1453 net1505 vssd1 vssd1 vccd1 vccd1 net1453 sky130_fd_sc_hd__clkbuf_4
XANTENNA__15257__B1 net50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1464 net1465 vssd1 vssd1 vccd1 vccd1 net1464 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_50_1840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1475 net1477 vssd1 vssd1 vccd1 vccd1 net1475 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_122_4033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19612_ clknet_leaf_120_clk _00556_ net1392 vssd1 vssd1 vccd1 vccd1 control.body\[778\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_50_1851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16824_ ag2.body\[231\] net933 vssd1 vssd1 vccd1 vccd1 _02503_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_122_4044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1486 net1493 vssd1 vssd1 vccd1 vccd1 net1486 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_50_1862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1497 net1498 vssd1 vssd1 vccd1 vccd1 net1497 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_122_4055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_1405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12958__B _07639_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_1420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19543_ clknet_leaf_118_clk _00487_ net1388 vssd1 vssd1 vccd1 vccd1 control.body\[853\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_31_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09613__A net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16755_ obsg2.obstacleArray\[44\] net490 net481 obsg2.obstacleArray\[45\] _02433_
+ vssd1 vssd1 vccd1 vccd1 _02434_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_31_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13967_ ag2.body\[106\] net189 _08157_ ag2.body\[98\] vssd1 vssd1 vccd1 vccd1 _00187_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__15009__B1 _01552_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17549__A2 net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15706_ ag2.body\[370\] net141 _01629_ ag2.body\[362\] vssd1 vssd1 vccd1 vccd1 _00964_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__17830__A net824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11294__A1 net742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19474_ clknet_leaf_110_clk net2151 net1418 vssd1 vssd1 vccd1 vccd1 control.body\[912\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12918_ net679 _07656_ vssd1 vssd1 vccd1 vccd1 _07657_ sky130_fd_sc_hd__nor2_1
X_16686_ net358 _02266_ _02270_ _02212_ vssd1 vssd1 vccd1 vccd1 _02365_ sky130_fd_sc_hd__a31o_1
XFILLER_0_0_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11294__B2 _06240_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13898_ ag2.body\[45\] net85 _08149_ ag2.body\[37\] vssd1 vssd1 vccd1 vccd1 _00126_
+ sky130_fd_sc_hd__a22o_1
X_18425_ _08135_ _03913_ _03800_ vssd1 vssd1 vccd1 vccd1 _03914_ sky130_fd_sc_hd__o21ai_1
X_15637_ ag2.body\[436\] net125 _01622_ ag2.body\[428\] vssd1 vssd1 vccd1 vccd1 _00902_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_115_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12849_ net239 _07625_ _07626_ net1990 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[180\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__14232__A1 net996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_4427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14232__B2 net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_135_4438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_4449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18356_ net464 _03785_ vssd1 vssd1 vccd1 vccd1 _03851_ sky130_fd_sc_hd__nor2_1
X_15568_ ag2.body\[503\] net185 _01614_ ag2.body\[495\] vssd1 vssd1 vccd1 vccd1 _00841_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_44_1655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1194 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17307_ ag2.body\[397\] net949 vssd1 vssd1 vccd1 vccd1 _02986_ sky130_fd_sc_hd__nand2_1
XFILLER_0_84_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12794__A1 net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14519_ net821 ag2.body\[315\] ag2.body\[317\] net809 vssd1 vssd1 vccd1 vccd1 _08680_
+ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_20_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18287_ net323 net321 vssd1 vssd1 vccd1 vccd1 _03783_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_25_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15499_ ag2.body\[553\] net113 _01607_ ag2.body\[545\] vssd1 vssd1 vccd1 vccd1 _00779_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_128_1501 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17238_ _02911_ _02912_ _02916_ vssd1 vssd1 vccd1 vccd1 _02917_ sky130_fd_sc_hd__or3_2
XFILLER_0_114_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19540__CLK clknet_leaf_113_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_94_3180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_94_3191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold903 _00607_ vssd1 vssd1 vccd1 vccd1 net2465 sky130_fd_sc_hd__dlygate4sd3_1
Xhold914 img_gen.updater.commands.count\[1\] vssd1 vssd1 vccd1 vccd1 net2476 sky130_fd_sc_hd__dlygate4sd3_1
X_17169_ _02838_ _02845_ _02846_ _02847_ vssd1 vssd1 vccd1 vccd1 _02848_ sky130_fd_sc_hd__or4b_1
XFILLER_0_128_1589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold925 control.body\[637\] vssd1 vssd1 vccd1 vccd1 net2487 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_3055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold936 _00514_ vssd1 vssd1 vccd1 vccd1 net2498 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_720 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_3066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_53_clk_X clknet_leaf_53_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold947 control.body\[860\] vssd1 vssd1 vccd1 vccd1 net2509 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_3077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20180_ clknet_leaf_87_clk _01124_ net1460 vssd1 vssd1 vccd1 vccd1 ag2.body\[210\]
+ sky130_fd_sc_hd__dfrtp_4
Xhold958 _00379_ vssd1 vssd1 vccd1 vccd1 net2520 sky130_fd_sc_hd__dlygate4sd3_1
Xhold969 control.body\[827\] vssd1 vssd1 vccd1 vccd1 net2531 sky130_fd_sc_hd__dlygate4sd3_1
X_09991_ net1193 _04240_ control.body\[735\] net743 _04963_ vssd1 vssd1 vccd1 vccd1
+ _04964_ sky130_fd_sc_hd__a221o_1
XANTENNA__10941__B net1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14299__B2 net814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_11__f_clk_X clknet_4_11__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08942_ ag2.body\[2\] vssd1 vssd1 vccd1 vccd1 _03967_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14417__A1_N net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout194_A net196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_105_3530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09523__A net1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_111_clk_X clknet_leaf_111_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout361_A _02222_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_3405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14471__A1 net975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_3416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_545 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14471__B2 net1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1549 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11117__X _06090_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16748__B1 net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09425_ score_detect.sig_out\[1\] track.last_collision score_detect.N\[1\] vssd1
+ vssd1 vccd1 vccd1 _04402_ sky130_fd_sc_hd__or3b_4
XANTENNA__14223__B2 net833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout247_X net247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1368_A net1369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_118_3913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18638__CLK clknet_leaf_131_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_118_3924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09356_ sound_gen.osc1.stayCount\[15\] sound_gen.osc1.stayCount\[14\] sound_gen.osc1.stayCount\[13\]
+ _04357_ vssd1 vssd1 vccd1 vccd1 _04358_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_118_3935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09287_ _04308_ vssd1 vssd1 vccd1 vccd1 sound_gen.osc1.freq_nxt\[2\] sky130_fd_sc_hd__inv_2
XANTENNA_fanout414_X net414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout1156_X net1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20516_ clknet_leaf_113_clk track.nextHighScore\[6\] net1403 vssd1 vssd1 vccd1 vccd1
+ track.highScore\[6\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16920__B1 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16803__B net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20447_ clknet_leaf_42_clk _01334_ net1371 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[83\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_120_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_1021 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14604__A net1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10200_ ag2.body\[115\] net1164 vssd1 vssd1 vccd1 vccd1 _05173_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_73_2541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11180_ net1154 ag2.body\[179\] vssd1 vssd1 vccd1 vccd1 _06153_ sky130_fd_sc_hd__and2b_1
XFILLER_0_82_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20378_ clknet_leaf_25_clk _01265_ net1345 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[14\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_73_2552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout783_X net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15487__B1 _01605_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10131_ net1148 control.body\[819\] vssd1 vssd1 vccd1 vccd1 _05104_ sky130_fd_sc_hd__xor2_1
XANTENNA__09417__B net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10062_ _05030_ _05032_ _05033_ _05034_ vssd1 vssd1 vccd1 vccd1 _05035_ sky130_fd_sc_hd__or4_2
XANTENNA_fanout950_X net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17634__B net961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15239__B1 _01578_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14870_ net2145 net182 _01537_ control.body\[1106\] vssd1 vssd1 vccd1 vccd1 _00220_
+ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout62_X net62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17353__C ag2.body\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10720__B1 net1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13821_ control.body_update.direction\[2\] control.body_update.direction\[1\] vssd1
+ vssd1 vccd1 vccd1 _08118_ sky130_fd_sc_hd__nand2b_2
XANTENNA__09433__A net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19413__CLK clknet_leaf_103_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_2356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_2367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16540_ net494 _02203_ vssd1 vssd1 vccd1 vccd1 _02219_ sky130_fd_sc_hd__nor2_1
XFILLER_0_15_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10079__A2 net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_2378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13752_ _07240_ _08070_ vssd1 vssd1 vccd1 vccd1 _08071_ sky130_fd_sc_hd__or2_1
XANTENNA__16739__B1 net487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10964_ net919 _04555_ _04599_ _04614_ vssd1 vssd1 vccd1 vccd1 _05937_ sky130_fd_sc_hd__o31ai_1
XANTENNA__14993__B net65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09720__X _04693_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12703_ net310 _07555_ vssd1 vssd1 vccd1 vccd1 _07556_ sky130_fd_sc_hd__nand2_1
X_16471_ net403 _02140_ _02142_ net366 vssd1 vssd1 vccd1 vccd1 _02150_ sky130_fd_sc_hd__o211a_1
XANTENNA__14214__A1 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13683_ _04944_ _05697_ vssd1 vssd1 vccd1 vccd1 _08027_ sky130_fd_sc_hd__and2_1
XANTENNA__14214__B2 net793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14338__X _08499_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10895_ _05862_ _05863_ _05865_ _05867_ vssd1 vssd1 vccd1 vccd1 _05868_ sky130_fd_sc_hd__a211o_1
X_18210_ _03652_ net40 vssd1 vssd1 vccd1 vccd1 _03744_ sky130_fd_sc_hd__nor2_1
X_15422_ control.body\[629\] net84 _01598_ ag2.body\[621\] vssd1 vssd1 vccd1 vccd1
+ _00711_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_14_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12634_ net307 _07519_ vssd1 vssd1 vccd1 vccd1 _07520_ sky130_fd_sc_hd__nor2_1
X_19190_ clknet_leaf_53_clk _00134_ net1366 vssd1 vssd1 vccd1 vccd1 ag2.body\[53\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_14_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_773 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_1443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_14_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18141_ net529 _03709_ vssd1 vssd1 vccd1 vccd1 _01318_ sky130_fd_sc_hd__and2_1
XFILLER_0_109_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15353_ net2658 net72 _01591_ control.body\[687\] vssd1 vssd1 vccd1 vccd1 _00649_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_108_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_1121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12565_ net268 _07481_ _07482_ net1983 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[40\]
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_130_4302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_1555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14304_ net846 ag2.body\[216\] _04070_ net1011 vssd1 vssd1 vccd1 vccd1 _08465_ sky130_fd_sc_hd__o22a_1
XANTENNA__11203__A net1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11516_ net1125 _06471_ _06485_ _06488_ vssd1 vssd1 vccd1 vccd1 _06489_ sky130_fd_sc_hd__o211a_1
X_18072_ net300 _03589_ vssd1 vssd1 vccd1 vccd1 _03664_ sky130_fd_sc_hd__nand2_1
X_15284_ control.body\[745\] net78 _01584_ control.body\[737\] vssd1 vssd1 vccd1 vccd1
+ _00587_ sky130_fd_sc_hd__a22o_1
X_12496_ net617 net440 net473 net560 vssd1 vssd1 vccd1 vccd1 _07442_ sky130_fd_sc_hd__or4_1
XANTENNA__16911__B1 net710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12018__B net1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17023_ _02693_ _02694_ _02695_ _02701_ vssd1 vssd1 vccd1 vccd1 _02702_ sky130_fd_sc_hd__a211o_1
X_14235_ net1042 _04176_ _04177_ net1007 vssd1 vssd1 vccd1 vccd1 _08396_ sky130_fd_sc_hd__a22o_1
X_11447_ _06416_ _06417_ _06418_ _06419_ vssd1 vssd1 vccd1 vccd1 _06420_ sky130_fd_sc_hd__a22o_1
XANTENNA__14514__A net985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09608__A net1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11378_ _04427_ _04695_ net642 vssd1 vssd1 vccd1 vccd1 _06351_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_0_225 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14166_ net980 _04064_ _04066_ net1019 _08326_ vssd1 vssd1 vccd1 vccd1 _08327_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_128_4220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_4231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_4242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13117_ net683 _07750_ vssd1 vssd1 vccd1 vccd1 _07751_ sky130_fd_sc_hd__nor2_1
X_10329_ net638 _04571_ net643 vssd1 vssd1 vccd1 vccd1 _05302_ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_52_1902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14097_ _08249_ _08250_ _08255_ _08257_ vssd1 vssd1 vccd1 vccd1 _08258_ sky130_fd_sc_hd__or4b_1
XTAP_TAPCELL_ROW_52_1913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18974_ clknet_leaf_8_clk img_gen.tracker.next_frame\[412\] net1270 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[412\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_52_1924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_4106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_4117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17925_ _03540_ _03557_ vssd1 vssd1 vccd1 vccd1 _03558_ sky130_fd_sc_hd__and2_1
XFILLER_0_98_1640 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13048_ net387 _07306_ _07638_ vssd1 vssd1 vccd1 vccd1 _07718_ sky130_fd_sc_hd__and3_2
XTAP_TAPCELL_ROW_33_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12969__A net341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1250 net1333 vssd1 vssd1 vccd1 vccd1 net1250 sky130_fd_sc_hd__buf_2
XANTENNA__12700__A1 net258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1261 net1262 vssd1 vssd1 vccd1 vccd1 net1261 sky130_fd_sc_hd__clkbuf_4
XANTENNA__15345__A _05827_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17856_ _03509_ _03510_ vssd1 vssd1 vccd1 vccd1 _01232_ sky130_fd_sc_hd__nor2_1
XANTENNA__09614__Y _04587_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1272 net1287 vssd1 vssd1 vccd1 vccd1 net1272 sky130_fd_sc_hd__buf_2
Xfanout1283 net1286 vssd1 vssd1 vccd1 vccd1 net1283 sky130_fd_sc_hd__clkbuf_2
Xfanout1294 net1296 vssd1 vssd1 vccd1 vccd1 net1294 sky130_fd_sc_hd__clkbuf_4
X_16807_ _04000_ net865 net701 ag2.body\[70\] _02485_ vssd1 vssd1 vccd1 vccd1 _02486_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_59_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17787_ _03461_ _03460_ vssd1 vssd1 vccd1 vccd1 _03464_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_89_843 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14999_ control.body\[1005\] net153 _01551_ control.body\[997\] vssd1 vssd1 vccd1
+ vccd1 _00335_ sky130_fd_sc_hd__a22o_1
XFILLER_0_88_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_80_clk_A clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16738_ obsg2.obstacleArray\[51\] net501 net482 obsg2.obstacleArray\[49\] vssd1 vssd1
+ vccd1 vccd1 _02417_ sky130_fd_sc_hd__a22o_1
XFILLER_0_92_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19526_ clknet_leaf_120_clk _00470_ net1394 vssd1 vssd1 vccd1 vccd1 control.body\[868\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_92_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_1717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20070__CLK clknet_leaf_73_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_46_1728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19457_ clknet_leaf_109_clk _00401_ net1420 vssd1 vssd1 vccd1 vccd1 control.body\[943\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_48_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16669_ obsg2.obstacleArray\[16\] obsg2.obstacleArray\[17\] net447 vssd1 vssd1 vccd1
+ vccd1 _02348_ sky130_fd_sc_hd__mux2_1
XANTENNA__14205__A1 net843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14205__B2 net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15402__B1 _01581_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09210_ net895 vssd1 vssd1 vccd1 vccd1 _04235_ sky130_fd_sc_hd__inv_2
XFILLER_0_57_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18408_ _03890_ _03891_ _03897_ vssd1 vssd1 vccd1 vccd1 _03898_ sky130_fd_sc_hd__a21o_1
X_19388_ clknet_leaf_112_clk _00332_ net1430 vssd1 vssd1 vccd1 vccd1 control.body\[1002\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_17_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_1543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_913 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09141_ ag2.body\[467\] vssd1 vssd1 vccd1 vccd1 _04166_ sky130_fd_sc_hd__inv_2
XFILLER_0_5_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_95_clk_A clknet_4_11__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18339_ _08140_ _03834_ vssd1 vssd1 vccd1 vccd1 _03835_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_96_3242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_96_3253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17155__B1 net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20391__RESET_B net1374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_96_3264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_1606 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_92_3117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09072_ ag2.body\[293\] vssd1 vssd1 vccd1 vccd1 _04097_ sky130_fd_sc_hd__inv_2
XFILLER_0_44_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_92_3128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_92_3139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12519__A1 net226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20301_ clknet_leaf_36_clk net1519 net1347 vssd1 vssd1 vccd1 vccd1 control.divider.count\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_128_1342 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11990__A2 net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold700 control.body\[835\] vssd1 vssd1 vccd1 vccd1 net2262 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout207_A net210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_854 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold711 _00648_ vssd1 vssd1 vccd1 vccd1 net2273 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14424__A net1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13192__A1 net241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12870__C _07444_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold722 control.body\[1033\] vssd1 vssd1 vccd1 vccd1 net2284 sky130_fd_sc_hd__dlygate4sd3_1
X_20232_ clknet_leaf_66_clk _01176_ net1476 vssd1 vssd1 vccd1 vccd1 ag2.body\[166\]
+ sky130_fd_sc_hd__dfrtp_4
Xhold733 control.body\[860\] vssd1 vssd1 vccd1 vccd1 net2295 sky130_fd_sc_hd__dlygate4sd3_1
Xhold744 control.body\[926\] vssd1 vssd1 vccd1 vccd1 net2306 sky130_fd_sc_hd__dlygate4sd3_1
Xhold755 control.body\[1099\] vssd1 vssd1 vccd1 vccd1 net2317 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15469__B1 _01603_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold766 control.body\[885\] vssd1 vssd1 vccd1 vccd1 net2328 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__16666__C1 net360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold777 control.body\[1030\] vssd1 vssd1 vccd1 vccd1 net2339 sky130_fd_sc_hd__dlygate4sd3_1
Xhold788 control.body\[706\] vssd1 vssd1 vccd1 vccd1 net2350 sky130_fd_sc_hd__dlygate4sd3_1
X_20163_ clknet_leaf_82_clk _01107_ net1480 vssd1 vssd1 vccd1 vccd1 ag2.body\[225\]
+ sky130_fd_sc_hd__dfrtp_4
X_09974_ _04632_ _04695_ vssd1 vssd1 vccd1 vccd1 _04947_ sky130_fd_sc_hd__nor2_2
Xhold799 control.body\[754\] vssd1 vssd1 vccd1 vccd1 net2361 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1116_A net1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_33_clk_A clknet_4_5__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13982__B net61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17454__B net960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20094_ clknet_leaf_76_clk _01038_ net1492 vssd1 vssd1 vccd1 vccd1 ag2.body\[300\]
+ sky130_fd_sc_hd__dfrtp_2
XPHY_EDGE_ROW_110_Left_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14692__A1 net1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout576_A net577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14692__B2 net830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16969__B1 net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16433__A2 _02059_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1302 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout364_X net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10399__A net1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout743_A net744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1485_A net1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19586__CLK clknet_leaf_118_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_62_2220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout531_X net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17394__B1 net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout629_X net629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09408_ _04387_ vssd1 vssd1 vccd1 vccd1 _04388_ sky130_fd_sc_hd__inv_2
XANTENNA__15944__A1 ag2.body\[166\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10680_ ag2.body\[349\] net1113 vssd1 vssd1 vccd1 vccd1 _05653_ sky130_fd_sc_hd__or2_1
XANTENNA__09700__B net1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__20408__RESET_B net1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12758__A1 net237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13955__B1 net67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09339_ sound_gen.osc1.stayCount\[3\] sound_gen.osc1.stayCount\[2\] _04342_ vssd1
+ vssd1 vccd1 vccd1 _04343_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_109_Right_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09623__A1 net783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09623__B2 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_106_clk_A clknet_4_10__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12350_ _07304_ _07316_ vssd1 vssd1 vccd1 vccd1 _07317_ sky130_fd_sc_hd__nor2_1
XANTENNA__10233__A2 _05191_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_2603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_193 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__20061__RESET_B net1502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout998_X net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_2614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_75_2625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11301_ net1168 control.body\[682\] vssd1 vssd1 vccd1 vccd1 _06274_ sky130_fd_sc_hd__xor2_1
X_12281_ img_gen.updater.commands.cmd_num\[1\] _07232_ _07248_ _07250_ vssd1 vssd1
+ vccd1 vccd1 _07251_ sky130_fd_sc_hd__a22o_2
XFILLER_0_105_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_56_2024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_2035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_174 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_399 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14020_ _08174_ _08176_ _08179_ _08180_ vssd1 vssd1 vccd1 vccd1 _08181_ sky130_fd_sc_hd__or4b_2
X_11232_ _06195_ _06196_ _06202_ _06203_ vssd1 vssd1 vccd1 vccd1 _06205_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_56_2046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09926__A2 net1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11677__B net1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10581__B net1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11163_ _06124_ _06125_ _06133_ _06134_ vssd1 vssd1 vccd1 vccd1 _06136_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_8_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10114_ _05072_ _05085_ _05086_ _05076_ vssd1 vssd1 vccd1 vccd1 _05087_ sky130_fd_sc_hd__or4b_2
XTAP_TAPCELL_ROW_8_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13892__B net52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15971_ ag2.body\[142\] net212 _01658_ ag2.body\[134\] vssd1 vssd1 vccd1 vccd1 _01200_
+ sky130_fd_sc_hd__a22o_1
X_11094_ ag2.body\[424\] net1224 vssd1 vssd1 vccd1 vccd1 _06067_ sky130_fd_sc_hd__xnor2_1
XANTENNA__14683__A1 net808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17710_ net396 _03388_ _03387_ net362 vssd1 vssd1 vccd1 vccd1 _03389_ sky130_fd_sc_hd__a211o_1
XANTENNA__14683__B2 net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10045_ net1157 control.body\[899\] vssd1 vssd1 vccd1 vccd1 _05018_ sky130_fd_sc_hd__xor2_1
X_14922_ control.body\[1064\] net170 _01543_ net2195 vssd1 vssd1 vccd1 vccd1 _00266_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_69_2418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18690_ clknet_leaf_28_clk img_gen.tracker.next_frame\[128\] net1337 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[128\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_69_2429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold60 img_gen.tracker.frame\[449\] vssd1 vssd1 vccd1 vccd1 net1622 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_117_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19929__CLK clknet_leaf_51_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold71 img_gen.tracker.frame\[514\] vssd1 vssd1 vccd1 vccd1 net1633 sky130_fd_sc_hd__dlygate4sd3_1
X_17641_ ag2.body\[160\] net738 net697 ag2.body\[166\] vssd1 vssd1 vccd1 vccd1 _03320_
+ sky130_fd_sc_hd__a22o_1
Xhold82 img_gen.tracker.frame\[510\] vssd1 vssd1 vccd1 vccd1 net1644 sky130_fd_sc_hd__dlygate4sd3_1
X_14853_ _08836_ _08842_ _01523_ _08574_ vssd1 vssd1 vccd1 vccd1 _01524_ sky130_fd_sc_hd__o211a_1
Xhold93 img_gen.tracker.frame\[528\] vssd1 vssd1 vccd1 vccd1 net1655 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_1278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13804_ net777 _06505_ _06557_ net1167 _06560_ vssd1 vssd1 vccd1 vccd1 _08106_ sky130_fd_sc_hd__o221a_1
XANTENNA__15452__X _01602_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17572_ _03245_ _03246_ _03249_ _03250_ vssd1 vssd1 vccd1 vccd1 _03251_ sky130_fd_sc_hd__or4_2
XANTENNA__10102__A net638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14784_ _01451_ _01452_ _01448_ _01450_ vssd1 vssd1 vccd1 vccd1 _01455_ sky130_fd_sc_hd__a211o_1
XFILLER_0_98_684 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11996_ img_gen.tracker.frame\[421\] net617 net583 img_gen.tracker.frame\[430\] _06967_
+ vssd1 vssd1 vccd1 vccd1 _06968_ sky130_fd_sc_hd__o221a_1
XFILLER_0_97_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19311_ clknet_leaf_99_clk _00255_ net1445 vssd1 vssd1 vccd1 vccd1 control.body\[1085\]
+ sky130_fd_sc_hd__dfrtp_1
X_16523_ _02139_ _02170_ _02201_ vssd1 vssd1 vccd1 vccd1 _02202_ sky130_fd_sc_hd__and3b_1
XFILLER_0_133_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13735_ _04391_ _07243_ _08056_ _07229_ vssd1 vssd1 vccd1 vccd1 _00056_ sky130_fd_sc_hd__a22o_1
X_10947_ _05074_ _05238_ vssd1 vssd1 vccd1 vccd1 _05920_ sky130_fd_sc_hd__nor2_1
XFILLER_0_58_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18953__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19242_ clknet_leaf_76_clk _00186_ net1481 vssd1 vssd1 vccd1 vccd1 ag2.body\[105\]
+ sky130_fd_sc_hd__dfrtp_4
X_16454_ _02129_ _02131_ _02132_ net365 vssd1 vssd1 vccd1 vccd1 _02133_ sky130_fd_sc_hd__a22o_1
X_13666_ net998 net989 net818 _08016_ _08013_ vssd1 vssd1 vccd1 vccd1 obsrand1.next_randY\[1\]
+ sky130_fd_sc_hd__o221a_1
XANTENNA__15935__B2 ag2.body\[165\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_1639 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10878_ ag2.body\[533\] net1108 vssd1 vssd1 vccd1 vccd1 _05851_ sky130_fd_sc_hd__xor2_1
XANTENNA__20149__RESET_B net1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14228__B net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15405_ net2356 net80 _01581_ net2378 vssd1 vssd1 vccd1 vccd1 _00696_ sky130_fd_sc_hd__a22o_1
X_19173_ clknet_leaf_21_clk _00117_ net1363 vssd1 vssd1 vccd1 vccd1 ag2.body\[36\]
+ sky130_fd_sc_hd__dfrtp_4
X_12617_ net250 _07509_ _07510_ net2007 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[64\]
+ sky130_fd_sc_hd__a22o_1
X_16385_ _02061_ _02062_ vssd1 vssd1 vccd1 vccd1 _02064_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_22_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13597_ control.divider.count\[15\] _07949_ _07969_ _07970_ _07971_ vssd1 vssd1 vccd1
+ vccd1 _07972_ sky130_fd_sc_hd__o2111a_1
XANTENNA__11957__C1 net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18124_ net352 net38 _03638_ obsg2.obstacleArray\[62\] vssd1 vssd1 vccd1 vccd1 _03698_
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_5_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15336_ _05283_ net52 vssd1 vssd1 vccd1 vccd1 _01590_ sky130_fd_sc_hd__nor2_2
X_12548_ net306 _07472_ vssd1 vssd1 vccd1 vccd1 _07473_ sky130_fd_sc_hd__or2_1
XFILLER_0_124_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18055_ net43 _03652_ vssd1 vssd1 vccd1 vccd1 _03653_ sky130_fd_sc_hd__nor2_1
XANTENNA__11972__A2 net583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15267_ control.body\[762\] net108 _01582_ net2361 vssd1 vssd1 vccd1 vccd1 _00572_
+ sky130_fd_sc_hd__a22o_1
XANTENNA_2 _03230_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12479_ net1654 _07432_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[4\] sky130_fd_sc_hd__and2_1
XANTENNA__14244__A net1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17006_ _04181_ net963 net952 _04182_ _02684_ vssd1 vssd1 vccd1 vccd1 _02685_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_39_1521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14218_ net819 ag2.body\[395\] ag2.body\[396\] net813 vssd1 vssd1 vccd1 vccd1 _08379_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_123_185 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11587__B net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_1559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15198_ net2251 net94 _01573_ control.body\[822\] vssd1 vssd1 vccd1 vccd1 _00512_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__10491__B net1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11185__B1 net782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12921__A1 net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11724__A2 net624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1093 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14149_ net824 ag2.body\[594\] ag2.body\[596\] net811 _08306_ vssd1 vssd1 vccd1 vccd1
+ _08310_ sky130_fd_sc_hd__o221a_1
XFILLER_0_61_1558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17274__B net849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18957_ clknet_leaf_5_clk img_gen.tracker.next_frame\[395\] net1269 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[395\] sky130_fd_sc_hd__dfrtp_1
X_17908_ net352 _03533_ vssd1 vssd1 vccd1 vccd1 _03543_ sky130_fd_sc_hd__nand2_1
XFILLER_0_94_1312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09690_ ag2.body\[68\] net1139 vssd1 vssd1 vccd1 vccd1 _04663_ sky130_fd_sc_hd__nand2_1
X_18888_ clknet_leaf_27_clk img_gen.tracker.next_frame\[326\] net1341 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[326\] sky130_fd_sc_hd__dfrtp_1
Xfanout1080 net1082 vssd1 vssd1 vccd1 vccd1 net1080 sky130_fd_sc_hd__buf_4
Xfanout1091 net1092 vssd1 vssd1 vccd1 vccd1 net1091 sky130_fd_sc_hd__buf_4
X_17839_ ag2.apple_cord\[6\] _03489_ _03496_ net685 vssd1 vssd1 vccd1 vccd1 _01229_
+ sky130_fd_sc_hd__a211o_1
XANTENNA__12211__B net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__20586__CLK clknet_leaf_105_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12437__B1 _06490_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13026__C _07638_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14831__D1 _08268_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09801__A net1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19509_ clknet_leaf_121_clk _00453_ net1403 vssd1 vssd1 vccd1 vccd1 control.body\[883\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__16179__A1 net373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10947__A _05074_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_3304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_1221 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_3315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_3326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_436 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11660__A1 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20501__RESET_B net1362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1066_A net1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09124_ ag2.body\[418\] vssd1 vssd1 vccd1 vccd1 _04149_ sky130_fd_sc_hd__inv_2
XFILLER_0_17_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12881__B _07639_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11963__A2 net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09055_ ag2.body\[249\] vssd1 vssd1 vccd1 vccd1 _04080_ sky130_fd_sc_hd__inv_2
XFILLER_0_60_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1233_A net1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13165__A1 net232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold530 img_gen.tracker.frame\[561\] vssd1 vssd1 vccd1 vccd1 net2092 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout693_A net694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold541 control.body\[772\] vssd1 vssd1 vccd1 vccd1 net2103 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold552 img_gen.tracker.frame\[430\] vssd1 vssd1 vccd1 vccd1 net2114 sky130_fd_sc_hd__dlygate4sd3_1
X_20215_ clknet_leaf_60_clk _01159_ net1466 vssd1 vssd1 vccd1 vccd1 ag2.body\[181\]
+ sky130_fd_sc_hd__dfrtp_4
Xhold563 control.body\[1118\] vssd1 vssd1 vccd1 vccd1 net2125 sky130_fd_sc_hd__dlygate4sd3_1
Xhold574 control.body\[704\] vssd1 vssd1 vccd1 vccd1 net2136 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__17300__B1 net944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1021_X net1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1400_A net1404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10923__B1 net754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold585 img_gen.tracker.frame\[339\] vssd1 vssd1 vccd1 vccd1 net2147 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1119_X net1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18826__CLK clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold596 _00218_ vssd1 vssd1 vccd1 vccd1 net2158 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20146_ clknet_leaf_101_clk _01090_ net1444 vssd1 vssd1 vccd1 vccd1 ag2.body\[240\]
+ sky130_fd_sc_hd__dfrtp_4
X_09957_ _04421_ _04603_ _04572_ vssd1 vssd1 vccd1 vccd1 _04930_ sky130_fd_sc_hd__o21ai_2
XANTENNA__17184__B net859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout860_A net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout481_X net481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout958_A net968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout579_X net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20077_ clknet_leaf_77_clk _01021_ net1491 vssd1 vssd1 vccd1 vccd1 ag2.body\[315\]
+ sky130_fd_sc_hd__dfrtp_4
X_09888_ _04632_ _04860_ vssd1 vssd1 vccd1 vccd1 _04861_ sky130_fd_sc_hd__or2_2
XFILLER_0_77_1554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17912__B _03542_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15614__B1 _01620_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14417__B2 net844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout746_X net746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11850_ net466 _06673_ vssd1 vssd1 vccd1 vccd1 _06822_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_68_813 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12979__A1 net225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10801_ ag2.body\[39\] net1054 vssd1 vssd1 vccd1 vccd1 _05774_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_16_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10857__A net1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11781_ img_gen.tracker.frame\[191\] net587 net548 img_gen.tracker.frame\[188\] _06752_
+ vssd1 vssd1 vccd1 vccd1 _06753_ sky130_fd_sc_hd__o221a_1
XFILLER_0_135_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_0_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13520_ net2129 net655 _07919_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[558\]
+ sky130_fd_sc_hd__and3_1
XANTENNA__09430__B net1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10732_ ag2.body\[254\] net1086 vssd1 vssd1 vccd1 vccd1 _05705_ sky130_fd_sc_hd__and2_1
XANTENNA__10576__B net1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13451_ net682 _07892_ vssd1 vssd1 vccd1 vccd1 _07893_ sky130_fd_sc_hd__nor2_1
X_10663_ net1099 control.body\[885\] vssd1 vssd1 vccd1 vccd1 _05636_ sky130_fd_sc_hd__xor2_1
XANTENNA__20309__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_1601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12402_ _07278_ _07330_ _07348_ _07282_ vssd1 vssd1 vccd1 vccd1 _07366_ sky130_fd_sc_hd__o31a_1
X_16170_ net378 _01848_ _01847_ net347 vssd1 vssd1 vccd1 vccd1 _01849_ sky130_fd_sc_hd__a211o_1
XFILLER_0_49_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10594_ net1100 control.body\[829\] vssd1 vssd1 vccd1 vccd1 _05567_ sky130_fd_sc_hd__xor2_1
XFILLER_0_35_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13382_ _07542_ net304 vssd1 vssd1 vccd1 vccd1 _07866_ sky130_fd_sc_hd__nor2_1
XFILLER_0_36_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15121_ control.body\[889\] net103 _01565_ net2503 vssd1 vssd1 vccd1 vccd1 _00443_
+ sky130_fd_sc_hd__a22o_1
X_12333_ _07294_ _07298_ _07284_ vssd1 vssd1 vccd1 vccd1 _07300_ sky130_fd_sc_hd__o21a_2
XFILLER_0_133_461 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19601__CLK clknet_leaf_118_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10592__A net1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_3_3_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_3_3_0_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__13156__A1 net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15052_ net2630 net164 _01558_ control.body\[947\] vssd1 vssd1 vccd1 vccd1 _00381_
+ sky130_fd_sc_hd__a22o_1
X_12264_ _07191_ _07233_ vssd1 vssd1 vccd1 vccd1 _07234_ sky130_fd_sc_hd__or2_1
XFILLER_0_120_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14003_ net1031 ag2.body\[509\] vssd1 vssd1 vccd1 vccd1 _08164_ sky130_fd_sc_hd__xor2_1
XFILLER_0_43_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11706__A2 net606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11215_ net1076 control.body\[846\] vssd1 vssd1 vccd1 vccd1 _06188_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_31_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12195_ _07155_ _07156_ _07159_ _07160_ vssd1 vssd1 vccd1 vccd1 _07167_ sky130_fd_sc_hd__a22o_1
X_19860_ clknet_leaf_94_clk _00804_ net1436 vssd1 vssd1 vccd1 vccd1 ag2.body\[530\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_120_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_881 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18811_ clknet_leaf_3_clk img_gen.tracker.next_frame\[249\] net1259 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[249\] sky130_fd_sc_hd__dfrtp_1
X_11146_ ag2.body\[411\] net768 net749 ag2.body\[414\] _06114_ vssd1 vssd1 vccd1 vccd1
+ _06119_ sky130_fd_sc_hd__a221o_1
XFILLER_0_128_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19791_ clknet_leaf_128_clk _00735_ net1329 vssd1 vssd1 vccd1 vccd1 ag2.body\[605\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__14656__A1 net839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14656__B2 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15954_ ag2.body\[159\] net199 _01656_ ag2.body\[151\] vssd1 vssd1 vccd1 vccd1 _01185_
+ sky130_fd_sc_hd__a22o_1
X_11077_ _06045_ _06046_ _06048_ _06049_ vssd1 vssd1 vccd1 vccd1 _06050_ sky130_fd_sc_hd__and4_1
XFILLER_0_95_1610 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18742_ clknet_leaf_143_clk img_gen.tracker.next_frame\[180\] net1256 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[180\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_120_1489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10355__A_N ag2.body\[290\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12131__A2 net588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10028_ _04999_ _05000_ _04998_ vssd1 vssd1 vccd1 vccd1 _05001_ sky130_fd_sc_hd__a21o_1
X_14905_ control.body\[1081\] net177 _01541_ control.body\[1073\] vssd1 vssd1 vccd1
+ vccd1 _00251_ sky130_fd_sc_hd__a22o_1
X_18673_ clknet_leaf_27_clk img_gen.tracker.next_frame\[111\] net1340 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[111\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__13127__B _07587_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14408__A1 net998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15885_ ag2.body\[209\] net184 _01649_ ag2.body\[201\] vssd1 vssd1 vccd1 vccd1 _01123_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_91_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15605__B1 _01619_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_1638 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15623__A _06314_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17624_ ag2.body\[185\] net872 vssd1 vssd1 vccd1 vccd1 _03303_ sky130_fd_sc_hd__xor2_1
XANTENNA__17070__A2 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14836_ _08585_ _08587_ _08593_ _08884_ _08467_ vssd1 vssd1 vccd1 vccd1 _01507_ sky130_fd_sc_hd__o311a_1
XANTENNA__11890__A1 net576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_1447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17555_ _04126_ net865 net693 ag2.body\[359\] _03233_ vssd1 vssd1 vccd1 vccd1 _03234_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_59_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14767_ net1001 ag2.body\[96\] vssd1 vssd1 vccd1 vccd1 _08928_ sky130_fd_sc_hd__xor2_1
X_11979_ _06947_ _06948_ _06950_ net564 vssd1 vssd1 vccd1 vccd1 _06951_ sky130_fd_sc_hd__a22o_1
XFILLER_0_58_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16506_ obsg2.obstacleArray\[8\] obsg2.obstacleArray\[9\] net456 vssd1 vssd1 vccd1
+ vccd1 _02185_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_1335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11642__A1 net505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13718_ track.nextHighScore\[6\] vssd1 vssd1 vccd1 vccd1 _08052_ sky130_fd_sc_hd__inv_2
XFILLER_0_128_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17486_ _04129_ net888 net728 ag2.body\[362\] vssd1 vssd1 vccd1 vccd1 _03165_ sky130_fd_sc_hd__a22o_1
X_14698_ net1023 ag2.body\[326\] vssd1 vssd1 vccd1 vccd1 _08859_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_6_1171 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_849 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16437_ net399 _02115_ vssd1 vssd1 vccd1 vccd1 _02116_ sky130_fd_sc_hd__or2_1
X_19225_ clknet_leaf_75_clk _00169_ net1483 vssd1 vssd1 vccd1 vccd1 ag2.body\[88\]
+ sky130_fd_sc_hd__dfrtp_4
X_13649_ control.divider.count\[17\] _08005_ net221 vssd1 vssd1 vccd1 vccd1 _08007_
+ sky130_fd_sc_hd__o21ai_1
XANTENNA__16581__A1 net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13395__A1 net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19156_ clknet_leaf_50_clk _00100_ net1367 vssd1 vssd1 vccd1 vccd1 ag2.body\[20\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_125_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16368_ _01896_ _01918_ _01929_ vssd1 vssd1 vccd1 vccd1 _02047_ sky130_fd_sc_hd__and3_1
XFILLER_0_125_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19538__Q control.body\[848\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18107_ net353 _03621_ vssd1 vssd1 vccd1 vccd1 _03687_ sky130_fd_sc_hd__nand2_1
X_15319_ _05036_ net63 vssd1 vssd1 vccd1 vccd1 _01589_ sky130_fd_sc_hd__and2_2
XFILLER_0_28_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11945__A2 net618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16333__A1 net371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15136__A2 net107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19087_ clknet_leaf_9_clk img_gen.tracker.next_frame\[525\] net1271 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[525\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_129_1470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16299_ net371 _01973_ net368 vssd1 vssd1 vccd1 vccd1 _01978_ sky130_fd_sc_hd__o21a_1
Xclkbuf_leaf_120_clk clknet_4_8__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_120_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_41_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13147__A1 net231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18849__CLK clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18038_ _03543_ net42 vssd1 vssd1 vccd1 vccd1 _03642_ sky130_fd_sc_hd__nor2_1
XFILLER_0_112_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16884__A2 net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14702__A net1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20000_ clknet_leaf_58_clk _00944_ net1472 vssd1 vssd1 vccd1 vccd1 ag2.body\[398\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__16097__B1 _01729_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout306 net307 vssd1 vssd1 vccd1 vccd1 net306 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_26_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09811_ net1181 control.body\[1050\] vssd1 vssd1 vccd1 vccd1 _04784_ sky130_fd_sc_hd__xor2_1
Xfanout328 net331 vssd1 vssd1 vccd1 vccd1 net328 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_10_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout339 net340 vssd1 vssd1 vccd1 vccd1 net339 sky130_fd_sc_hd__buf_4
X_19989_ clknet_leaf_64_clk _00933_ net1475 vssd1 vssd1 vccd1 vccd1 ag2.body\[403\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA_clkload11_A clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15844__B1 _01644_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17572__X _03251_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09742_ ag2.body\[355\] net1163 vssd1 vssd1 vccd1 vccd1 _04715_ sky130_fd_sc_hd__xor2_1
XFILLER_0_94_53 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10373__B_N net920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_97 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13037__B _07542_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09673_ net923 _04634_ vssd1 vssd1 vccd1 vccd1 _04646_ sky130_fd_sc_hd__or2_4
XANTENNA__11483__D _06455_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10013__Y _04986_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout274_A net279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1441 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17061__A2 net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1017 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10684__A2 _04695_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10948__Y _05921_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12876__B net311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09531__A net1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout441_A net443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1183_A net1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13053__A net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1350_A net1351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12892__A net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout706_A net708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1069_X net1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1448_A net1452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11397__B1 _06369_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09107_ ag2.body\[370\] vssd1 vssd1 vccd1 vccd1 _04132_ sky130_fd_sc_hd__inv_2
XANTENNA__11936__A2 net621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17747__X _03426_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13500__B net304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_111_clk clknet_4_10__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_111_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_32_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1236_X net1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16875__A2 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09038_ ag2.body\[201\] vssd1 vssd1 vccd1 vccd1 _04063_ sky130_fd_sc_hd__inv_2
XFILLER_0_103_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17907__B net485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout696_X net696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13689__A2 net434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11020__B net1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold360 img_gen.tracker.frame\[159\] vssd1 vssd1 vccd1 vccd1 net1922 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16303__S net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1403_X net1403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold371 img_gen.tracker.frame\[270\] vssd1 vssd1 vccd1 vccd1 net1933 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold382 img_gen.tracker.frame\[82\] vssd1 vssd1 vccd1 vccd1 net1944 sky130_fd_sc_hd__dlygate4sd3_1
X_11000_ _05253_ _05964_ _05967_ _05972_ vssd1 vssd1 vccd1 vccd1 _05973_ sky130_fd_sc_hd__or4_4
XFILLER_0_99_1020 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold393 img_gen.tracker.frame\[131\] vssd1 vssd1 vccd1 vccd1 net1955 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout863_X net863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10372__A1 net767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14638__A1 net840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14638__B2 net832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout840 net847 vssd1 vssd1 vccd1 vccd1 net840 sky130_fd_sc_hd__clkbuf_4
Xfanout851 net852 vssd1 vssd1 vccd1 vccd1 net851 sky130_fd_sc_hd__buf_2
XFILLER_0_79_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20129_ clknet_leaf_81_clk _01073_ net1485 vssd1 vssd1 vccd1 vccd1 ag2.body\[271\]
+ sky130_fd_sc_hd__dfrtp_4
Xfanout862 net867 vssd1 vssd1 vccd1 vccd1 net862 sky130_fd_sc_hd__buf_4
XANTENNA__10204__X _05177_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout873 net875 vssd1 vssd1 vccd1 vccd1 net873 sky130_fd_sc_hd__clkbuf_4
Xfanout884 net889 vssd1 vssd1 vccd1 vccd1 net884 sky130_fd_sc_hd__clkbuf_8
XANTENNA__12113__A2 net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout895 control.body_update.curr_length\[7\] vssd1 vssd1 vccd1 vccd1 net895 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12489__D _07312_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12951_ net293 _07670_ _07671_ net1604 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[236\]
+ sky130_fd_sc_hd__a22o_1
Xhold1060 control.body\[914\] vssd1 vssd1 vccd1 vccd1 net2622 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11321__B1 net1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1071 control.body\[878\] vssd1 vssd1 vccd1 vccd1 net2633 sky130_fd_sc_hd__dlygate4sd3_1
X_11902_ _06870_ _06873_ net471 vssd1 vssd1 vccd1 vccd1 _06874_ sky130_fd_sc_hd__a21o_1
X_15670_ ag2.body\[401\] net195 _01626_ ag2.body\[393\] vssd1 vssd1 vccd1 vccd1 _00931_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_119_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold1082 control.body\[729\] vssd1 vssd1 vccd1 vccd1 net2644 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11872__A1 net563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1093 control.body\[873\] vssd1 vssd1 vccd1 vccd1 net2655 sky130_fd_sc_hd__dlygate4sd3_1
X_12882_ net680 _07641_ vssd1 vssd1 vccd1 vccd1 _07642_ sky130_fd_sc_hd__nor2_1
X_14621_ _08776_ _08777_ _08781_ vssd1 vssd1 vccd1 vccd1 _08782_ sky130_fd_sc_hd__and3_1
XANTENNA__11690__B net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11833_ img_gen.tracker.frame\[539\] net579 net541 img_gen.tracker.frame\[536\] _06804_
+ vssd1 vssd1 vccd1 vccd1 _06805_ sky130_fd_sc_hd__o221a_1
XANTENNA__10587__A net1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09817__A1 net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14810__A1 net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09817__B2 net755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14810__B2 net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17340_ net927 net709 vssd1 vssd1 vccd1 vccd1 _03019_ sky130_fd_sc_hd__nand2_1
XFILLER_0_95_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14552_ net1040 ag2.body\[68\] vssd1 vssd1 vccd1 vccd1 _08713_ sky130_fd_sc_hd__xor2_1
XFILLER_0_90_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11764_ net1215 net1190 img_gen.tracker.frame\[62\] vssd1 vssd1 vccd1 vccd1 _06736_
+ sky130_fd_sc_hd__or3_1
XFILLER_0_16_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13503_ net250 _07912_ _07913_ net1886 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[547\]
+ sky130_fd_sc_hd__a22o_1
X_10715_ ag2.body\[619\] net1152 vssd1 vssd1 vccd1 vccd1 _05688_ sky130_fd_sc_hd__xor2_1
X_17271_ _02944_ _02949_ vssd1 vssd1 vccd1 vccd1 _02950_ sky130_fd_sc_hd__nand2b_1
X_14483_ _08636_ _08637_ _08638_ _08640_ vssd1 vssd1 vccd1 vccd1 _08644_ sky130_fd_sc_hd__or4_1
X_11695_ _06662_ _06664_ _06666_ net572 net473 vssd1 vssd1 vccd1 vccd1 _06667_ sky130_fd_sc_hd__a221o_1
XFILLER_0_138_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19010_ clknet_leaf_1_clk img_gen.tracker.next_frame\[448\] net1244 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[448\] sky130_fd_sc_hd__dfrtp_1
X_16222_ _01725_ _01888_ _01900_ vssd1 vssd1 vccd1 vccd1 _01901_ sky130_fd_sc_hd__o21a_1
XANTENNA__11689__Y _06661_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13434_ net281 _07884_ _07885_ net1947 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[506\]
+ sky130_fd_sc_hd__a22o_1
X_10646_ _05529_ _05558_ _05587_ _05618_ vssd1 vssd1 vccd1 vccd1 _05619_ sky130_fd_sc_hd__nand4_1
XFILLER_0_107_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16153_ obsg2.obstacleArray\[5\] net431 vssd1 vssd1 vccd1 vccd1 _01832_ sky130_fd_sc_hd__or2_1
XFILLER_0_84_1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16315__A1 net415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_102_clk clknet_4_10__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_102_clk
+ sky130_fd_sc_hd__clkbuf_8
X_13365_ net249 _07858_ _07859_ net1830 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[463\]
+ sky130_fd_sc_hd__a22o_1
X_10577_ ag2.body\[186\] net1177 vssd1 vssd1 vccd1 vccd1 _05550_ sky130_fd_sc_hd__nand2_1
XFILLER_0_126_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10060__B1 net1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11211__A net1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15104_ net2093 net145 _01564_ control.body\[897\] vssd1 vssd1 vccd1 vccd1 _00427_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_11_407 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12316_ _07264_ _07273_ _07271_ vssd1 vssd1 vccd1 vccd1 _07283_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_23_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16084_ net373 _01760_ _01762_ net346 vssd1 vssd1 vccd1 vccd1 _01763_ sky130_fd_sc_hd__a211o_1
X_13296_ net255 _07831_ _07832_ net1738 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[421\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_126_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19912_ clknet_leaf_54_clk _00856_ net1457 vssd1 vssd1 vccd1 vccd1 ag2.body\[486\]
+ sky130_fd_sc_hd__dfrtp_4
X_15035_ control.body\[971\] net165 _01557_ net2436 vssd1 vssd1 vccd1 vccd1 _00365_
+ sky130_fd_sc_hd__a22o_1
X_12247_ _07203_ _07214_ _07216_ _07209_ vssd1 vssd1 vccd1 vccd1 _07217_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_20_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09616__A net1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19843_ clknet_leaf_92_clk _00787_ net1412 vssd1 vssd1 vccd1 vccd1 ag2.body\[545\]
+ sky130_fd_sc_hd__dfrtp_4
X_12178_ net480 _07147_ vssd1 vssd1 vccd1 vccd1 _07150_ sky130_fd_sc_hd__nand2_1
XANTENNA__10363__A1 net773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15826__B1 _01643_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10363__B2 net753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17833__A net662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11129_ _06098_ _06099_ _06100_ _06101_ vssd1 vssd1 vccd1 vccd1 _06102_ sky130_fd_sc_hd__or4_1
XFILLER_0_3_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10114__X _05087_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19774_ clknet_leaf_19_clk _00718_ net1331 vssd1 vssd1 vccd1 vccd1 ag2.body\[620\]
+ sky130_fd_sc_hd__dfrtp_4
X_16986_ _04021_ net942 net692 ag2.body\[95\] vssd1 vssd1 vccd1 vccd1 _02665_ sky130_fd_sc_hd__a22o_1
XANTENNA__12104__A2 net628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13301__A1 net256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09903__X _04876_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18725_ clknet_leaf_142_clk img_gen.tracker.next_frame\[163\] net1257 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[163\] sky130_fd_sc_hd__dfrtp_1
X_15937_ ag2.body\[175\] net126 _01655_ ag2.body\[167\] vssd1 vssd1 vccd1 vccd1 _01169_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__17552__B net888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18656_ clknet_leaf_130_clk img_gen.tracker.next_frame\[94\] net1317 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[94\] sky130_fd_sc_hd__dfrtp_1
X_15868_ ag2.body\[226\] net160 _01647_ ag2.body\[218\] vssd1 vssd1 vccd1 vccd1 _01108_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_133_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14819_ net845 ag2.body\[152\] ag2.body\[155\] net822 vssd1 vssd1 vccd1 vccd1 _01490_
+ sky130_fd_sc_hd__o22a_1
X_17607_ _03277_ _03280_ _03281_ _03285_ vssd1 vssd1 vccd1 vccd1 _03286_ sky130_fd_sc_hd__or4_4
X_15799_ ag2.body\[292\] net205 _01640_ ag2.body\[284\] vssd1 vssd1 vccd1 vccd1 _01046_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__09808__A1 _04551_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18587_ clknet_leaf_14_clk img_gen.tracker.next_frame\[25\] net1280 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[25\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_114_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11615__A1 net508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17538_ ag2.body\[278\] net699 net936 _04095_ _03216_ vssd1 vssd1 vccd1 vccd1 _03217_
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_50_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_715 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17469_ _04193_ net874 net700 ag2.body\[534\] vssd1 vssd1 vccd1 vccd1 _03148_ sky130_fd_sc_hd__o22a_1
XFILLER_0_131_1382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17751__B1 _03333_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19208_ clknet_leaf_86_clk _00152_ net1459 vssd1 vssd1 vccd1 vccd1 ag2.body\[71\]
+ sky130_fd_sc_hd__dfrtp_4
X_20480_ clknet_leaf_39_clk _01367_ net1355 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[116\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__11379__B1 net1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_1531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11918__A2 net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19139_ clknet_leaf_132_clk img_gen.control.next\[1\] net1303 vssd1 vssd1 vccd1 vccd1
+ img_gen.control.current\[1\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_15_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17503__B1 net726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11121__A net1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12591__A2 net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_114_3790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_965 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_110_3665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_3676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_110_3687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1029_A ag2.randCord\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout103 net104 vssd1 vssd1 vccd1 vccd1 net103 sky130_fd_sc_hd__buf_2
XANTENNA__09526__A net1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout114 net219 vssd1 vssd1 vccd1 vccd1 net114 sky130_fd_sc_hd__buf_2
Xfanout125 net127 vssd1 vssd1 vccd1 vccd1 net125 sky130_fd_sc_hd__buf_2
XANTENNA_fanout391_A net393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout136 net139 vssd1 vssd1 vccd1 vccd1 net136 sky130_fd_sc_hd__clkbuf_4
Xfanout147 net154 vssd1 vssd1 vccd1 vccd1 net147 sky130_fd_sc_hd__buf_2
XFILLER_0_129_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout158 net161 vssd1 vssd1 vccd1 vccd1 net158 sky130_fd_sc_hd__buf_2
XANTENNA__13048__A net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19177__CLK clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13828__C1 _08113_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout169 net171 vssd1 vssd1 vccd1 vccd1 net169 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_138_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09725_ _04695_ net634 vssd1 vssd1 vccd1 vccd1 _04698_ sky130_fd_sc_hd__or2_1
XANTENNA__17462__B net853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12887__A net678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout277_X net277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout656_A net657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1569 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15263__A _04573_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16468__S1 net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09656_ _04619_ _04620_ _04622_ _04623_ vssd1 vssd1 vccd1 vccd1 _04629_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_2_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout823_A _03968_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16793__A1 net399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09587_ net1227 control.body\[904\] vssd1 vssd1 vccd1 vccd1 _04560_ sky130_fd_sc_hd__or2_1
XFILLER_0_136_1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17990__B1 net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1186_X net1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16806__B net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11015__B net1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout611_X net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout709_X net709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10500_ _05453_ _05457_ _05462_ _05472_ _05302_ vssd1 vssd1 vccd1 vccd1 _05473_ sky130_fd_sc_hd__a32o_1
XFILLER_0_68_1317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_1466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11480_ ag2.body\[492\] net1138 vssd1 vssd1 vccd1 vccd1 _06453_ sky130_fd_sc_hd__xor2_1
XFILLER_0_68_1339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11909__A2 net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10431_ net786 control.body\[1064\] _05402_ _05403_ net742 vssd1 vssd1 vccd1 vccd1
+ _05404_ sky130_fd_sc_hd__a221o_1
XFILLER_0_116_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09578__A3 net908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_420 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11031__A net1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13150_ net277 _07764_ _07765_ net1892 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[341\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_21_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout980_X net980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10362_ _05305_ _05312_ _05319_ _05323_ _05334_ vssd1 vssd1 vccd1 vccd1 _05335_ sky130_fd_sc_hd__o32a_2
X_12101_ img_gen.tracker.frame\[375\] net610 net555 img_gen.tracker.frame\[378\] _07072_
+ vssd1 vssd1 vccd1 vccd1 _07073_ sky130_fd_sc_hd__a221o_1
X_10293_ ag2.body\[331\] net1165 vssd1 vssd1 vccd1 vccd1 _05266_ sky130_fd_sc_hd__xor2_1
XFILLER_0_108_1384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10870__A ag2.body\[534\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13081_ net291 _07731_ _07732_ net1858 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[305\]
+ sky130_fd_sc_hd__a22o_1
XANTENNA__14342__A net979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12334__A2 _06985_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09735__B1 net1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12032_ img_gen.tracker.frame\[30\] net556 _07003_ vssd1 vssd1 vccd1 vccd1 _07004_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_104_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold190 img_gen.tracker.frame\[530\] vssd1 vssd1 vccd1 vccd1 net1752 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121_1540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15808__B1 _01641_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16840_ _02512_ _02514_ _02517_ _02518_ vssd1 vssd1 vccd1 vccd1 _02519_ sky130_fd_sc_hd__nand4_1
XFILLER_0_121_1595 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout670 net672 vssd1 vssd1 vccd1 vccd1 net670 sky130_fd_sc_hd__clkbuf_4
Xfanout681 _04393_ vssd1 vssd1 vccd1 vccd1 net681 sky130_fd_sc_hd__buf_2
XANTENNA__17372__B net926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16771_ obsg2.obstacleArray\[15\] net501 net487 obsg2.obstacleArray\[14\] vssd1 vssd1
+ vccd1 vccd1 _02450_ sky130_fd_sc_hd__a22o_1
Xfanout692 net695 vssd1 vssd1 vccd1 vccd1 net692 sky130_fd_sc_hd__buf_4
X_13983_ ag2.body\[120\] net211 _08159_ ag2.body\[112\] vssd1 vssd1 vccd1 vccd1 _00201_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_57_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12797__A net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13834__A2 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15722_ _04719_ _01631_ vssd1 vssd1 vccd1 vccd1 _01632_ sky130_fd_sc_hd__and2b_2
XFILLER_0_73_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18510_ net1513 net1507 vssd1 vssd1 vccd1 vccd1 _00041_ sky130_fd_sc_hd__or2_1
XFILLER_0_92_1635 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12934_ net290 _07662_ _07663_ net1813 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[227\]
+ sky130_fd_sc_hd__a22o_1
X_19490_ clknet_leaf_113_clk _00434_ net1399 vssd1 vssd1 vccd1 vccd1 control.body\[896\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_16_Right_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09171__A ag2.body\[534\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15653_ ag2.body\[418\] net139 _01624_ ag2.body\[410\] vssd1 vssd1 vccd1 vccd1 _00916_
+ sky130_fd_sc_hd__a22o_1
X_18441_ track.nextHighScore\[7\] _03913_ _03785_ vssd1 vssd1 vccd1 vccd1 _03930_
+ sky130_fd_sc_hd__a21o_1
X_12865_ net383 net309 _07633_ vssd1 vssd1 vccd1 vccd1 _07634_ sky130_fd_sc_hd__and3_1
XANTENNA__16784__A1 net462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17981__B1 net523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11519__A_N net1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14604_ net1012 ag2.body\[135\] vssd1 vssd1 vccd1 vccd1 _08765_ sky130_fd_sc_hd__nand2_1
XFILLER_0_29_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18372_ net1951 _03864_ _08024_ vssd1 vssd1 vccd1 vccd1 _01394_ sky130_fd_sc_hd__mux2_1
X_11816_ img_gen.tracker.frame\[407\] net584 vssd1 vssd1 vccd1 vccd1 _06788_ sky130_fd_sc_hd__or2_1
XANTENNA__15901__A _05543_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15584_ ag2.body\[484\] net130 _01617_ ag2.body\[476\] vssd1 vssd1 vccd1 vccd1 _00854_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__10110__A net1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12796_ _07423_ _07501_ net308 net341 vssd1 vssd1 vccd1 vccd1 _07601_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_95_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17323_ _02995_ _02997_ _03000_ _03001_ vssd1 vssd1 vccd1 vccd1 _03002_ sky130_fd_sc_hd__or4_1
XFILLER_0_16_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14535_ net1030 _04083_ ag2.body\[254\] net804 vssd1 vssd1 vccd1 vccd1 _08696_ sky130_fd_sc_hd__a22o_1
XFILLER_0_83_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11747_ _06690_ _06717_ _06718_ _06705_ net387 vssd1 vssd1 vccd1 vccd1 _06719_ sky130_fd_sc_hd__a311o_1
XFILLER_0_126_512 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17733__B1 _03411_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_137_4491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14517__A net1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13421__A net682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17254_ ag2.body\[547\] net716 net689 ag2.body\[551\] vssd1 vssd1 vccd1 vccd1 _02933_
+ sky130_fd_sc_hd__a22o_1
X_14466_ net838 ag2.body\[265\] ag2.body\[267\] net820 vssd1 vssd1 vccd1 vccd1 _08627_
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_55_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_133_4366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_1439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11678_ net1174 net1123 vssd1 vssd1 vccd1 vccd1 _06650_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_133_4377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10764__B net1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16205_ _01743_ _01883_ _01878_ _01728_ vssd1 vssd1 vccd1 vccd1 _01884_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_133_4388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13140__B _07639_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13417_ net236 _07878_ _07879_ net1778 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[495\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_70_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10629_ net1045 control.body\[671\] vssd1 vssd1 vccd1 vccd1 _05602_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_42_1594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17185_ ag2.body\[569\] net869 vssd1 vssd1 vccd1 vccd1 _02864_ sky130_fd_sc_hd__xor2_1
X_14397_ net821 ag2.body\[123\] ag2.body\[126\] net803 vssd1 vssd1 vccd1 vccd1 _08558_
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_109_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_25_Right_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16136_ net882 net870 net860 vssd1 vssd1 vccd1 vccd1 _01815_ sky130_fd_sc_hd__a21o_1
XANTENNA__16839__A2 net735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13348_ net664 _07852_ vssd1 vssd1 vccd1 vccd1 _07853_ sky130_fd_sc_hd__nor2_1
XFILLER_0_51_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17547__B net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11781__B1 net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16067_ obsg2.obstacleArray\[106\] obsg2.obstacleArray\[107\] net421 vssd1 vssd1
+ vccd1 vccd1 _01746_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_1315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10780__A net1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13279_ net671 _07825_ vssd1 vssd1 vccd1 vccd1 _07826_ sky130_fd_sc_hd__nor2_1
XFILLER_0_27_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_968 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09726__B1 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15018_ control.body\[990\] net169 _01553_ control.body\[982\] vssd1 vssd1 vccd1
+ vccd1 _00352_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_55_1988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19826_ clknet_leaf_124_clk _00770_ net1407 vssd1 vssd1 vccd1 vccd1 ag2.body\[560\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__17264__A2 net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1489 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_1072 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__20345__RESET_B net1293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16472__B1 _02075_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09633__X _04606_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15354__Y _01592_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19757_ clknet_leaf_129_clk _00701_ net1326 vssd1 vssd1 vccd1 vccd1 control.body\[635\]
+ sky130_fd_sc_hd__dfrtp_1
X_16969_ ag2.body\[410\] net724 net709 ag2.body\[412\] vssd1 vssd1 vccd1 vccd1 _02648_
+ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_34_Right_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09510_ ag2.body\[401\] net781 net1113 _04145_ _04475_ vssd1 vssd1 vccd1 vccd1 _04483_
+ sky130_fd_sc_hd__a221o_1
X_18708_ clknet_leaf_144_clk img_gen.tracker.next_frame\[146\] net1255 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[146\] sky130_fd_sc_hd__dfrtp_1
X_19688_ clknet_leaf_136_clk net2266 net1302 vssd1 vssd1 vccd1 vccd1 control.body\[710\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12500__A _07443_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10939__B net1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09441_ _04407_ _04408_ _04409_ _04412_ vssd1 vssd1 vccd1 vccd1 _04414_ sky130_fd_sc_hd__or4_1
X_18639_ clknet_leaf_131_clk img_gen.tracker.next_frame\[77\] net1311 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[77\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_52_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16373__A_N net956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14632__A1_N net798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09372_ _04368_ _04371_ vssd1 vssd1 vccd1 vccd1 _01418_ sky130_fd_sc_hd__nor2_1
XFILLER_0_34_1541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20601_ net1533 vssd1 vssd1 vccd1 vccd1 gpio_oeb[13] sky130_fd_sc_hd__buf_2
XFILLER_0_75_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16118__S net377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkload125_A clknet_leaf_83_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14427__A net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout237_A net238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20532_ clknet_leaf_114_clk _01397_ net1398 vssd1 vssd1 vccd1 vccd1 toggle1.bcd_ones\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10674__B net1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_43_Right_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_116_3852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_116_3863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20463_ clknet_leaf_28_clk _01350_ net1337 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[99\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_7_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12013__A1 net385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_116_3874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_112_3727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1146_A net1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_3738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10024__B1 _04986_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_1248 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_112_3749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09808__X _04781_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20394_ clknet_leaf_38_clk _01281_ net1354 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[30\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_63_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16361__B net409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11772__B1 net608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__15502__A2 net113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13513__A1 net288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__09717__B1 net1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout394_X net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout773_A net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_2480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_2491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1101_X net1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_52_Right_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17192__B net929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout940_A net941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout561_X net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13065__X _07726_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13506__A net664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09708_ _04075_ net1232 net779 ag2.body\[241\] _04680_ vssd1 vssd1 vccd1 vccd1 _04681_
+ sky130_fd_sc_hd__a221o_1
XANTENNA__09703__B net1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11827__A1 net571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10980_ net1150 control.body\[755\] vssd1 vssd1 vccd1 vccd1 _05953_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout52_A net55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10849__B net1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09639_ net1206 _04251_ control.body\[1020\] net761 vssd1 vssd1 vccd1 vccd1 _04612_
+ sky130_fd_sc_hd__o22a_1
XANTENNA_fanout1470_X net1470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16766__A1 obsg2.obstacleArray\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_2874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout826_X net826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_2885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15721__A _04418_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_2896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12650_ net678 _07529_ vssd1 vssd1 vccd1 vccd1 _07530_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_80_2749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_65_2295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11601_ _06572_ _06573_ net507 vssd1 vssd1 vccd1 vccd1 _06574_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11055__A2 _04758_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16518__A1 net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12581_ net307 _07490_ vssd1 vssd1 vccd1 vccd1 _07491_ sky130_fd_sc_hd__nor2_1
XFILLER_0_33_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_61_Right_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14320_ net1008 ag2.body\[455\] vssd1 vssd1 vccd1 vccd1 _08481_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_93_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11532_ net1222 net1174 vssd1 vssd1 vccd1 vccd1 _06505_ sky130_fd_sc_hd__nand2_2
XFILLER_0_68_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12004__A1 net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14251_ _08404_ _08405_ _08406_ _08409_ vssd1 vssd1 vccd1 vccd1 _08412_ sky130_fd_sc_hd__or4_1
X_11463_ _04085_ net1237 net1164 _04088_ vssd1 vssd1 vccd1 vccd1 _06436_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_22_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_2689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13202_ net383 _07621_ vssd1 vssd1 vccd1 vccd1 _07791_ sky130_fd_sc_hd__nor2_1
Xwire389 _03164_ vssd1 vssd1 vccd1 vccd1 net389 sky130_fd_sc_hd__buf_1
XFILLER_0_104_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10414_ _05364_ _05368_ _05374_ _05386_ vssd1 vssd1 vccd1 vccd1 _05387_ sky130_fd_sc_hd__o31a_2
XFILLER_0_61_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19269__RESET_B net1503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14182_ net811 ag2.body\[196\] vssd1 vssd1 vccd1 vccd1 _08343_ sky130_fd_sc_hd__nor2_1
X_11394_ net1047 control.body\[647\] vssd1 vssd1 vccd1 vccd1 _06367_ sky130_fd_sc_hd__xor2_1
XFILLER_0_81_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17935__X _03566_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13133_ _07486_ net329 net340 vssd1 vssd1 vccd1 vccd1 _07758_ sky130_fd_sc_hd__and3b_1
XANTENNA__17494__A2 net713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10345_ _05306_ _05307_ _05317_ vssd1 vssd1 vccd1 vccd1 _05318_ sky130_fd_sc_hd__a21o_1
XFILLER_0_103_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14072__A net984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18990_ clknet_leaf_8_clk img_gen.tracker.next_frame\[428\] net1270 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[428\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_103_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13504__A1 net276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09708__B1 net779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17941_ net48 net296 _03570_ vssd1 vssd1 vccd1 vccd1 _03571_ sky130_fd_sc_hd__and3_1
X_13064_ net293 _07723_ _07724_ net1748 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[296\]
+ sky130_fd_sc_hd__a22o_1
X_10276_ ag2.body\[138\] net1186 vssd1 vssd1 vccd1 vccd1 _05249_ sky130_fd_sc_hd__xor2_1
XFILLER_0_123_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_70_Right_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12015_ _06986_ vssd1 vssd1 vccd1 vccd1 _06987_ sky130_fd_sc_hd__inv_2
Xfanout1410 net1415 vssd1 vssd1 vccd1 vccd1 net1410 sky130_fd_sc_hd__clkbuf_4
Xfanout1421 net1423 vssd1 vssd1 vccd1 vccd1 net1421 sky130_fd_sc_hd__clkbuf_2
XANTENNA__17246__A2 net730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10105__A net1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17872_ _03505_ _03515_ vssd1 vssd1 vccd1 vccd1 _01243_ sky130_fd_sc_hd__and2b_1
Xfanout1432 net1433 vssd1 vssd1 vccd1 vccd1 net1432 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_126_4170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14800__A net1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1443 net1444 vssd1 vssd1 vccd1 vccd1 net1443 sky130_fd_sc_hd__clkbuf_4
Xfanout1454 net1455 vssd1 vssd1 vccd1 vccd1 net1454 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_126_4181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18198__B net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19611_ clknet_leaf_119_clk _00555_ net1391 vssd1 vssd1 vccd1 vccd1 control.body\[777\]
+ sky130_fd_sc_hd__dfrtp_1
X_16823_ ag2.body\[225\] net873 vssd1 vssd1 vccd1 vccd1 _02502_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_50_1841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1465 net1478 vssd1 vssd1 vccd1 vccd1 net1465 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_122_4034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1476 net1477 vssd1 vssd1 vccd1 vccd1 net1476 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_79_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10599__X _05572_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_4045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1487 net1488 vssd1 vssd1 vccd1 vccd1 net1487 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_50_1863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1498 net1499 vssd1 vssd1 vccd1 vccd1 net1498 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_122_4056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_1298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19542_ clknet_leaf_115_clk _00486_ net1389 vssd1 vssd1 vccd1 vccd1 control.body\[852\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13416__A net672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16754_ obsg2.obstacleArray\[47\] net500 net486 obsg2.obstacleArray\[46\] vssd1 vssd1
+ vccd1 vccd1 _02433_ sky130_fd_sc_hd__a22o_1
X_13966_ ag2.body\[105\] net202 _08157_ ag2.body\[97\] vssd1 vssd1 vccd1 vccd1 _00186_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_88_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_31_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1514 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15705_ ag2.body\[369\] net141 _01629_ ag2.body\[361\] vssd1 vssd1 vccd1 vccd1 _00963_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_92_1465 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11207__Y _06180_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12917_ _07463_ net340 net335 vssd1 vssd1 vccd1 vccd1 _07656_ sky130_fd_sc_hd__and3b_1
X_16685_ _02212_ _02241_ _02252_ _02363_ _02244_ vssd1 vssd1 vccd1 vccd1 _02364_ sky130_fd_sc_hd__o221a_1
X_19473_ clknet_leaf_109_clk net2359 net1416 vssd1 vssd1 vccd1 vccd1 control.body\[927\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11294__A2 _04859_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13897_ ag2.body\[44\] net118 _08149_ ag2.body\[36\] vssd1 vssd1 vccd1 vccd1 _00125_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_1372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18424_ _03788_ _03801_ vssd1 vssd1 vccd1 vccd1 _03913_ sky130_fd_sc_hd__or2_1
X_15636_ ag2.body\[435\] net126 _01622_ ag2.body\[427\] vssd1 vssd1 vccd1 vccd1 _00901_
+ sky130_fd_sc_hd__a22o_1
X_12848_ net675 _07625_ vssd1 vssd1 vccd1 vccd1 _07626_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_14_Left_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_48_1781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_4428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_48_1792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_135_4439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15567_ ag2.body\[502\] net186 _01614_ ag2.body\[494\] vssd1 vssd1 vccd1 vccd1 _00840_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_84_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18355_ net2233 _08024_ _03818_ net464 _03850_ vssd1 vssd1 vccd1 vccd1 _01391_ sky130_fd_sc_hd__o221a_1
X_12779_ net307 _07592_ vssd1 vssd1 vccd1 vccd1 _07593_ sky130_fd_sc_hd__nor2_1
XFILLER_0_28_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_925 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_1667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17306_ ag2.body\[398\] net940 vssd1 vssd1 vccd1 vccd1 _02985_ sky130_fd_sc_hd__xor2_1
XFILLER_0_124_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14518_ net845 ag2.body\[312\] ag2.body\[319\] net796 _08674_ vssd1 vssd1 vccd1 vccd1
+ _08679_ sky130_fd_sc_hd__a221o_1
XFILLER_0_86_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18286_ net326 net325 vssd1 vssd1 vccd1 vccd1 _03782_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_25_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15498_ ag2.body\[552\] net113 _01607_ ag2.body\[544\] vssd1 vssd1 vccd1 vccd1 _00778_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_86_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_1513 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_25_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17237_ _02910_ _02913_ _02914_ _02915_ vssd1 vssd1 vccd1 vccd1 _02916_ sky130_fd_sc_hd__or4bb_1
XANTENNA__15193__B1 _01573_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14449_ net975 ag2.body\[227\] vssd1 vssd1 vccd1 vccd1 _08610_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_9_69 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_94_3181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold904 control.body\[811\] vssd1 vssd1 vccd1 vccd1 net2466 sky130_fd_sc_hd__dlygate4sd3_1
X_17168_ ag2.body\[594\] net722 net715 ag2.body\[595\] vssd1 vssd1 vccd1 vccd1 _02847_
+ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_94_3192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17277__B net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold915 control.body\[827\] vssd1 vssd1 vccd1 vccd1 net2477 sky130_fd_sc_hd__dlygate4sd3_1
Xhold926 _00703_ vssd1 vssd1 vccd1 vccd1 net2488 sky130_fd_sc_hd__dlygate4sd3_1
X_16119_ obsg2.obstacleArray\[77\] net430 vssd1 vssd1 vccd1 vccd1 _01798_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_90_3056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold937 control.body\[946\] vssd1 vssd1 vccd1 vccd1 net2499 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_3067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold948 _00478_ vssd1 vssd1 vccd1 vccd1 net2510 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_3078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17099_ _04098_ net854 net700 ag2.body\[302\] _02777_ vssd1 vssd1 vccd1 vccd1 _02778_
+ sky130_fd_sc_hd__a221o_1
Xhold959 control.body\[677\] vssd1 vssd1 vccd1 vccd1 net2521 sky130_fd_sc_hd__dlygate4sd3_1
X_09990_ net1217 control.body\[728\] vssd1 vssd1 vccd1 vccd1 _04963_ sky130_fd_sc_hd__xor2_1
XFILLER_0_110_732 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_23_Left_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_1608 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_08941_ net985 vssd1 vssd1 vccd1 vccd1 _03966_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16401__S net452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_1590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09804__A net1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19809_ clknet_leaf_124_clk _00753_ net1405 vssd1 vssd1 vccd1 vccd1 ag2.body\[591\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_105_3520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_105_3531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout187_A net218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11809__A1 net558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_3406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_3417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13045__B net646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_32_Left_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1096_A net1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_91_clk clknet_4_11__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_91_clk
+ sky130_fd_sc_hd__clkbuf_8
X_09424_ _04401_ net1726 _04399_ vssd1 vssd1 vccd1 vccd1 _00000_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_118_3914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09355_ sound_gen.osc1.stayCount\[12\] sound_gen.osc1.stayCount\[11\] _04355_ vssd1
+ vssd1 vccd1 vccd1 _04357_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout521_A net528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09635__C1 _04607_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_118_3925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_3936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_843 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout619_A net620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1263_A net1333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_1561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19365__CLK clknet_leaf_102_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09286_ sound_gen.osc1.freq\[1\] _04284_ _04286_ sound_gen.posDetector1.N\[0\] vssd1
+ vssd1 vccd1 vccd1 _04308_ sky130_fd_sc_hd__o22ai_4
XANTENNA_clkbuf_leaf_7_clk_A clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11993__B1 net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20515_ clknet_leaf_113_clk track.nextHighScore\[5\] net1403 vssd1 vssd1 vccd1 vccd1
+ track.highScore\[5\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_105_526 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_584 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout407_X net407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1430_A net1435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1051_X net1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13734__A1 net687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1149_X net1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20446_ clknet_leaf_42_clk _01333_ net1371 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[82\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__17187__B net938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout890_A net891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_41_Left_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout988_A net995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_1033 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17755__X _03434_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_2542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20377_ clknet_leaf_26_clk _01264_ net1344 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[13\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_73_2553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_2564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16684__B1 _02211_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10130_ _05099_ _05100_ _05101_ _05102_ vssd1 vssd1 vccd1 vccd1 _05103_ sky130_fd_sc_hd__or4_1
XANTENNA__17915__B _03531_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout776_X net776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10061_ ag2.body\[480\] net784 net744 ag2.body\[487\] vssd1 vssd1 vccd1 vccd1 _05034_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12170__B1 net544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout943_X net943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_86_2936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13820_ _08113_ _08114_ vssd1 vssd1 vccd1 vccd1 _08117_ sky130_fd_sc_hd__and2b_1
XANTENNA__09433__B net1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17931__A net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18189__B1 net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09469__A2 net1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout55_X net55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10579__B net1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_2357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_2368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_134_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13751_ net687 _08062_ net320 vssd1 vssd1 vccd1 vccd1 _08070_ sky130_fd_sc_hd__a21o_1
X_10963_ _05922_ _05935_ _05919_ vssd1 vssd1 vccd1 vccd1 _05936_ sky130_fd_sc_hd__o21ai_1
XANTENNA__17650__B net937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_2379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_82_clk clknet_4_14__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_82_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_98_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12702_ net344 net329 _07438_ vssd1 vssd1 vccd1 vccd1 _07555_ sky130_fd_sc_hd__and3_1
X_16470_ obsg2.obstacleArray\[52\] obsg2.obstacleArray\[53\] obsg2.obstacleArray\[54\]
+ obsg2.obstacleArray\[55\] net454 net397 vssd1 vssd1 vccd1 vccd1 _02149_ sky130_fd_sc_hd__mux4_1
XANTENNA__10484__B1 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1472 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13682_ net906 net434 _08025_ _08022_ vssd1 vssd1 vccd1 vccd1 track.nextCurrScore\[4\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_70_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10894_ _05859_ _05861_ _05864_ _05866_ vssd1 vssd1 vccd1 vccd1 _05867_ sky130_fd_sc_hd__or4_1
X_15421_ net2248 net81 _01598_ ag2.body\[620\] vssd1 vssd1 vccd1 vccd1 _00710_ sky130_fd_sc_hd__a22o_1
X_12633_ net388 _07518_ vssd1 vssd1 vccd1 vccd1 _07519_ sky130_fd_sc_hd__or2_2
XFILLER_0_112_1347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14067__A net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10595__A net1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_14_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18140_ net48 _03558_ _03704_ obsg2.obstacleArray\[67\] vssd1 vssd1 vccd1 vccd1 _03709_
+ sky130_fd_sc_hd__a31o_1
X_15352_ control.body\[694\] net72 _01591_ net2272 vssd1 vssd1 vccd1 vccd1 _00648_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_38_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12564_ net245 _07481_ _07482_ net1945 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[39\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_81_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_130_4303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_1060 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14303_ net828 ag2.body\[218\] _04070_ net1011 _08459_ vssd1 vssd1 vccd1 vccd1 _08464_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_13_1499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11984__B1 net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_1133 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11515_ net504 _06486_ _06487_ net759 vssd1 vssd1 vccd1 vccd1 _06488_ sky130_fd_sc_hd__a211o_1
XFILLER_0_108_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18071_ obsg2.obstacleArray\[43\] _03663_ net521 vssd1 vssd1 vccd1 vccd1 _01294_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_48_1507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18732__CLK clknet_leaf_141_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15283_ control.body\[744\] net78 _01584_ net2314 vssd1 vssd1 vccd1 vccd1 _00586_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__10882__X _05855_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19858__CLK clknet_leaf_93_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12495_ net292 _07440_ _07441_ net2056 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[11\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_124_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17022_ ag2.body\[329\] net736 net694 ag2.body\[335\] _02700_ vssd1 vssd1 vccd1 vccd1
+ _02701_ sky130_fd_sc_hd__a221o_1
XFILLER_0_123_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14234_ net1025 ag2.body\[485\] vssd1 vssd1 vccd1 vccd1 _08395_ sky130_fd_sc_hd__or2_1
XANTENNA__09448__X _04421_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11446_ net1134 control.body\[956\] vssd1 vssd1 vccd1 vccd1 _06419_ sky130_fd_sc_hd__or2_1
XANTENNA__14922__B1 _01543_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14165_ net1035 ag2.body\[204\] vssd1 vssd1 vccd1 vccd1 _08326_ sky130_fd_sc_hd__xor2_1
X_11377_ ag2.body\[473\] net778 _06345_ _06347_ _06349_ vssd1 vssd1 vccd1 vccd1 _06350_
+ sky130_fd_sc_hd__a2111o_1
XFILLER_0_0_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_128_4221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_128_4232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13116_ _07581_ _07639_ vssd1 vssd1 vccd1 vccd1 _07750_ sky130_fd_sc_hd__nor2_1
X_10328_ _05283_ _05286_ _05287_ _05300_ vssd1 vssd1 vccd1 vccd1 _05301_ sky130_fd_sc_hd__o22a_1
X_14096_ net820 ag2.body\[283\] ag2.body\[284\] net816 _08256_ vssd1 vssd1 vccd1 vccd1
+ _08257_ sky130_fd_sc_hd__o221a_1
X_18973_ clknet_leaf_8_clk img_gen.tracker.next_frame\[411\] net1270 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[411\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_52_1903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_4107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_4118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17924_ net539 net537 net460 net957 vssd1 vssd1 vccd1 vccd1 _03557_ sky130_fd_sc_hd__and4b_1
XANTENNA__17219__A2 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13047_ net225 _07716_ _07717_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[287\]
+ sky130_fd_sc_hd__o21bai_1
X_10259_ net767 control.body\[787\] control.body\[789\] net753 _05228_ vssd1 vssd1
+ vccd1 vccd1 _05232_ sky130_fd_sc_hd__a221oi_1
XTAP_TAPCELL_ROW_33_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14530__A net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12161__B1 net585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1240 net1243 vssd1 vssd1 vccd1 vccd1 net1240 sky130_fd_sc_hd__clkbuf_2
Xfanout1251 net1254 vssd1 vssd1 vccd1 vccd1 net1251 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_59_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17855_ _04280_ _07317_ img_gen.updater.commands.rR1.rainbowRNG\[1\] vssd1 vssd1
+ vccd1 vccd1 _03510_ sky130_fd_sc_hd__o21ba_1
Xfanout1262 net1263 vssd1 vssd1 vccd1 vccd1 net1262 sky130_fd_sc_hd__clkbuf_4
XANTENNA__15345__B net52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1273 net1275 vssd1 vssd1 vccd1 vccd1 net1273 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_94_1538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout1284 net1286 vssd1 vssd1 vccd1 vccd1 net1284 sky130_fd_sc_hd__clkbuf_4
X_16806_ ag2.body\[69\] net953 vssd1 vssd1 vccd1 vccd1 _02485_ sky130_fd_sc_hd__xor2_1
XANTENNA__13146__A net667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1295 net1296 vssd1 vssd1 vccd1 vccd1 net1295 sky130_fd_sc_hd__clkbuf_4
X_17786_ net1036 net1027 _03460_ vssd1 vssd1 vccd1 vccd1 _03463_ sky130_fd_sc_hd__and3_1
X_14998_ control.body\[1004\] net151 _01551_ control.body\[996\] vssd1 vssd1 vccd1
+ vccd1 _00334_ sky130_fd_sc_hd__a22o_1
XFILLER_0_89_855 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19525_ clknet_leaf_120_clk net2434 net1395 vssd1 vssd1 vccd1 vccd1 control.body\[867\]
+ sky130_fd_sc_hd__dfrtp_1
X_16737_ obsg2.obstacleArray\[54\] net487 net482 obsg2.obstacleArray\[53\] _02415_
+ vssd1 vssd1 vccd1 vccd1 _02416_ sky130_fd_sc_hd__a221o_1
X_13949_ ag2.body\[90\] net190 _08155_ ag2.body\[82\] vssd1 vssd1 vccd1 vccd1 _00171_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12985__A net337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_73_clk clknet_4_15__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_73_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_89_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_1718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19456_ clknet_leaf_109_clk net2410 net1420 vssd1 vssd1 vccd1 vccd1 control.body\[942\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_46_1729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_1403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16668_ obsg2.obstacleArray\[19\] net451 net393 vssd1 vssd1 vccd1 vccd1 _02347_ sky130_fd_sc_hd__o21a_1
XANTENNA__16176__B net424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18407_ _04639_ _03834_ _03896_ vssd1 vssd1 vccd1 vccd1 _03897_ sky130_fd_sc_hd__a21oi_1
X_15619_ ag2.body\[452\] net123 _01613_ ag2.body\[444\] vssd1 vssd1 vccd1 vccd1 _00886_
+ sky130_fd_sc_hd__a22o_1
X_19387_ clknet_leaf_102_clk _00331_ net1426 vssd1 vssd1 vccd1 vccd1 control.body\[1001\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__15953__A2 net196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16599_ net361 _02273_ _02277_ net357 vssd1 vssd1 vccd1 vccd1 _02278_ sky130_fd_sc_hd__o211a_1
XFILLER_0_130_1469 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09140_ ag2.body\[466\] vssd1 vssd1 vccd1 vccd1 _04165_ sky130_fd_sc_hd__inv_2
XANTENNA__20365__CLK clknet_leaf_21_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18338_ _04642_ _08026_ _08028_ vssd1 vssd1 vccd1 vccd1 _03834_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_44_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_96_3243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_1577 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_96_3254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11975__B1 net575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_96_3265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16904__B net885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09071_ ag2.body\[285\] vssd1 vssd1 vccd1 vccd1 _04096_ sky130_fd_sc_hd__inv_2
XFILLER_0_60_906 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16363__C1 net370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_3118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18269_ net516 _03773_ vssd1 vssd1 vccd1 vccd1 _01382_ sky130_fd_sc_hd__nor2_1
XANTENNA__10792__X _05765_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1618 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_3129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14705__A net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20300_ clknet_leaf_36_clk net1518 net1347 vssd1 vssd1 vccd1 vccd1 control.divider.count\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_128_1354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold701 img_gen.updater.commands.rR1.rainbowRNG\[11\] vssd1 vssd1 vccd1 vccd1 net2263
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10952__B net1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold712 control.body\[649\] vssd1 vssd1 vccd1 vccd1 net2274 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11727__B1 net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold723 control.body\[1048\] vssd1 vssd1 vccd1 vccd1 net2285 sky130_fd_sc_hd__dlygate4sd3_1
X_20231_ clknet_leaf_66_clk _01175_ net1476 vssd1 vssd1 vccd1 vccd1 ag2.body\[165\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_13_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_1353 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold734 control.body\[964\] vssd1 vssd1 vccd1 vccd1 net2296 sky130_fd_sc_hd__dlygate4sd3_1
Xhold745 control.body\[700\] vssd1 vssd1 vccd1 vccd1 net2307 sky130_fd_sc_hd__dlygate4sd3_1
Xhold756 control.body\[892\] vssd1 vssd1 vccd1 vccd1 net2318 sky130_fd_sc_hd__dlygate4sd3_1
Xhold767 sound_gen.osc1.stayCount\[0\] vssd1 vssd1 vccd1 vccd1 net2329 sky130_fd_sc_hd__dlygate4sd3_1
Xhold778 control.body\[1041\] vssd1 vssd1 vccd1 vccd1 net2340 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20162_ clknet_leaf_95_clk _01106_ net1441 vssd1 vssd1 vccd1 vccd1 ag2.body\[224\]
+ sky130_fd_sc_hd__dfrtp_4
X_09973_ net914 _04420_ net910 vssd1 vssd1 vccd1 vccd1 _04946_ sky130_fd_sc_hd__or3b_2
XFILLER_0_110_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold789 control.body\[1060\] vssd1 vssd1 vccd1 vccd1 net2351 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_1640 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20093_ clknet_leaf_78_clk _01037_ net1490 vssd1 vssd1 vccd1 vccd1 ag2.body\[299\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA_fanout1011_A net1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12152__B1 net579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1109_A ag2.x\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout471_A net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17091__B1 net964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_2_Right_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_1037 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_2800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1380_A net1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout736_A _04263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_64_clk clknet_4_13__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_64_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_94_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout1478_A net1505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1099_X net1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_2210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_2221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_81 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09407_ img_gen.updater.commands.mode\[0\] img_gen.updater.commands.mode\[1\] vssd1
+ vssd1 vccd1 vccd1 _04387_ sky130_fd_sc_hd__nor2_1
XANTENNA__18755__CLK clknet_leaf_15_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout524_X net524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15944__A2 net195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout903_A control.body_update.curr_length\[5\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_75_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13955__A1 _04421_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09338_ sound_gen.osc1.stayCount\[1\] sound_gen.osc1.stayCount\[0\] _04305_ vssd1
+ vssd1 vccd1 vccd1 _04342_ sky130_fd_sc_hd__and3_1
XFILLER_0_8_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_1220 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_2740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11023__B net1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09269_ sound_gen.osc1.stayCount\[11\] _04290_ net535 _04287_ sound_gen.osc1.stayCount\[12\]
+ vssd1 vssd1 vccd1 vccd1 _04292_ sky130_fd_sc_hd__o32a_1
XANTENNA__14615__A net987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_2604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_2615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11300_ net1096 control.body\[685\] vssd1 vssd1 vccd1 vccd1 _06273_ sky130_fd_sc_hd__xor2_1
X_12280_ _04272_ img_gen.updater.commands.cmd_num\[0\] _07240_ _07249_ vssd1 vssd1
+ vccd1 vccd1 _07250_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_65_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_1405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_2025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_2036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14380__A1 net834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11231_ net1171 _04244_ control.body\[863\] net744 _06194_ vssd1 vssd1 vccd1 vccd1
+ _06204_ sky130_fd_sc_hd__a221o_1
XANTENNA__14380__B2 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17449__A2 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16106__C1 _01743_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17926__A net48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20429_ clknet_leaf_23_clk _01316_ net1359 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[65\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_132_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16657__B1 net394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11162_ _06123_ _06130_ _06131_ _06132_ vssd1 vssd1 vccd1 vccd1 _06135_ sky130_fd_sc_hd__or4_2
XANTENNA__17645__B net868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_8_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10113_ _05079_ _05080_ _05081_ _05082_ _04551_ vssd1 vssd1 vccd1 vccd1 _05086_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_8_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09715__Y _04688_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14350__A net1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15970_ ag2.body\[141\] net198 _01658_ ag2.body\[133\] vssd1 vssd1 vccd1 vccd1 _01199_
+ sky130_fd_sc_hd__a22o_1
X_11093_ _04980_ _05920_ _06028_ vssd1 vssd1 vccd1 vccd1 _06066_ sky130_fd_sc_hd__a21o_1
XANTENNA__16409__B1 net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10044_ net1179 control.body\[898\] vssd1 vssd1 vccd1 vccd1 _05017_ sky130_fd_sc_hd__xor2_1
X_14921_ net895 _05399_ net66 vssd1 vssd1 vccd1 vccd1 _01543_ sky130_fd_sc_hd__and3_2
XTAP_TAPCELL_ROW_69_2419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15880__B2 ag2.body\[213\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12694__A1 net238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold50 img_gen.tracker.frame\[499\] vssd1 vssd1 vccd1 vccd1 net1612 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold61 img_gen.tracker.frame\[52\] vssd1 vssd1 vccd1 vccd1 net1623 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17640_ net691 ag2.body\[167\] _04050_ net872 vssd1 vssd1 vccd1 vccd1 _03319_ sky130_fd_sc_hd__a2bb2o_1
Xhold72 img_gen.tracker.frame\[102\] vssd1 vssd1 vccd1 vccd1 net1634 sky130_fd_sc_hd__dlygate4sd3_1
X_14852_ _08485_ _08489_ _08732_ _01522_ vssd1 vssd1 vccd1 vccd1 _01523_ sky130_fd_sc_hd__o211a_1
Xhold83 img_gen.tracker.frame\[61\] vssd1 vssd1 vccd1 vccd1 net1645 sky130_fd_sc_hd__dlygate4sd3_1
Xhold94 img_gen.tracker.frame\[527\] vssd1 vssd1 vccd1 vccd1 net1656 sky130_fd_sc_hd__dlygate4sd3_1
X_13803_ net625 net589 _08104_ _08105_ net1192 vssd1 vssd1 vccd1 vccd1 _00075_ sky130_fd_sc_hd__a32o_1
XANTENNA__17380__B net962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17571_ ag2.body\[576\] net879 vssd1 vssd1 vccd1 vccd1 _03250_ sky130_fd_sc_hd__xor2_1
X_14783_ net975 _04094_ _04095_ net1010 _01449_ vssd1 vssd1 vccd1 vccd1 _01454_ sky130_fd_sc_hd__a221o_1
X_11995_ img_gen.tracker.frame\[424\] net599 vssd1 vssd1 vccd1 vccd1 _06967_ sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_55_clk clknet_4_12__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_55_clk
+ sky130_fd_sc_hd__clkbuf_8
X_19310_ clknet_leaf_99_clk _00254_ net1445 vssd1 vssd1 vccd1 vccd1 control.body\[1084\]
+ sky130_fd_sc_hd__dfrtp_1
X_16522_ _02086_ _02199_ _02200_ _02107_ vssd1 vssd1 vccd1 vccd1 _02201_ sky130_fd_sc_hd__a211o_1
X_13734_ net687 _07202_ _07242_ _07259_ vssd1 vssd1 vccd1 vccd1 _00055_ sky130_fd_sc_hd__a22o_1
X_10946_ _05909_ _05910_ _05914_ _05918_ vssd1 vssd1 vccd1 vccd1 _05919_ sky130_fd_sc_hd__or4_4
XFILLER_0_42_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_52_clk_X clknet_leaf_52_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19241_ clknet_leaf_84_clk _00185_ net1481 vssd1 vssd1 vccd1 vccd1 ag2.body\[104\]
+ sky130_fd_sc_hd__dfrtp_4
X_13665_ net818 _08014_ _08015_ net998 vssd1 vssd1 vccd1 vccd1 obsrand1.next_randY\[0\]
+ sky130_fd_sc_hd__o31ai_1
X_16453_ obsg2.obstacleArray\[84\] obsg2.obstacleArray\[85\] obsg2.obstacleArray\[86\]
+ obsg2.obstacleArray\[87\] net458 net399 vssd1 vssd1 vccd1 vccd1 _02132_ sky130_fd_sc_hd__mux4_1
XANTENNA__15935__A2 net138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10877_ ag2.body\[530\] net1180 vssd1 vssd1 vccd1 vccd1 _05850_ sky130_fd_sc_hd__xor2_1
XFILLER_0_26_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12616_ net230 _07509_ _07510_ net2140 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[63\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_6_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15404_ net2315 net80 _01581_ net2480 vssd1 vssd1 vccd1 vccd1 _00695_ sky130_fd_sc_hd__a22o_1
XANTENNA__14228__C net1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16384_ _02061_ _02062_ vssd1 vssd1 vccd1 vccd1 _02063_ sky130_fd_sc_hd__and2_1
XFILLER_0_94_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19172_ clknet_leaf_53_clk _00116_ net1366 vssd1 vssd1 vccd1 vccd1 ag2.body\[35\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_6_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13596_ control.divider.count\[14\] control.divider.count\[13\] _07953_ vssd1 vssd1
+ vccd1 vccd1 _07971_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_22_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09614__A2 _04586_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18123_ obsg2.obstacleArray\[61\] _03697_ net524 vssd1 vssd1 vccd1 vccd1 _01312_
+ sky130_fd_sc_hd__o21a_1
X_15335_ control.body\[711\] net73 _01587_ net2454 vssd1 vssd1 vccd1 vccd1 _00633_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_42_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12547_ net334 _07471_ vssd1 vssd1 vccd1 vccd1 _07472_ sky130_fd_sc_hd__nand2_2
XFILLER_0_136_492 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14525__A net992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16896__B1 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18054_ net301 _03570_ vssd1 vssd1 vccd1 vccd1 _03652_ sky130_fd_sc_hd__nand2_1
XANTENNA__09619__A net1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15266_ net2591 net96 _01582_ net2061 vssd1 vssd1 vccd1 vccd1 _00571_ sky130_fd_sc_hd__a22o_1
XFILLER_0_13_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12478_ net1639 _07432_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[3\] sky130_fd_sc_hd__and2_1
XANTENNA_3 _03230_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_827 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_1500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14217_ _08373_ _08375_ _08377_ vssd1 vssd1 vccd1 vccd1 _08378_ sky130_fd_sc_hd__or3b_2
X_17005_ ag2.body\[499\] net853 vssd1 vssd1 vccd1 vccd1 _02684_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_39_1511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11429_ ag2.body\[394\] net1185 vssd1 vssd1 vccd1 vccd1 _06402_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_39_1522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15197_ control.body\[829\] net94 _01573_ net2518 vssd1 vssd1 vccd1 vccd1 _00511_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_65_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_197 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14148_ net987 ag2.body\[593\] vssd1 vssd1 vccd1 vccd1 _08309_ sky130_fd_sc_hd__xor2_1
XANTENNA__10932__A1 net775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10932__B2 net750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18956_ clknet_leaf_5_clk img_gen.tracker.next_frame\[394\] net1269 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[394\] sky130_fd_sc_hd__dfrtp_1
X_14079_ net988 ag2.body\[561\] vssd1 vssd1 vccd1 vccd1 _08240_ sky130_fd_sc_hd__xor2_1
XANTENNA__18628__CLK clknet_leaf_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12134__B1 net546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17907_ _01890_ net485 net381 vssd1 vssd1 vccd1 vccd1 _03542_ sky130_fd_sc_hd__and3b_2
XANTENNA__15075__B _04586_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18887_ clknet_leaf_25_clk img_gen.tracker.next_frame\[325\] net1343 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[325\] sky130_fd_sc_hd__dfrtp_1
Xfanout1070 net1071 vssd1 vssd1 vccd1 vccd1 net1070 sky130_fd_sc_hd__clkbuf_4
Xfanout1081 net1082 vssd1 vssd1 vccd1 vccd1 net1081 sky130_fd_sc_hd__clkbuf_4
X_17838_ net798 net224 vssd1 vssd1 vccd1 vccd1 _03496_ sky130_fd_sc_hd__nor2_1
Xfanout1092 net1093 vssd1 vssd1 vccd1 vccd1 net1092 sky130_fd_sc_hd__buf_4
XFILLER_0_83_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16820__B1 net706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12437__A1 net1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17769_ _02533_ _02837_ _03446_ _03447_ vssd1 vssd1 vccd1 vccd1 _03448_ sky130_fd_sc_hd__and4_1
XFILLER_0_77_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_46_clk clknet_4_7__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_46_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA__14831__C1 _01501_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1509 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19508_ clknet_leaf_113_clk _00452_ net1396 vssd1 vssd1 vccd1 vccd1 control.body\[882\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_18_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_3305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10947__B _05238_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_3316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19439_ clknet_leaf_108_clk _00383_ net1422 vssd1 vssd1 vccd1 vccd1 control.body\[957\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_130_1233 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_3327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11660__A2 net743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15926__A2 net124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_1277 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16634__B net445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_109 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11948__B1 net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09123_ ag2.body\[417\] vssd1 vssd1 vccd1 vccd1 _04148_ sky130_fd_sc_hd__inv_2
XFILLER_0_128_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17679__A2 net725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12070__C1 net561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16126__S net428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14435__A net980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20619__1562 vssd1 vssd1 vccd1 vccd1 net1562 _20619__1562/LO sky130_fd_sc_hd__conb_1
XFILLER_0_5_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1059_A net1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09054_ ag2.body\[248\] vssd1 vssd1 vccd1 vccd1 _04079_ sky130_fd_sc_hd__inv_2
XANTENNA__10682__B net1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_153 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19403__CLK clknet_leaf_103_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold520 img_gen.tracker.frame\[18\] vssd1 vssd1 vccd1 vccd1 net2082 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__14722__X _08883_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16650__A obsg2.obstacleArray\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold531 control.body\[905\] vssd1 vssd1 vccd1 vccd1 net2093 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1226_A net1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold542 _00558_ vssd1 vssd1 vccd1 vccd1 net2104 sky130_fd_sc_hd__dlygate4sd3_1
X_20214_ clknet_leaf_60_clk _01158_ net1466 vssd1 vssd1 vccd1 vccd1 ag2.body\[180\]
+ sky130_fd_sc_hd__dfrtp_4
Xhold553 img_gen.tracker.frame\[191\] vssd1 vssd1 vccd1 vccd1 net2115 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__17465__B net932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold564 _00224_ vssd1 vssd1 vccd1 vccd1 net2126 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__16103__A2 net426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_493 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold575 img_gen.tracker.frame\[87\] vssd1 vssd1 vccd1 vccd1 net2137 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10007__A_N net898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_1471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold586 img_gen.tracker.frame\[358\] vssd1 vssd1 vccd1 vccd1 net2148 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold597 control.divider.count\[0\] vssd1 vssd1 vccd1 vccd1 net2159 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout686_A _04393_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1235 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_1493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09956_ _04926_ _04927_ _04928_ vssd1 vssd1 vccd1 vccd1 _04929_ sky130_fd_sc_hd__or3_1
X_20145_ clknet_leaf_96_clk _01089_ net1449 vssd1 vssd1 vccd1 vccd1 ag2.body\[255\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA_fanout1014_X net1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12125__B1 net541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19553__CLK clknet_leaf_115_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20076_ clknet_leaf_77_clk _01020_ net1492 vssd1 vssd1 vccd1 vccd1 ag2.body\[314\]
+ sky130_fd_sc_hd__dfrtp_4
X_09887_ net920 net916 net923 net912 vssd1 vssd1 vccd1 vccd1 _04860_ sky130_fd_sc_hd__o31a_1
XANTENNA_fanout853_A net857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_449 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17912__C net298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16811__B1 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11018__B net1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout641_X net641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1383_X net1383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_37_clk clknet_4_5__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_37_clk
+ sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout739_X net739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10800_ ag2.body\[39\] net1055 vssd1 vssd1 vccd1 vccd1 _05773_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_16_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11780_ img_gen.tracker.frame\[182\] net621 net603 img_gen.tracker.frame\[185\] vssd1
+ vssd1 vccd1 vccd1 _06752_ sky130_fd_sc_hd__o22a_1
XANTENNA__09711__B net1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15378__B1 _01594_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10731_ ag2.body\[250\] net1182 vssd1 vssd1 vccd1 vccd1 _05704_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_7_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_1453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_1149 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13450_ _07581_ net302 vssd1 vssd1 vccd1 vccd1 _07892_ sky130_fd_sc_hd__nor2_1
X_10662_ net1179 control.body\[882\] vssd1 vssd1 vccd1 vccd1 _05635_ sky130_fd_sc_hd__xor2_1
XFILLER_0_12_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__11939__B1 net548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12401_ _07221_ _07346_ _07218_ vssd1 vssd1 vccd1 vccd1 _07365_ sky130_fd_sc_hd__and3b_1
XFILLER_0_118_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16327__C1 net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13381_ net274 _07864_ _07865_ net1997 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[473\]
+ sky130_fd_sc_hd__a22o_1
X_10593_ net1226 control.body\[824\] vssd1 vssd1 vccd1 vccd1 _05566_ sky130_fd_sc_hd__xor2_1
XFILLER_0_69_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15120_ net2637 net107 _01565_ control.body\[880\] vssd1 vssd1 vccd1 vccd1 _00442_
+ sky130_fd_sc_hd__a22o_1
X_12332_ _07255_ _07287_ vssd1 vssd1 vccd1 vccd1 _07299_ sky130_fd_sc_hd__nor2_1
XFILLER_0_49_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15051_ control.body\[954\] net163 _01558_ net2499 vssd1 vssd1 vccd1 vccd1 _00380_
+ sky130_fd_sc_hd__a22o_1
X_12263_ img_gen.updater.commands.count\[6\] img_gen.updater.commands.count\[5\] img_gen.updater.commands.count\[7\]
+ vssd1 vssd1 vccd1 vccd1 _07233_ sky130_fd_sc_hd__or3b_1
XANTENNA__15550__B1 net61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14002_ net1011 ag2.body\[511\] vssd1 vssd1 vccd1 vccd1 _08163_ sky130_fd_sc_hd__xor2_1
XFILLER_0_82_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11214_ _06183_ _06184_ _06185_ _06186_ vssd1 vssd1 vccd1 vccd1 _06187_ sky130_fd_sc_hd__and4_1
XFILLER_0_31_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17827__C1 net686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12194_ _07157_ _07158_ _07163_ _07164_ vssd1 vssd1 vccd1 vccd1 _07166_ sky130_fd_sc_hd__a22o_1
XFILLER_0_120_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18810_ clknet_leaf_3_clk img_gen.tracker.next_frame\[248\] net1259 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[248\] sky130_fd_sc_hd__dfrtp_1
X_11145_ ag2.body\[411\] net768 net749 ag2.body\[414\] _06117_ vssd1 vssd1 vccd1 vccd1
+ _06118_ sky130_fd_sc_hd__o221ai_1
XFILLER_0_124_1593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09445__Y _04418_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19790_ clknet_leaf_127_clk _00734_ net1328 vssd1 vssd1 vccd1 vccd1 ag2.body\[604\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__14080__A net1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__12116__B1 net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18741_ clknet_leaf_141_clk img_gen.tracker.next_frame\[179\] net1262 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[179\] sky130_fd_sc_hd__dfrtp_1
X_15953_ ag2.body\[158\] net196 _01656_ ag2.body\[150\] vssd1 vssd1 vccd1 vccd1 _01184_
+ sky130_fd_sc_hd__a22o_1
X_11076_ _04130_ net1113 net747 ag2.body\[367\] _06042_ vssd1 vssd1 vccd1 vccd1 _06049_
+ sky130_fd_sc_hd__o221a_1
XANTENNA_clkbuf_leaf_94_clk_A clknet_4_11__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17055__B1 net701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14904_ control.body\[1080\] net178 _01541_ control.body\[1072\] vssd1 vssd1 vccd1
+ vccd1 _00250_ sky130_fd_sc_hd__a22o_1
X_10027_ ag2.body\[506\] net1184 vssd1 vssd1 vccd1 vccd1 _05000_ sky130_fd_sc_hd__or2_1
X_18672_ clknet_leaf_26_clk img_gen.tracker.next_frame\[110\] net1339 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[110\] sky130_fd_sc_hd__dfrtp_1
X_15884_ ag2.body\[208\] net184 _01649_ ag2.body\[200\] vssd1 vssd1 vccd1 vccd1 _01122_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_91_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17623_ ag2.body\[184\] net881 vssd1 vssd1 vccd1 vccd1 _03302_ sky130_fd_sc_hd__xor2_1
XANTENNA__15623__B net56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14835_ _01502_ _01503_ _01504_ _01505_ vssd1 vssd1 vccd1 vccd1 _01506_ sky130_fd_sc_hd__and4_1
Xclkbuf_leaf_28_clk clknet_4_4__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_28_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_118_1386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17554_ ag2.body\[353\] net877 vssd1 vssd1 vccd1 vccd1 _03233_ sky130_fd_sc_hd__xor2_1
XFILLER_0_93_1390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14766_ net992 ag2.body\[97\] vssd1 vssd1 vccd1 vccd1 _08927_ sky130_fd_sc_hd__xor2_1
XANTENNA__13092__A1 net265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11978_ img_gen.tracker.frame\[556\] net605 net588 img_gen.tracker.frame\[562\] _06949_
+ vssd1 vssd1 vccd1 vccd1 _06950_ sky130_fd_sc_hd__o221a_1
XFILLER_0_58_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_1363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16505_ obsg2.obstacleArray\[10\] obsg2.obstacleArray\[11\] net456 vssd1 vssd1 vccd1
+ vccd1 _02184_ sky130_fd_sc_hd__mux2_1
XANTENNA__15369__B1 _01593_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13717_ track.highScore\[6\] _08030_ net356 vssd1 vssd1 vccd1 vccd1 track.nextHighScore\[6\]
+ sky130_fd_sc_hd__mux2_4
X_10929_ net780 control.body\[1033\] _05901_ vssd1 vssd1 vccd1 vccd1 _05902_ sky130_fd_sc_hd__a21oi_1
XANTENNA__15910__Y _01652_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17485_ _03157_ _03158_ _03162_ _03163_ _03154_ vssd1 vssd1 vccd1 vccd1 _03164_ sky130_fd_sc_hd__a2111oi_1
X_14697_ net993 _04110_ _04111_ net1041 _08857_ vssd1 vssd1 vccd1 vccd1 _08858_ sky130_fd_sc_hd__o221a_1
X_19224_ clknet_leaf_75_clk _00168_ net1494 vssd1 vssd1 vccd1 vccd1 ag2.body\[87\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_6_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13711__X track.nextHighScore\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16436_ obsg2.obstacleArray\[88\] obsg2.obstacleArray\[89\] net458 vssd1 vssd1 vccd1
+ vccd1 _02115_ sky130_fd_sc_hd__mux2_1
XANTENNA__10850__B1 net1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13648_ control.divider.count\[16\] _08004_ _08006_ net221 vssd1 vssd1 vccd1 vccd1
+ control.divider.next_count\[16\] sky130_fd_sc_hd__o211a_1
XFILLER_0_128_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_32_clk_A clknet_4_5__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14592__A1 net829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19155_ clknet_leaf_52_clk _00099_ net1367 vssd1 vssd1 vccd1 vccd1 ag2.body\[19\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__19426__CLK clknet_leaf_111_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13579_ _07953_ vssd1 vssd1 vccd1 vccd1 _07954_ sky130_fd_sc_hd__inv_2
X_16367_ net416 _02043_ _02045_ net372 vssd1 vssd1 vccd1 vccd1 _02046_ sky130_fd_sc_hd__a211o_1
XANTENNA__10783__A net1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14255__A net994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18106_ obsg2.obstacleArray\[55\] _03686_ net524 vssd1 vssd1 vccd1 vccd1 _01306_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_87_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15318_ control.body\[727\] net74 _01588_ net2322 vssd1 vssd1 vccd1 vccd1 _00617_
+ sky130_fd_sc_hd__a22o_1
X_16298_ net418 _01976_ _01975_ net369 vssd1 vssd1 vccd1 vccd1 _01977_ sky130_fd_sc_hd__a211o_1
XFILLER_0_81_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19086_ clknet_leaf_9_clk img_gen.tracker.next_frame\[524\] net1272 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[524\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_112_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18037_ obsg2.obstacleArray\[31\] _03641_ net532 vssd1 vssd1 vccd1 vccd1 _01282_
+ sky130_fd_sc_hd__o21a_1
XANTENNA_clkbuf_leaf_47_clk_A clknet_4_7__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_1410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15249_ control.body\[779\] net99 _01579_ net2135 vssd1 vssd1 vccd1 vccd1 _00557_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_23_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_99_Right_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17285__B net966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16097__A1 _01742_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10007__B net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout307 _07445_ vssd1 vssd1 vccd1 vccd1 net307 sky130_fd_sc_hd__buf_4
X_09810_ _04418_ _04723_ _04782_ _04694_ _04711_ vssd1 vssd1 vccd1 vccd1 _04783_ sky130_fd_sc_hd__o2111a_1
Xfanout318 _01818_ vssd1 vssd1 vccd1 vccd1 net318 sky130_fd_sc_hd__clkbuf_4
X_19988_ clknet_leaf_66_clk _00932_ net1475 vssd1 vssd1 vccd1 vccd1 ag2.body\[402\]
+ sky130_fd_sc_hd__dfrtp_4
Xfanout329 net330 vssd1 vssd1 vccd1 vccd1 net329 sky130_fd_sc_hd__buf_2
XANTENNA__12107__B1 net593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09741_ ag2.body\[357\] net1113 vssd1 vssd1 vccd1 vccd1 _04714_ sky130_fd_sc_hd__xnor2_1
X_18939_ clknet_leaf_143_clk img_gen.tracker.next_frame\[377\] net1288 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[377\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__12658__A1 net240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13855__B1 _08134_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_65 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17046__B1 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_105_clk_A clknet_4_10__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11119__A net1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09672_ _04643_ _04644_ vssd1 vssd1 vccd1 vccd1 _04645_ sky130_fd_sc_hd__or2_1
XFILLER_0_119_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15533__B net62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_1453 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_6_Left_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_19_clk clknet_4_3__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_19_clk
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_90_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout267_A net268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11618__C1 net1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1497 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_1452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10677__B net1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16557__C1 net359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1176_A net1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16309__C1 net418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout601_A net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14165__A net1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09106_ ag2.body\[369\] vssd1 vssd1 vccd1 vccd1 _04131_ sky130_fd_sc_hd__inv_2
XFILLER_0_72_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_1500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19919__CLK clknet_leaf_52_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14335__A1 net818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09037_ ag2.body\[200\] vssd1 vssd1 vccd1 vccd1 _04062_ sky130_fd_sc_hd__inv_2
XFILLER_0_130_421 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14335__B2 net812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1131_X net1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17907__C net381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1229_X net1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09546__X _04519_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17195__B net852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold350 img_gen.tracker.frame\[209\] vssd1 vssd1 vccd1 vccd1 net1912 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout970_A net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold361 toggle1.bcd_tens\[2\] vssd1 vssd1 vccd1 vccd1 net1923 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout591_X net591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16088__A1 net348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold372 img_gen.tracker.frame\[32\] vssd1 vssd1 vccd1 vccd1 net1934 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout689_X net689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17763__X _03442_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold383 img_gen.tracker.frame\[39\] vssd1 vssd1 vccd1 vccd1 net1945 sky130_fd_sc_hd__dlygate4sd3_1
Xhold394 img_gen.tracker.frame\[258\] vssd1 vssd1 vccd1 vccd1 net1956 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout830 net831 vssd1 vssd1 vccd1 vccd1 net830 sky130_fd_sc_hd__clkbuf_4
Xfanout841 net847 vssd1 vssd1 vccd1 vccd1 net841 sky130_fd_sc_hd__clkbuf_2
Xfanout852 net857 vssd1 vssd1 vccd1 vccd1 net852 sky130_fd_sc_hd__buf_4
XFILLER_0_99_1065 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_20128_ clknet_leaf_80_clk _01072_ net1485 vssd1 vssd1 vccd1 vccd1 ag2.body\[270\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__19976__RESET_B net1470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09939_ ag2.body\[24\] net784 net768 ag2.body\[27\] _04906_ vssd1 vssd1 vccd1 vccd1
+ _04912_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout856_X net856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout863 net867 vssd1 vssd1 vccd1 vccd1 net863 sky130_fd_sc_hd__buf_4
Xfanout874 net878 vssd1 vssd1 vccd1 vccd1 net874 sky130_fd_sc_hd__buf_4
XANTENNA__17037__B1 net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout885 net886 vssd1 vssd1 vccd1 vccd1 net885 sky130_fd_sc_hd__buf_4
XANTENNA__11029__A net1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout896 net897 vssd1 vssd1 vccd1 vccd1 net896 sky130_fd_sc_hd__clkbuf_4
X_12950_ _07672_ net266 _07670_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[235\]
+ sky130_fd_sc_hd__mux2_1
X_20059_ clknet_leaf_72_clk _01003_ net1501 vssd1 vssd1 vccd1 vccd1 ag2.body\[329\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__19905__RESET_B net1464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1050 control.body\[699\] vssd1 vssd1 vccd1 vccd1 net2612 sky130_fd_sc_hd__dlygate4sd3_1
X_11901_ img_gen.tracker.frame\[58\] net580 net558 _06872_ vssd1 vssd1 vccd1 vccd1
+ _06873_ sky130_fd_sc_hd__o211ai_1
Xhold1061 control.body\[930\] vssd1 vssd1 vccd1 vccd1 net2623 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1072 control.body\[891\] vssd1 vssd1 vccd1 vccd1 net2634 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11971__B net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15599__B1 _01619_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1083 control.body\[1012\] vssd1 vssd1 vccd1 vccd1 net2645 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__15443__B net54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12881_ _07434_ _07639_ vssd1 vssd1 vccd1 vccd1 _07641_ sky130_fd_sc_hd__nor2_1
Xhold1094 control.body\[1002\] vssd1 vssd1 vccd1 vccd1 net2656 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_119_1673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14620_ net1025 _03997_ ag2.body\[63\] net790 _08775_ vssd1 vssd1 vccd1 vccd1 _08781_
+ sky130_fd_sc_hd__o221a_1
X_11832_ img_gen.tracker.frame\[530\] net613 net596 img_gen.tracker.frame\[533\] vssd1
+ vssd1 vccd1 vccd1 _06804_ sky130_fd_sc_hd__o22a_1
XFILLER_0_90_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14551_ _08700_ _08701_ _08702_ _08703_ _08711_ vssd1 vssd1 vccd1 vccd1 _08712_ sky130_fd_sc_hd__a221o_2
X_11763_ _06732_ _06734_ net559 vssd1 vssd1 vccd1 vccd1 _06735_ sky130_fd_sc_hd__mux2_1
XANTENNA__12821__A1 net278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13502_ net230 _07912_ _07913_ net1829 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[546\]
+ sky130_fd_sc_hd__a22o_1
X_10714_ ag2.body\[616\] net1219 vssd1 vssd1 vccd1 vccd1 _05687_ sky130_fd_sc_hd__xor2_1
X_14482_ net998 _04156_ _04159_ net1008 _08641_ vssd1 vssd1 vccd1 vccd1 _08643_ sky130_fd_sc_hd__a221o_1
X_17270_ _02946_ _02947_ _02948_ vssd1 vssd1 vccd1 vccd1 _02949_ sky130_fd_sc_hd__and3_1
XFILLER_0_83_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11694_ img_gen.tracker.frame\[119\] net586 net547 img_gen.tracker.frame\[116\] _06665_
+ vssd1 vssd1 vccd1 vccd1 _06666_ sky130_fd_sc_hd__o221a_1
XFILLER_0_138_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16221_ net956 _01888_ vssd1 vssd1 vccd1 vccd1 _01900_ sky130_fd_sc_hd__nand2_1
X_13433_ net257 _07884_ _07885_ net1914 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[505\]
+ sky130_fd_sc_hd__a22o_1
X_10645_ _05588_ _05598_ _05600_ _05610_ _05617_ vssd1 vssd1 vccd1 vccd1 _05618_ sky130_fd_sc_hd__o32a_2
XFILLER_0_130_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16152_ net379 _01830_ _01829_ net349 vssd1 vssd1 vccd1 vccd1 _01831_ sky130_fd_sc_hd__a211o_1
XANTENNA__19599__CLK clknet_leaf_118_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13364_ net228 _07858_ _07859_ net2020 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[462\]
+ sky130_fd_sc_hd__a22o_1
X_10576_ ag2.body\[186\] net1177 vssd1 vssd1 vccd1 vccd1 _05549_ sky130_fd_sc_hd__or2_1
XANTENNA__14326__A1 net842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15103_ net2150 net183 _01564_ control.body\[896\] vssd1 vssd1 vccd1 vccd1 _00426_
+ sky130_fd_sc_hd__a22o_1
X_12315_ _07271_ _07277_ _07281_ net687 vssd1 vssd1 vccd1 vccd1 _07282_ sky130_fd_sc_hd__o31a_1
XFILLER_0_126_1633 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14326__B2 net800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16083_ obsg2.obstacleArray\[99\] net430 net376 _01761_ vssd1 vssd1 vccd1 vccd1 _01762_
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_133_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_1498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13295_ net234 _07831_ _07832_ net1741 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[420\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_122_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10108__A net1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19911_ clknet_leaf_54_clk _00855_ net1457 vssd1 vssd1 vccd1 vccd1 ag2.body\[485\]
+ sky130_fd_sc_hd__dfrtp_4
X_15034_ control.body\[970\] net163 _01557_ net2218 vssd1 vssd1 vccd1 vccd1 _00364_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_32_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_1677 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12246_ img_gen.updater.commands.cmd_num\[0\] _07215_ img_gen.updater.commands.cmd_num\[1\]
+ vssd1 vssd1 vccd1 vccd1 _07216_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12888__A1 net245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1605 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19842_ clknet_leaf_92_clk _00786_ net1412 vssd1 vssd1 vccd1 vccd1 ag2.body\[544\]
+ sky130_fd_sc_hd__dfrtp_4
X_12177_ net317 _07147_ net480 vssd1 vssd1 vccd1 vccd1 _07149_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_23_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11128_ control.body\[867\] net1148 vssd1 vssd1 vccd1 vccd1 _06101_ sky130_fd_sc_hd__and2b_1
X_19773_ clknet_leaf_19_clk _00717_ net1331 vssd1 vssd1 vccd1 vccd1 ag2.body\[619\]
+ sky130_fd_sc_hd__dfrtp_4
X_16985_ ag2.body\[94\] net700 net932 _04022_ vssd1 vssd1 vccd1 vccd1 _02664_ sky130_fd_sc_hd__a22o_1
XFILLER_0_3_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18724_ clknet_leaf_142_clk img_gen.tracker.next_frame\[162\] net1257 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[162\] sky130_fd_sc_hd__dfrtp_1
X_11059_ ag2.body\[433\] net1198 vssd1 vssd1 vccd1 vccd1 _06032_ sky130_fd_sc_hd__xnor2_1
X_15936_ ag2.body\[174\] net138 _01655_ ag2.body\[166\] vssd1 vssd1 vccd1 vccd1 _01168_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__18010__A net351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20618__1561 vssd1 vssd1 vccd1 vccd1 net1561 _20618__1561/LO sky130_fd_sc_hd__conb_1
XFILLER_0_91_1305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18655_ clknet_leaf_16_clk img_gen.tracker.next_frame\[93\] net1315 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[93\] sky130_fd_sc_hd__dfrtp_1
X_15867_ ag2.body\[225\] net201 _01647_ ag2.body\[217\] vssd1 vssd1 vccd1 vccd1 _01107_
+ sky130_fd_sc_hd__a22o_1
X_17606_ _04149_ net867 _03283_ _03284_ vssd1 vssd1 vccd1 vccd1 _03285_ sky130_fd_sc_hd__a211o_1
XFILLER_0_56_1469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14818_ _01480_ _01481_ _01482_ _01488_ vssd1 vssd1 vccd1 vccd1 _01489_ sky130_fd_sc_hd__or4_4
XFILLER_0_34_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18586_ clknet_leaf_14_clk img_gen.tracker.next_frame\[24\] net1276 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[24\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_133_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15798_ ag2.body\[291\] net207 _01640_ ag2.body\[283\] vssd1 vssd1 vccd1 vccd1 _01045_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__09808__A2 _04759_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16002__A_N net883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11076__B1 net747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17049__A2_N net711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17537_ ag2.body\[275\] net854 vssd1 vssd1 vccd1 vccd1 _03216_ sky130_fd_sc_hd__xnor2_1
X_14749_ net839 ag2.body\[105\] ag2.body\[111\] net796 _08905_ vssd1 vssd1 vccd1 vccd1
+ _08910_ sky130_fd_sc_hd__o221a_1
XFILLER_0_8_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16003__A1 net539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_1609 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17200__B1 net931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17468_ _04193_ net874 net863 _04194_ _03146_ vssd1 vssd1 vccd1 vccd1 _03147_ sky130_fd_sc_hd__a221o_1
XFILLER_0_117_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__20133__RESET_B net1449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19207_ clknet_leaf_86_clk _00151_ net1459 vssd1 vssd1 vccd1 vccd1 ag2.body\[70\]
+ sky130_fd_sc_hd__dfrtp_4
X_16419_ net401 _02097_ net366 vssd1 vssd1 vccd1 vccd1 _02098_ sky130_fd_sc_hd__o21a_1
XFILLER_0_89_1289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17399_ _04185_ net863 net692 ag2.body\[511\] _03076_ vssd1 vssd1 vccd1 vccd1 _03078_
+ sky130_fd_sc_hd__a221o_1
X_19138_ clknet_leaf_132_clk img_gen.control.next\[0\] net1303 vssd1 vssd1 vccd1 vccd1
+ img_gen.control.current\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_70_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12040__A2 net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18528__RESET_B net1292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18966__CLK clknet_leaf_5_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19069_ clknet_leaf_28_clk img_gen.tracker.next_frame\[507\] net1336 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[507\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__09992__B2 net758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16404__S net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_8_clk clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_8_clk
+ sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_114_3791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10960__B net1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_3666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_110_3677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_1198 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_110_3688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17267__B1 net707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout104 net114 vssd1 vssd1 vccd1 vccd1 net104 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_59_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout115 net117 vssd1 vssd1 vccd1 vccd1 net115 sky130_fd_sc_hd__buf_2
Xfanout126 net127 vssd1 vssd1 vccd1 vccd1 net126 sky130_fd_sc_hd__buf_2
Xfanout137 net139 vssd1 vssd1 vccd1 vccd1 net137 sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout148 net154 vssd1 vssd1 vccd1 vccd1 net148 sky130_fd_sc_hd__buf_2
XANTENNA__13048__B _07306_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout159 net161 vssd1 vssd1 vccd1 vccd1 net159 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_129_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16490__A1 _02075_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09724_ net894 net899 net902 net907 vssd1 vssd1 vccd1 vccd1 _04697_ sky130_fd_sc_hd__or4_4
XANTENNA__14247__A1_N net837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09542__A net1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09655_ net1121 control.body\[748\] vssd1 vssd1 vccd1 vccd1 _04628_ sky130_fd_sc_hd__xor2_1
XANTENNA__15263__B net52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19316__RESET_B net1435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout551_A net552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11854__A2 net590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1293_A net1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11136__X _06109_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_3_2_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_3_2_0_clk sky130_fd_sc_hd__clkbuf_8
X_09586_ net1157 control.body\[907\] vssd1 vssd1 vccd1 vccd1 _04559_ sky130_fd_sc_hd__xor2_1
XANTENNA__11067__B1 _06039_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12803__A1 net239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10200__B net1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1081_X net1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1460_A net1461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout816_A _03969_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout437_X net437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1179_X net1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09680__B1 net1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16094__B net425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_1329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_1489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10430_ net1110 control.body\[1069\] vssd1 vssd1 vccd1 vccd1 _05403_ sky130_fd_sc_hd__or2_1
XFILLER_0_116_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1020 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12031__A2 net611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10361_ _04983_ _05325_ _05329_ _05333_ vssd1 vssd1 vccd1 vccd1 _05334_ sky130_fd_sc_hd__or4_2
XFILLER_0_103_432 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14623__A net1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12100_ img_gen.tracker.frame\[372\] net628 net595 img_gen.tracker.frame\[381\] vssd1
+ vssd1 vccd1 vccd1 _07072_ sky130_fd_sc_hd__a22o_1
X_13080_ _07733_ net265 _07731_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[304\]
+ sky130_fd_sc_hd__mux2_1
X_10292_ _05261_ _05262_ _05263_ _05264_ vssd1 vssd1 vccd1 vccd1 _05265_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout973_X net973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19194__Q ag2.body\[57\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10870__B net1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12031_ img_gen.tracker.frame\[27\] net611 net576 _07002_ vssd1 vssd1 vccd1 vccd1
+ _07003_ sky130_fd_sc_hd__a211o_1
Xhold180 img_gen.tracker.frame\[50\] vssd1 vssd1 vccd1 vccd1 net1742 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09436__B net1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold191 img_gen.tracker.frame\[210\] vssd1 vssd1 vccd1 vccd1 net1753 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__19121__CLK clknet_leaf_141_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18101__Y _03683_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout660 net661 vssd1 vssd1 vccd1 vccd1 net660 sky130_fd_sc_hd__clkbuf_2
Xfanout671 net672 vssd1 vssd1 vccd1 vccd1 net671 sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_69_Left_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16770_ obsg2.obstacleArray\[8\] net493 net484 obsg2.obstacleArray\[9\] _02448_ vssd1
+ vssd1 vccd1 vccd1 _02449_ sky130_fd_sc_hd__a221o_1
Xfanout682 net684 vssd1 vssd1 vccd1 vccd1 net682 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12098__A2 net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13982_ _06240_ net61 vssd1 vssd1 vccd1 vccd1 _08159_ sky130_fd_sc_hd__nor2_2
Xfanout693 net694 vssd1 vssd1 vccd1 vccd1 net693 sky130_fd_sc_hd__clkbuf_4
XANTENNA__13295__A1 net234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09499__B1 net642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15721_ _04418_ net60 vssd1 vssd1 vccd1 vccd1 _01631_ sky130_fd_sc_hd__nor2_2
XANTENNA__17940__Y _03570_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12933_ _07664_ net266 _07662_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[226\]
+ sky130_fd_sc_hd__mux2_1
XANTENNA__11845__A2 net617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_1647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_1521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18440_ _03912_ _03928_ _03791_ vssd1 vssd1 vccd1 vccd1 _03929_ sky130_fd_sc_hd__a21oi_1
X_15652_ ag2.body\[417\] net139 _01624_ ag2.body\[409\] vssd1 vssd1 vccd1 vccd1 _00915_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__13047__A1 net225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_1554 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12864_ _06672_ _07545_ vssd1 vssd1 vccd1 vccd1 _07633_ sky130_fd_sc_hd__nor2_1
XANTENNA__18839__CLK clknet_leaf_4_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_953 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_1345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14603_ net985 _04034_ ag2.body\[132\] net815 _08763_ vssd1 vssd1 vccd1 vccd1 _08764_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_5_1418 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18371_ net464 _08143_ _03823_ _03863_ vssd1 vssd1 vccd1 vccd1 _03864_ sky130_fd_sc_hd__a31o_1
X_11815_ net568 _06786_ _06784_ vssd1 vssd1 vccd1 vccd1 _06787_ sky130_fd_sc_hd__a21oi_1
XANTENNA__15901__B net55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15583_ ag2.body\[483\] net130 _01617_ ag2.body\[475\] vssd1 vssd1 vccd1 vccd1 _00853_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_9_1598 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12795_ net278 _07599_ _07600_ net2037 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[152\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_96_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_1389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17322_ net719 ag2.body\[219\] _04069_ net863 vssd1 vssd1 vccd1 vccd1 _03001_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_51_1355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11746_ net576 _06711_ _06713_ _06716_ net474 vssd1 vssd1 vccd1 vccd1 _06718_ sky130_fd_sc_hd__a311o_1
X_14534_ net846 ag2.body\[248\] ag2.body\[253\] net808 _08694_ vssd1 vssd1 vccd1 vccd1
+ _08695_ sky130_fd_sc_hd__a221o_1
XFILLER_0_3_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_137_4492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_78_Left_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_1399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17253_ ag2.body\[548\] net962 vssd1 vssd1 vccd1 vccd1 _02932_ sky130_fd_sc_hd__xor2_1
XANTENNA__18989__CLK clknet_leaf_8_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14465_ net1001 ag2.body\[264\] vssd1 vssd1 vccd1 vccd1 _08626_ sky130_fd_sc_hd__or2_1
X_11677_ net1174 net1123 vssd1 vssd1 vccd1 vccd1 _06649_ sky130_fd_sc_hd__xor2_4
XFILLER_0_24_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_133_4367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_133_4378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16204_ _01881_ _01882_ net346 vssd1 vssd1 vccd1 vccd1 _01883_ sky130_fd_sc_hd__mux2_1
XANTENNA__11222__A net1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_133_4389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10628_ net1045 control.body\[671\] vssd1 vssd1 vccd1 vccd1 _05601_ sky130_fd_sc_hd__nand2_1
X_13416_ net672 _07878_ vssd1 vssd1 vccd1 vccd1 _07879_ sky130_fd_sc_hd__nor2_1
X_14396_ net839 ag2.body\[121\] _04030_ net985 _08556_ vssd1 vssd1 vccd1 vccd1 _08557_
+ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_12_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12022__A2 net612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17184_ ag2.body\[570\] net859 vssd1 vssd1 vccd1 vccd1 _02863_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_12_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16135_ net737 net732 _01691_ vssd1 vssd1 vccd1 vccd1 _01814_ sky130_fd_sc_hd__and3_1
XFILLER_0_3_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13347_ net332 _07515_ _07813_ vssd1 vssd1 vccd1 vccd1 _07852_ sky130_fd_sc_hd__and3_1
X_10559_ _04191_ net1132 _04416_ _05530_ _05531_ vssd1 vssd1 vccd1 vccd1 _05532_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_126_1441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16066_ obsg2.obstacleArray\[104\] net421 net373 _01744_ vssd1 vssd1 vccd1 vccd1
+ _01745_ sky130_fd_sc_hd__o211a_1
XFILLER_0_45_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13278_ net384 _07464_ vssd1 vssd1 vccd1 vccd1 _07825_ sky130_fd_sc_hd__nor2_2
XANTENNA__19898__RESET_B net1464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_1485 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_12229_ img_gen.updater.commands.cmd_num\[3\] _07197_ vssd1 vssd1 vccd1 vccd1 _07199_
+ sky130_fd_sc_hd__or2_1
X_15017_ control.body\[989\] net167 _01553_ control.body\[981\] vssd1 vssd1 vccd1
+ vccd1 _00351_ sky130_fd_sc_hd__a22o_1
XFILLER_0_27_1593 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_87_Left_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19825_ clknet_leaf_124_clk _00769_ net1408 vssd1 vssd1 vccd1 vccd1 ag2.body\[575\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_55_1989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17563__B net950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16472__A1 net364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19756_ clknet_leaf_129_clk _00700_ net1326 vssd1 vssd1 vccd1 vccd1 control.body\[634\]
+ sky130_fd_sc_hd__dfrtp_1
X_16968_ ag2.body\[408\] net884 vssd1 vssd1 vccd1 vccd1 _02647_ sky130_fd_sc_hd__xor2_1
XANTENNA__13286__A1 net255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12089__A2 net630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18707_ clknet_leaf_143_clk img_gen.tracker.next_frame\[145\] net1255 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[145\] sky130_fd_sc_hd__dfrtp_1
X_15919_ _04831_ net61 vssd1 vssd1 vccd1 vccd1 _01653_ sky130_fd_sc_hd__nor2_2
XFILLER_0_91_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19687_ clknet_leaf_135_clk _00631_ net1302 vssd1 vssd1 vccd1 vccd1 control.body\[709\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11836__A2 net622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16899_ _02572_ _02577_ vssd1 vssd1 vccd1 vccd1 _02578_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_79_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17421__B1 net720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09440_ _04403_ _04404_ _04410_ _04411_ _04405_ vssd1 vssd1 vccd1 vccd1 _04413_ sky130_fd_sc_hd__a221o_1
XFILLER_0_56_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18638_ clknet_leaf_131_clk img_gen.tracker.next_frame\[76\] net1312 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[76\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_1581 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10301__A net1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19764__CLK clknet_leaf_127_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16775__A2 net503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_103_3470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09371_ sound_gen.osc1.stayCount\[19\] _04361_ net270 vssd1 vssd1 vccd1 vccd1 _04371_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_47_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14786__A1 net991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18569_ clknet_leaf_15_clk img_gen.tracker.next_frame\[7\] net1313 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[7\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__14786__B2 net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20600_ net1532 vssd1 vssd1 vccd1 vccd1 gpio_oeb[12] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_96_Left_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_1597 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10955__B net1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20531_ clknet_leaf_114_clk _01396_ net1398 vssd1 vssd1 vccd1 vccd1 toggle1.bcd_ones\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_74_477 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout132_A net144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1649 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_116_3853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_116_3864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20462_ clknet_leaf_28_clk _01349_ net1336 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[98\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__13210__A1 net241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_116_3875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10024__A1 _04967_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_3728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_1313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10024__B2 _04996_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_112_3739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20393_ clknet_leaf_38_clk _01280_ net1355 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[29\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_113_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10971__A net1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14443__A net1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1041_A net1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_1661 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19144__CLK clknet_leaf_51_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1139_A net1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09537__A net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10690__B net1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13059__A net338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout599_A net602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17754__A _03428_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1693 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout1306_A net1310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_71_2481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17473__B net953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_71_2492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout387_X net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_1301 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13277__A1 net280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_1345 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09707_ ag2.body\[246\] net1085 vssd1 vssd1 vccd1 vccd1 _04680_ sky130_fd_sc_hd__xor2_1
XANTENNA__19150__RESET_B net1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout933_A net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout554_X net554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1378 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17412__B1 net740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_1621 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__10211__A net1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13029__A1 net259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09638_ net745 control.body\[1023\] control.body\[1020\] net761 vssd1 vssd1 vccd1
+ vccd1 _04611_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_69_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16766__A2 net502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_2875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout45_A net46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17963__A1 net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20055__RESET_B net1502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_2886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_1665 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_84_2897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14777__A1 net983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout721_X net721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15721__B net60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09569_ ag2.body\[202\] net776 net762 ag2.body\[204\] vssd1 vssd1 vccd1 vccd1 _04542_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__15974__B1 net663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14777__B2 net795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout819_X net819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_2296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11600_ obsg2.obstacleArray\[18\] obsg2.obstacleArray\[22\] net514 vssd1 vssd1 vccd1
+ vccd1 _06573_ sky130_fd_sc_hd__mux2_1
XANTENNA__13522__A net226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12580_ _06671_ _07310_ vssd1 vssd1 vccd1 vccd1 _07490_ sky130_fd_sc_hd__or2_2
XFILLER_0_66_956 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10865__B _05781_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_1705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_1304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11531_ net777 _06492_ vssd1 vssd1 vccd1 vccd1 _06504_ sky130_fd_sc_hd__or2_1
XANTENNA__17929__A net463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10263__B2 _05235_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14250_ net984 _04197_ _04198_ net1021 _08408_ vssd1 vssd1 vccd1 vccd1 _08411_ sky130_fd_sc_hd__a221o_1
X_11462_ ag2.body\[256\] net789 net764 ag2.body\[260\] _06434_ vssd1 vssd1 vccd1 vccd1
+ _06435_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_22_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17648__B net959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13201_ net287 _07788_ _07789_ net1961 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[368\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_61_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10413_ net742 _05375_ _05382_ _05385_ vssd1 vssd1 vccd1 vccd1 _05386_ sky130_fd_sc_hd__or4_1
X_14181_ net988 _04060_ ag2.body\[198\] net799 vssd1 vssd1 vccd1 vccd1 _08342_ sky130_fd_sc_hd__o22a_1
XANTENNA__11358__A4 _05075_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20617__1560 vssd1 vssd1 vccd1 vccd1 net1560 _20617__1560/LO sky130_fd_sc_hd__conb_1
XFILLER_0_34_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11393_ net1169 control.body\[642\] vssd1 vssd1 vccd1 vccd1 _06366_ sky130_fd_sc_hd__xor2_1
XANTENNA__14353__A net1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18140__A1 net48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10566__A2 net1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_694 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13132_ net291 _07755_ _07756_ net1632 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[332\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_104_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_1348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10344_ ag2.body\[520\] net1231 vssd1 vssd1 vccd1 vccd1 _05317_ sky130_fd_sc_hd__xor2_1
XFILLER_0_123_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_1024 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19637__CLK clknet_leaf_124_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17940_ net345 _03569_ vssd1 vssd1 vccd1 vccd1 _03570_ sky130_fd_sc_hd__nor2_2
XFILLER_0_29_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_13063_ _07725_ net268 _07723_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[295\]
+ sky130_fd_sc_hd__mux2_1
X_10275_ ag2.body\[136\] net1235 vssd1 vssd1 vccd1 vccd1 _05248_ sky130_fd_sc_hd__or2_1
XANTENNA__19920__RESET_B net1368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11515__A1 net504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1400 net1404 vssd1 vssd1 vccd1 vccd1 net1400 sky130_fd_sc_hd__clkbuf_2
X_12014_ _06932_ _06985_ vssd1 vssd1 vccd1 vccd1 _06986_ sky130_fd_sc_hd__nor2_2
XFILLER_0_44_1192 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1411 net1415 vssd1 vssd1 vccd1 vccd1 net1411 sky130_fd_sc_hd__clkbuf_2
XANTENNA__17383__B net942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1422 net1423 vssd1 vssd1 vccd1 vccd1 net1422 sky130_fd_sc_hd__clkbuf_4
X_17871_ img_gen.updater.commands.rR1.rainbowRNG\[11\] img_gen.updater.commands.rR1.rainbowRNG\[10\]
+ _03503_ img_gen.updater.commands.rR1.rainbowRNG\[12\] vssd1 vssd1 vccd1 vccd1 _03515_
+ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_126_4160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14800__B ag2.body\[294\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1433 net1434 vssd1 vssd1 vccd1 vccd1 net1433 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_126_4171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19610_ clknet_leaf_120_clk _00554_ net1394 vssd1 vssd1 vccd1 vccd1 control.body\[776\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout1444 net1452 vssd1 vssd1 vccd1 vccd1 net1444 sky130_fd_sc_hd__clkbuf_4
XANTENNA__16454__B2 net365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16822_ _02497_ _02498_ _02500_ vssd1 vssd1 vccd1 vccd1 _02501_ sky130_fd_sc_hd__and3b_1
XFILLER_0_94_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17651__B1 net928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1455 net1465 vssd1 vssd1 vccd1 vccd1 net1455 sky130_fd_sc_hd__clkbuf_4
Xfanout1466 net1468 vssd1 vssd1 vccd1 vccd1 net1466 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_50_1842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1477 net1478 vssd1 vssd1 vccd1 vccd1 net1477 sky130_fd_sc_hd__buf_2
XANTENNA__12601__A net328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_1853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_122_4035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout490 net492 vssd1 vssd1 vccd1 vccd1 net490 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_6_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18661__CLK clknet_leaf_13_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_122_4046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09533__A_N net1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19787__CLK clknet_leaf_127_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1488 net1489 vssd1 vssd1 vccd1 vccd1 net1488 sky130_fd_sc_hd__buf_2
Xfanout1499 net1504 vssd1 vssd1 vccd1 vccd1 net1499 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_122_4057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_1400 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_19541_ clknet_leaf_118_clk _00485_ net1388 vssd1 vssd1 vccd1 vccd1 control.body\[851\]
+ sky130_fd_sc_hd__dfrtp_1
X_16753_ obsg2.obstacleArray\[40\] net490 net481 obsg2.obstacleArray\[41\] _02431_
+ vssd1 vssd1 vccd1 vccd1 _02432_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_31_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13965_ ag2.body\[104\] net202 _08157_ ag2.body\[96\] vssd1 vssd1 vccd1 vccd1 _00185_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_31_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11818__A2 net545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15704_ ag2.body\[368\] net141 _01629_ ag2.body\[360\] vssd1 vssd1 vccd1 vccd1 _00962_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_88_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11217__A net1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_1526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19472_ clknet_leaf_110_clk _00416_ net1417 vssd1 vssd1 vccd1 vccd1 control.body\[926\]
+ sky130_fd_sc_hd__dfrtp_1
X_12916_ net290 _07654_ _07655_ net1670 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[218\]
+ sky130_fd_sc_hd__a22o_1
X_16684_ net358 _02256_ _02260_ _02211_ vssd1 vssd1 vccd1 vccd1 _02363_ sky130_fd_sc_hd__a31o_1
XANTENNA__10121__A net1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13896_ ag2.body\[43\] net118 _08149_ ag2.body\[35\] vssd1 vssd1 vccd1 vccd1 _00124_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__16727__B net957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output26_A net26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18423_ _03811_ _03911_ vssd1 vssd1 vccd1 vccd1 _03912_ sky130_fd_sc_hd__nand2_1
X_15635_ ag2.body\[434\] net125 _01622_ ag2.body\[426\] vssd1 vssd1 vccd1 vccd1 _00900_
+ sky130_fd_sc_hd__a22o_1
X_12847_ _07431_ _07624_ vssd1 vssd1 vccd1 vccd1 _07625_ sky130_fd_sc_hd__nor2_1
XANTENNA__14528__A net1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_135_4429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18354_ _04402_ _07181_ _03849_ vssd1 vssd1 vccd1 vccd1 _03850_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_48_1793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15566_ ag2.body\[501\] net185 _01614_ ag2.body\[493\] vssd1 vssd1 vccd1 vccd1 _00839_
+ sky130_fd_sc_hd__a22o_1
X_12778_ _06672_ _07310_ vssd1 vssd1 vccd1 vccd1 _07592_ sky130_fd_sc_hd__or2_2
XTAP_TAPCELL_ROW_44_1657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10775__B net1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17305_ ag2.body\[394\] net862 vssd1 vssd1 vccd1 vccd1 _02984_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_51_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14517_ net1024 ag2.body\[318\] vssd1 vssd1 vccd1 vccd1 _08678_ sky130_fd_sc_hd__xor2_1
XFILLER_0_12_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18285_ net517 _03781_ vssd1 vssd1 vccd1 vccd1 _01390_ sky130_fd_sc_hd__nor2_1
XFILLER_0_72_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_44_1679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11729_ img_gen.tracker.frame\[209\] net608 net552 img_gen.tracker.frame\[212\] vssd1
+ vssd1 vccd1 vccd1 _06701_ sky130_fd_sc_hd__o22a_1
XFILLER_0_9_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15497_ _06290_ net54 vssd1 vssd1 vccd1 vccd1 _01607_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_25_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19167__CLK clknet_leaf_52_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_365 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17236_ ag2.body\[441\] net732 net960 _04158_ _02909_ vssd1 vssd1 vccd1 vccd1 _02915_
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_117_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_14448_ net846 ag2.body\[224\] ag2.body\[230\] net804 _08608_ vssd1 vssd1 vccd1 vccd1
+ _08609_ sky130_fd_sc_hd__a221o_1
XFILLER_0_128_1525 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17558__B net855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_94_3182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_981 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_17167_ ag2.body\[593\] net730 net715 ag2.body\[595\] vssd1 vssd1 vccd1 vccd1 _02846_
+ sky130_fd_sc_hd__a22o_1
X_14379_ _08535_ _08536_ _08537_ _08533_ vssd1 vssd1 vccd1 vccd1 _08540_ sky130_fd_sc_hd__a211o_1
XANTENNA__14263__A net989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_94_3193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold905 img_gen.updater.commands.rR1.rainbowRNG\[2\] vssd1 vssd1 vccd1 vccd1 net2467
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_1524 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold916 ag2.body\[584\] vssd1 vssd1 vccd1 vccd1 net2478 sky130_fd_sc_hd__dlygate4sd3_1
Xhold927 sound_gen.osc1.freq\[2\] vssd1 vssd1 vccd1 vccd1 net2489 sky130_fd_sc_hd__dlygate4sd3_1
X_16118_ _01795_ _01796_ net377 vssd1 vssd1 vccd1 vccd1 _01797_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_90_3057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold938 control.body\[640\] vssd1 vssd1 vccd1 vccd1 net2500 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_51_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_1568 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold949 ag2.body\[460\] vssd1 vssd1 vccd1 vccd1 net2511 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_90_3068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17098_ ag2.body\[298\] net726 net719 ag2.body\[299\] vssd1 vssd1 vccd1 vccd1 _02777_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_90_3079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08940_ net994 vssd1 vssd1 vccd1 vccd1 _03965_ sky130_fd_sc_hd__inv_2
XFILLER_0_110_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16049_ net460 _01727_ vssd1 vssd1 vccd1 vccd1 _01728_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_102_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17293__B net865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20294__CLK clknet_leaf_37_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10015__B net1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17642__B1 net695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19808_ clknet_leaf_125_clk _00752_ net1410 vssd1 vssd1 vccd1 vccd1 ag2.body\[590\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_58_1317 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_1590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_105_3521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_105_3532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19739_ clknet_leaf_129_clk _00683_ net1325 vssd1 vssd1 vccd1 vccd1 control.body\[649\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_56_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_101_3407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_101_3418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16748__A2 net501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09883__B1 net1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09423_ obsg2.obsNeeded\[0\] net516 vssd1 vssd1 vccd1 vccd1 _04401_ sky130_fd_sc_hd__or2_1
XFILLER_0_133_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14759__A1 net817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14759__B2 net1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10966__A net1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout347_A _01732_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14438__A net1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09354_ _04355_ vssd1 vssd1 vccd1 vccd1 _04356_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout1089_A net1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_118_3915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10685__B net1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_118_3926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_118_3937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_60_2160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_1413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15708__B1 _01629_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09285_ _04303_ _04304_ vssd1 vssd1 vccd1 vccd1 sound_gen.osc1.keepCounting_nxt sky130_fd_sc_hd__nor2_1
XFILLER_0_129_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout514_A net515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_1573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout135_X net135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20514_ clknet_leaf_113_clk net324 net1401 vssd1 vssd1 vccd1 vccd1 track.highScore\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09819__X _04792_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_596 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16920__A2 net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_324 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_1711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20445_ clknet_leaf_42_clk _01332_ net1373 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[81\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA_fanout1423_A net1435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11745__A1 net565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20376_ clknet_leaf_25_clk _01263_ net1344 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[12\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_63_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout883_A net884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16799__S net402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_2543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_1322 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_2554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16684__A1 net358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout1211_X net1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13498__A1 net250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10206__A net1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10060_ ag2.body\[483\] net768 net1057 _04177_ vssd1 vssd1 vccd1 vccd1 _05033_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout671_X net671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout769_X net769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10720__A2 net774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_2948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17931__B _03562_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_2959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout936_X net936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12140__B net599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_67_2358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10962_ _05927_ _05932_ _05933_ _05934_ vssd1 vssd1 vccd1 vccd1 _05935_ sky130_fd_sc_hd__or4_2
X_13750_ _08068_ vssd1 vssd1 vccd1 vccd1 _08069_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_67_2369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16739__A2 net491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout48_X net48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12701_ net283 net310 _07553_ _07554_ net1595 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[104\]
+ sky130_fd_sc_hd__a32o_1
XANTENNA__11681__B1 net601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10893_ net1047 control.body\[655\] vssd1 vssd1 vccd1 vccd1 _05866_ sky130_fd_sc_hd__xor2_1
X_13681_ net905 net639 vssd1 vssd1 vccd1 vccd1 _08026_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_38_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13252__A _06724_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15420_ control.body\[627\] net83 _01598_ ag2.body\[619\] vssd1 vssd1 vccd1 vccd1
+ _00709_ sky130_fd_sc_hd__a22o_1
X_12632_ net621 net436 net468 net574 vssd1 vssd1 vccd1 vccd1 _07518_ sky130_fd_sc_hd__or4_1
XFILLER_0_66_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13422__A1 net236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14067__B ag2.body\[209\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_1513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15351_ net2225 net72 _01591_ control.body\[685\] vssd1 vssd1 vccd1 vccd1 _00647_
+ sky130_fd_sc_hd__a22o_1
X_12563_ net678 _07481_ vssd1 vssd1 vccd1 vccd1 _07482_ sky130_fd_sc_hd__nor2_1
XFILLER_0_31_39 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__16563__A net350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11514_ obsg2.obstacleArray\[115\] net633 net509 obsg2.obstacleArray\[119\] net506
+ vssd1 vssd1 vccd1 vccd1 _06487_ sky130_fd_sc_hd__o221a_1
XANTENNA__11039__A_N net1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14302_ net838 ag2.body\[217\] ag2.body\[221\] net808 _08460_ vssd1 vssd1 vccd1 vccd1
+ _08463_ sky130_fd_sc_hd__a221o_1
XFILLER_0_110_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18070_ net42 _03662_ vssd1 vssd1 vccd1 vccd1 _03663_ sky130_fd_sc_hd__nor2_1
XFILLER_0_53_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12494_ net1658 _07441_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[10\]
+ sky130_fd_sc_hd__and2_1
X_15282_ _04606_ net55 vssd1 vssd1 vccd1 vccd1 _01584_ sky130_fd_sc_hd__nor2_2
XFILLER_0_48_1519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16911__A2 net869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17021_ ag2.body\[334\] net945 vssd1 vssd1 vccd1 vccd1 _02700_ sky130_fd_sc_hd__xor2_1
XFILLER_0_22_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18551__Q ag2.y\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14233_ net1025 ag2.body\[485\] vssd1 vssd1 vccd1 vccd1 _08394_ sky130_fd_sc_hd__nand2_1
X_11445_ net1134 control.body\[956\] vssd1 vssd1 vccd1 vccd1 _06418_ sky130_fd_sc_hd__nand2_1
XFILLER_0_62_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11500__A net1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14164_ net971 ag2.body\[203\] vssd1 vssd1 vccd1 vccd1 _08325_ sky130_fd_sc_hd__xor2_1
X_11376_ _04168_ net1197 net1080 _04171_ _06348_ vssd1 vssd1 vccd1 vccd1 _06349_ sky130_fd_sc_hd__a221o_1
XFILLER_0_21_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_128_4222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10327_ _05288_ _05289_ _05294_ _05299_ vssd1 vssd1 vccd1 vccd1 _05300_ sky130_fd_sc_hd__or4_2
X_13115_ net339 net285 net329 _07471_ _07749_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[323\]
+ sky130_fd_sc_hd__a41o_1
XTAP_TAPCELL_ROW_128_4233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14095_ net992 ag2.body\[281\] vssd1 vssd1 vccd1 vccd1 _08256_ sky130_fd_sc_hd__xnor2_1
X_18972_ clknet_leaf_7_clk img_gen.tracker.next_frame\[410\] net1265 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[410\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_123_1455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14811__A net1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10116__A net1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1541 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_1450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17923_ net516 _03556_ vssd1 vssd1 vccd1 vccd1 _01253_ sky130_fd_sc_hd__nor2_1
X_13046_ img_gen.tracker.frame\[287\] net646 _07716_ vssd1 vssd1 vccd1 vccd1 _07717_
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_37_1461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_124_4108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_1488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10258_ net767 control.body\[787\] _05226_ _05227_ _05230_ vssd1 vssd1 vccd1 vccd1
+ _05231_ sky130_fd_sc_hd__o2111a_1
XTAP_TAPCELL_ROW_124_4119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout1230 net1232 vssd1 vssd1 vccd1 vccd1 net1230 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_33_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout1241 net1242 vssd1 vssd1 vccd1 vccd1 net1241 sky130_fd_sc_hd__clkbuf_4
X_17854_ _07304_ _07316_ img_gen.updater.commands.rR1.rainbowRNG\[1\] img_gen.updater.commands.rR1.rainbowRNG\[0\]
+ vssd1 vssd1 vccd1 vccd1 _03509_ sky130_fd_sc_hd__o211a_1
Xfanout1252 net1254 vssd1 vssd1 vccd1 vccd1 net1252 sky130_fd_sc_hd__buf_2
X_10189_ net641 _04432_ vssd1 vssd1 vccd1 vccd1 _05162_ sky130_fd_sc_hd__nor2_2
Xfanout1263 net1333 vssd1 vssd1 vccd1 vccd1 net1263 sky130_fd_sc_hd__buf_2
XFILLER_0_59_1637 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xfanout1274 net1275 vssd1 vssd1 vccd1 vccd1 net1274 sky130_fd_sc_hd__clkbuf_4
XANTENNA__20321__Q obsg2.randCord\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16805_ _03999_ net877 net945 _04001_ _02483_ vssd1 vssd1 vccd1 vccd1 _02484_ sky130_fd_sc_hd__a221o_1
Xfanout1285 net1286 vssd1 vssd1 vccd1 vccd1 net1285 sky130_fd_sc_hd__clkbuf_4
Xfanout1296 net1311 vssd1 vssd1 vccd1 vccd1 net1296 sky130_fd_sc_hd__buf_2
X_17785_ _03460_ _03462_ net1036 vssd1 vssd1 vccd1 vccd1 _01210_ sky130_fd_sc_hd__mux2_1
X_14997_ control.body\[1003\] net151 _01551_ net2214 vssd1 vssd1 vccd1 vccd1 _00333_
+ sky130_fd_sc_hd__a22o_1
X_19524_ clknet_leaf_121_clk _00468_ net1401 vssd1 vssd1 vccd1 vccd1 control.body\[866\]
+ sky130_fd_sc_hd__dfrtp_1
X_16736_ obsg2.obstacleArray\[55\] net501 net491 obsg2.obstacleArray\[52\] vssd1 vssd1
+ vccd1 vccd1 _02415_ sky130_fd_sc_hd__a22o_1
X_13948_ ag2.body\[89\] net190 _08155_ ag2.body\[81\] vssd1 vssd1 vccd1 vccd1 _00170_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_89_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17927__A1 net318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12985__B net333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19455_ clknet_leaf_110_clk _00399_ net1422 vssd1 vssd1 vccd1 vccd1 control.body\[941\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_46_1719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16667_ obsg2.obstacleArray\[18\] net448 vssd1 vssd1 vccd1 vccd1 _02346_ sky130_fd_sc_hd__or2_1
X_13879_ ag2.body\[28\] net115 _08147_ ag2.body\[20\] vssd1 vssd1 vccd1 vccd1 _00109_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__10786__A net1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18406_ _03835_ _03894_ _03895_ _03891_ vssd1 vssd1 vccd1 vccd1 _03896_ sky130_fd_sc_hd__a31o_1
XFILLER_0_53_1269 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_1595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15618_ ag2.body\[451\] net127 _01613_ ag2.body\[443\] vssd1 vssd1 vccd1 vccd1 _00885_
+ sky130_fd_sc_hd__a22o_1
X_19386_ clknet_leaf_112_clk _00330_ net1425 vssd1 vssd1 vccd1 vccd1 control.body\[1000\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_1681 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13413__A1 net257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16598_ net395 _02276_ _02275_ net359 vssd1 vssd1 vccd1 vccd1 _02277_ sky130_fd_sc_hd__a211o_1
XANTENNA__18557__CLK clknet_leaf_43_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18337_ _04644_ _08025_ _03831_ vssd1 vssd1 vccd1 vccd1 _03833_ sky130_fd_sc_hd__o21a_1
XFILLER_0_17_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15549_ ag2.body\[519\] net188 _01580_ ag2.body\[511\] vssd1 vssd1 vccd1 vccd1 _00825_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_96_3244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17155__A2 net722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_41 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_96_3255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_1589 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_96_3266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_1023 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09070_ ag2.body\[279\] vssd1 vssd1 vccd1 vccd1 _04095_ sky130_fd_sc_hd__inv_2
X_18268_ net319 _03559_ obsg2.obstacleArray\[131\] vssd1 vssd1 vccd1 vccd1 _03773_
+ sky130_fd_sc_hd__a21oi_1
XANTENNA__17288__B net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_92_3119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_85 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17219_ ag2.body\[315\] net720 net707 ag2.body\[317\] vssd1 vssd1 vccd1 vccd1 _02898_
+ sky130_fd_sc_hd__a22o_1
X_18199_ obsg2.obstacleArray\[96\] _03738_ net521 vssd1 vssd1 vccd1 vccd1 _01347_
+ sky130_fd_sc_hd__o21a_1
XANTENNA__12506__A net387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold702 control.body\[912\] vssd1 vssd1 vccd1 vccd1 net2264 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_1452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20230_ clknet_leaf_66_clk _01174_ net1476 vssd1 vssd1 vccd1 vccd1 ag2.body\[164\]
+ sky130_fd_sc_hd__dfrtp_4
Xhold713 control.body\[1092\] vssd1 vssd1 vccd1 vccd1 net2275 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__16115__B1 _01729_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold724 control.body\[842\] vssd1 vssd1 vccd1 vccd1 net2286 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_4_1__f_clk_A clknet_3_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold735 control.body\[790\] vssd1 vssd1 vccd1 vccd1 net2297 sky130_fd_sc_hd__dlygate4sd3_1
Xhold746 control.body\[726\] vssd1 vssd1 vccd1 vccd1 net2308 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_64_1365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16666__A1 net396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold757 control.body\[1059\] vssd1 vssd1 vccd1 vccd1 net2319 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1653 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold768 control.body\[927\] vssd1 vssd1 vccd1 vccd1 net2330 sky130_fd_sc_hd__dlygate4sd3_1
X_20161_ clknet_leaf_96_clk _01105_ net1441 vssd1 vssd1 vccd1 vccd1 ag2.body\[239\]
+ sky130_fd_sc_hd__dfrtp_4
XPHY_EDGE_ROW_123_Right_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold779 control.body\[806\] vssd1 vssd1 vccd1 vccd1 net2341 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09972_ net639 _04427_ net899 vssd1 vssd1 vccd1 vccd1 _04945_ sky130_fd_sc_hd__a21o_1
XANTENNA__10928__A1_N net761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_1539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20092_ clknet_leaf_78_clk _01036_ net1490 vssd1 vssd1 vccd1 vccd1 ag2.body\[298\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_41_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13337__A net332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10313__X _05286_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1004_A net1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16969__A2 net724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20231__Q ag2.body\[165\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13056__B net660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_311 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout464_A net465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19332__CLK clknet_leaf_103_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_2801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09550__A net1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_2200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_2211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout252_X net252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_2222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout1373_A net1374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout729_A _04264_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13072__A net685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09406_ sound_gen.osc1.keepCounting_nxt _04304_ net2329 vssd1 vssd1 vccd1 vccd1 _01399_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_93 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__13404__A1 net284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_1679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13955__A2 net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09337_ sound_gen.at_max net1589 vssd1 vssd1 vccd1 vccd1 _01427_ sky130_fd_sc_hd__xor2_1
XFILLER_0_8_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout1161_X net1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16383__A net538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11966__A1 net560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_2730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_1443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09549__X _04522_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_2741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09268_ sound_gen.osc1.timer\[1\] sound_gen.osc1.timer\[2\] _04284_ _04285_ vssd1
+ vssd1 vccd1 vccd1 _04291_ sky130_fd_sc_hd__nor4_1
XFILLER_0_35_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_302 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__17198__B net861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14615__B ag2.body\[57\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_2605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_75_2616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_1287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09709__B net1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09199_ ag2.body\[620\] vssd1 vssd1 vccd1 vccd1 _04224_ sky130_fd_sc_hd__inv_2
XFILLER_0_69_1298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_2026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11230_ net1076 control.body\[862\] vssd1 vssd1 vccd1 vccd1 _06203_ sky130_fd_sc_hd__nand2_1
X_20428_ clknet_4_6__leaf_clk _01315_ net1370 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleArray\[64\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_56_2037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout886_X net886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11161_ ag2.body\[601\] net1196 vssd1 vssd1 vccd1 vccd1 _06134_ sky130_fd_sc_hd__nand2_1
X_20359_ clknet_leaf_22_clk _01250_ net1361 vssd1 vssd1 vccd1 vccd1 obsg2.obstacleCount\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__20417__RESET_B net1357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10112_ _05077_ _05078_ _05083_ _05084_ vssd1 vssd1 vccd1 vccd1 _05085_ sky130_fd_sc_hd__a22o_1
XANTENNA__09725__A _04695_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11092_ _06041_ _06047_ _06050_ net476 _05303_ vssd1 vssd1 vccd1 vccd1 _06065_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_8_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11974__B net550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10043_ net1202 control.body\[897\] vssd1 vssd1 vccd1 vccd1 _05016_ sky130_fd_sc_hd__xor2_1
X_14920_ control.body\[1079\] net171 _01542_ control.body\[1071\] vssd1 vssd1 vccd1
+ vccd1 _00265_ sky130_fd_sc_hd__a22o_1
XANTENNA__15880__A2 net192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09444__B net899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold40 ag2.body\[1\] vssd1 vssd1 vccd1 vccd1 net1602 sky130_fd_sc_hd__dlygate4sd3_1
Xhold51 img_gen.tracker.frame\[519\] vssd1 vssd1 vccd1 vccd1 net1613 sky130_fd_sc_hd__dlygate4sd3_1
Xhold62 img_gen.tracker.frame\[103\] vssd1 vssd1 vccd1 vccd1 net1624 sky130_fd_sc_hd__dlygate4sd3_1
Xhold73 img_gen.tracker.frame\[164\] vssd1 vssd1 vccd1 vccd1 net1635 sky130_fd_sc_hd__dlygate4sd3_1
X_14851_ _08509_ _08584_ _08683_ _08699_ vssd1 vssd1 vccd1 vccd1 _01522_ sky130_fd_sc_hd__and4_2
XFILLER_0_76_1247 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xhold84 img_gen.tracker.frame\[485\] vssd1 vssd1 vccd1 vccd1 net1646 sky130_fd_sc_hd__dlygate4sd3_1
Xhold95 img_gen.tracker.frame\[517\] vssd1 vssd1 vccd1 vccd1 net1657 sky130_fd_sc_hd__dlygate4sd3_1
X_13802_ _08104_ _08105_ net1217 vssd1 vssd1 vccd1 vccd1 _00074_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17570_ ag2.body\[582\] net938 vssd1 vssd1 vccd1 vccd1 _03249_ sky130_fd_sc_hd__xor2_1
XFILLER_0_98_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14782_ net838 ag2.body\[273\] ag2.body\[274\] net828 _01446_ vssd1 vssd1 vccd1 vccd1
+ _01453_ sky130_fd_sc_hd__a221o_1
X_11994_ img_gen.tracker.frame\[412\] net600 net584 img_gen.tracker.frame\[418\] _06965_
+ vssd1 vssd1 vccd1 vccd1 _06966_ sky130_fd_sc_hd__o221a_1
XANTENNA__16277__B net412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18031__B1 net531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16521_ _02181_ _02198_ _02086_ vssd1 vssd1 vccd1 vccd1 _02200_ sky130_fd_sc_hd__a21oi_1
XANTENNA_clkbuf_4_12__f_clk_A clknet_3_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09460__A net894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13733_ _04391_ _07228_ _08056_ _08055_ vssd1 vssd1 vccd1 vccd1 _00054_ sky130_fd_sc_hd__o31a_1
X_10945_ _05913_ _05915_ _05916_ _05917_ vssd1 vssd1 vccd1 vccd1 _05918_ sky130_fd_sc_hd__or4_1
XFILLER_0_58_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14078__A net971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19825__CLK clknet_leaf_124_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19240_ clknet_leaf_84_clk _00184_ net1481 vssd1 vssd1 vccd1 vccd1 ag2.body\[103\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_42_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16452_ net402 _02130_ net367 vssd1 vssd1 vccd1 vccd1 _02131_ sky130_fd_sc_hd__o21a_1
X_13664_ net972 _08014_ vssd1 vssd1 vccd1 vccd1 _08018_ sky130_fd_sc_hd__nand2_1
XFILLER_0_128_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10876_ _05845_ _05846_ _05847_ _05848_ vssd1 vssd1 vccd1 vccd1 _05849_ sky130_fd_sc_hd__a22o_1
X_15403_ control.body\[644\] net83 _01581_ net2424 vssd1 vssd1 vccd1 vccd1 _00694_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_54_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19171_ clknet_leaf_53_clk _00115_ net1366 vssd1 vssd1 vccd1 vccd1 ag2.body\[34\]
+ sky130_fd_sc_hd__dfrtp_4
X_12615_ net666 _07509_ vssd1 vssd1 vccd1 vccd1 _07510_ sky130_fd_sc_hd__nor2_1
X_16383_ net538 _02058_ vssd1 vssd1 vccd1 vccd1 _02062_ sky130_fd_sc_hd__nand2_1
XANTENNA__14228__D net1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13595_ control.divider.count\[14\] _07953_ control.divider.count\[12\] _03960_ vssd1
+ vssd1 vccd1 vccd1 _07970_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_53_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18122_ net46 _03696_ vssd1 vssd1 vccd1 vccd1 _03697_ sky130_fd_sc_hd__nor2_1
XFILLER_0_93_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_1343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15334_ control.body\[710\] net73 _01587_ net2265 vssd1 vssd1 vccd1 vccd1 _00632_
+ sky130_fd_sc_hd__a22o_1
X_12546_ net594 net436 net473 net561 vssd1 vssd1 vccd1 vccd1 _07471_ sky130_fd_sc_hd__and4_1
XFILLER_0_87_1376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16440__S0 net454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17676__X _03355_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18053_ net522 _03651_ vssd1 vssd1 vccd1 vccd1 _01288_ sky130_fd_sc_hd__and2_1
XANTENNA__16896__B2 ag2.body\[213\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15265_ net2549 net109 _01582_ control.body\[752\] vssd1 vssd1 vccd1 vccd1 _00570_
+ sky130_fd_sc_hd__a22o_1
X_12477_ _07425_ _07430_ net678 vssd1 vssd1 vccd1 vccd1 _07432_ sky130_fd_sc_hd__a21oi_1
X_17004_ _02678_ _02680_ _02682_ vssd1 vssd1 vccd1 vccd1 _02683_ sky130_fd_sc_hd__or3b_1
XANTENNA_4 _03230_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11230__A net1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20316__Q ag2.randCord\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14216_ net801 ag2.body\[414\] ag2.body\[415\] net793 _08376_ vssd1 vssd1 vccd1 vccd1
+ _08377_ sky130_fd_sc_hd__o221a_1
XFILLER_0_112_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_39_1512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11428_ ag2.body\[399\] net1056 vssd1 vssd1 vccd1 vccd1 _06401_ sky130_fd_sc_hd__or2_1
X_15196_ net2461 net95 _01573_ control.body\[820\] vssd1 vssd1 vccd1 vccd1 _00510_
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_39_1523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11185__A2 net784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11359_ net773 control.body\[810\] _04243_ net1049 vssd1 vssd1 vccd1 vccd1 _06332_
+ sky130_fd_sc_hd__o22a_1
X_14147_ net1015 ag2.body\[598\] vssd1 vssd1 vccd1 vccd1 _08308_ sky130_fd_sc_hd__xnor2_1
XANTENNA__12613__X _07508_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14541__A net1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18013__A net432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_57 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18955_ clknet_leaf_5_clk img_gen.tracker.next_frame\[393\] net1269 vssd1 vssd1 vccd1
+ vccd1 img_gen.tracker.frame\[393\] sky130_fd_sc_hd__dfrtp_1
X_14078_ net971 ag2.body\[563\] vssd1 vssd1 vccd1 vccd1 _08239_ sky130_fd_sc_hd__xor2_1
XFILLER_0_123_1296 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_60_Left_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17906_ _03533_ _03538_ vssd1 vssd1 vccd1 vccd1 _03541_ sky130_fd_sc_hd__or2_1
X_13029_ net259 _07708_ _07709_ net1970 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[277\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_59_1401 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18886_ clknet_leaf_26_clk img_gen.tracker.next_frame\[324\] net1339 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[324\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__15075__C net65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20051__Q ag2.body\[337\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1060 net1062 vssd1 vssd1 vccd1 vccd1 net1060 sky130_fd_sc_hd__clkbuf_4
Xfanout1071 net1072 vssd1 vssd1 vccd1 vccd1 net1071 sky130_fd_sc_hd__clkbuf_2
X_17837_ net662 _03495_ vssd1 vssd1 vccd1 vccd1 _01228_ sky130_fd_sc_hd__and2_1
XANTENNA_clkbuf_leaf_6_clk_A clknet_4_1__leaf_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1082 ag2.x\[2\] vssd1 vssd1 vccd1 vccd1 net1082 sky130_fd_sc_hd__clkbuf_4
XANTENNA__17571__B net879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout1093 ag2.x\[2\] vssd1 vssd1 vccd1 vccd1 net1093 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_59_1467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17768_ _02566_ _02755_ _02768_ _03140_ vssd1 vssd1 vccd1 vccd1 _03447_ sky130_fd_sc_hd__and4_1
XANTENNA__20332__CLK clknet_leaf_20_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_141 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__14831__B1 _01500_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16719_ obsg2.obstacleArray\[107\] net501 net487 obsg2.obstacleArray\[106\] vssd1
+ vssd1 vccd1 vccd1 _02398_ sky130_fd_sc_hd__a22o_1
XFILLER_0_72_1645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19507_ clknet_leaf_113_clk _00451_ net1396 vssd1 vssd1 vccd1 vccd1 control.body\[881\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_92_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17699_ obsg2.obstacleArray\[128\] obsg2.obstacleArray\[129\] obsg2.obstacleArray\[132\]
+ obsg2.obstacleArray\[133\] net410 net370 vssd1 vssd1 vccd1 vccd1 _03378_ sky130_fd_sc_hd__mux4_1
XFILLER_0_92_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_18_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_98_3306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_1689 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19438_ clknet_leaf_110_clk net2280 net1422 vssd1 vssd1 vccd1 vccd1 control.body\[956\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_98_3317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_1245 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16915__B net881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19369_ clknet_leaf_102_clk _00313_ net1438 vssd1 vssd1 vccd1 vccd1 control.body\[1031\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_72_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09122_ ag2.body\[407\] vssd1 vssd1 vccd1 vccd1 _04147_ sky130_fd_sc_hd__inv_2
XFILLER_0_130_1289 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1405 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_121 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_09053_ ag2.body\[247\] vssd1 vssd1 vccd1 vccd1 _04078_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_3 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkload100_A clknet_leaf_98_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16351__A3 _01996_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20226__Q ag2.body\[160\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_165 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold510 img_gen.tracker.frame\[241\] vssd1 vssd1 vccd1 vccd1 net2072 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold521 control.divider.count\[7\] vssd1 vssd1 vccd1 vccd1 net2083 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16650__B net446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17836__A0 net1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold532 _00419_ vssd1 vssd1 vccd1 vccd1 net2094 sky130_fd_sc_hd__dlygate4sd3_1
X_20213_ clknet_leaf_60_clk _01157_ net1466 vssd1 vssd1 vccd1 vccd1 ag2.body\[179\]
+ sky130_fd_sc_hd__dfrtp_4
Xhold543 img_gen.tracker.frame\[34\] vssd1 vssd1 vccd1 vccd1 net2105 sky130_fd_sc_hd__dlygate4sd3_1
Xhold554 img_gen.tracker.frame\[565\] vssd1 vssd1 vccd1 vccd1 net2116 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold565 img_gen.tracker.frame\[321\] vssd1 vssd1 vccd1 vccd1 net2127 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1121_A net1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold576 img_gen.tracker.frame\[75\] vssd1 vssd1 vccd1 vccd1 net2138 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__20510__RESET_B net1403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold587 img_gen.tracker.frame\[464\] vssd1 vssd1 vccd1 vccd1 net2149 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout1219_A net1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold598 control.divider.next_count\[1\] vssd1 vssd1 vccd1 vccd1 net2160 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_1314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20144_ clknet_leaf_97_clk _01088_ net1449 vssd1 vssd1 vccd1 vccd1 ag2.body\[254\]
+ sky130_fd_sc_hd__dfrtp_4
X_09955_ net783 control.body\[736\] control.body\[737\] net777 vssd1 vssd1 vccd1 vccd1
+ _04928_ sky130_fd_sc_hd__a22o_1
XFILLER_0_99_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout581_A net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout679_A net681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20075_ clknet_leaf_77_clk _01019_ net1491 vssd1 vssd1 vccd1 vccd1 ag2.body\[313\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__13873__A1 _07181_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09886_ _04446_ _04632_ vssd1 vssd1 vccd1 vccd1 _04859_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout1007_X net1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16498__S0 net458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17481__B net887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout846_A net847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout1490_A net1492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18722__CLK clknet_leaf_142_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout467_X net467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16811__A1 ag2.body\[66\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1578 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19848__CLK clknet_leaf_93_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15282__A _04606_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16811__B2 ag2.body\[67\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10697__Y _05670_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11636__B1 _06497_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13514__B _07807_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout634_X net634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_0_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10730_ ag2.body\[249\] net779 _05699_ _05700_ _05702_ vssd1 vssd1 vccd1 vccd1 _05703_
+ sky130_fd_sc_hd__a221o_1
XANTENNA__16575__B1 net391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18872__CLK clknet_leaf_22_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17772__C1 _02622_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16825__B net854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_177 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_10661_ net921 _04431_ _05051_ _05633_ vssd1 vssd1 vccd1 vccd1 _05634_ sky130_fd_sc_hd__o31a_1
XANTENNA_fanout801_X net801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14626__A net1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12400_ img_gen.updater.commands.rR1.rainbowRNG\[11\] _07319_ _07320_ _07360_ _07363_
+ vssd1 vssd1 vccd1 vccd1 _07364_ sky130_fd_sc_hd__a221o_1
XANTENNA__12061__B1 net609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13380_ net249 _07864_ _07865_ net1904 vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[472\]
+ sky130_fd_sc_hd__a22o_1
X_10592_ net1149 control.body\[827\] vssd1 vssd1 vccd1 vccd1 _05565_ sky130_fd_sc_hd__xor2_1
XFILLER_0_63_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19197__Q ag2.body\[60\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10873__B net1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_1625 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__19228__CLK clknet_leaf_75_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12331_ _07295_ _07297_ vssd1 vssd1 vccd1 vccd1 _07298_ sky130_fd_sc_hd__or2_1
XANTENNA__09439__B net1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10218__X _05191_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12262_ img_gen.updater.commands.mode\[2\] img_gen.updater.commands.mode\[0\] img_gen.updater.commands.mode\[1\]
+ vssd1 vssd1 vccd1 vccd1 _07232_ sky130_fd_sc_hd__or3b_2
X_15050_ net2519 net163 _01558_ control.body\[945\] vssd1 vssd1 vccd1 vccd1 _00379_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_133_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17656__B net934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15550__A1 _04416_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14001_ net844 ag2.body\[504\] ag2.body\[508\] net814 vssd1 vssd1 vccd1 vccd1 _08162_
+ sky130_fd_sc_hd__o22a_1
X_11213_ net1171 control.body\[842\] vssd1 vssd1 vccd1 vccd1 _06186_ sky130_fd_sc_hd__xnor2_1
X_12193_ _07153_ _07154_ _07161_ _07162_ vssd1 vssd1 vccd1 vccd1 _07165_ sky130_fd_sc_hd__a22o_1
Xoutput30 net30 vssd1 vssd1 vccd1 vccd1 gpio_out[5] sky130_fd_sc_hd__buf_2
XANTENNA__14361__A net1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11572__C1 net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11144_ ag2.body\[415\] net1056 vssd1 vssd1 vccd1 vccd1 _06117_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09455__A net901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_29 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_18740_ clknet_leaf_142_clk img_gen.tracker.next_frame\[178\] net1261 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[178\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_27 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_15952_ ag2.body\[157\] net199 _01656_ ag2.body\[149\] vssd1 vssd1 vccd1 vccd1 _01183_
+ sky130_fd_sc_hd__a22o_1
X_11075_ ag2.body\[364\] net763 net757 ag2.body\[365\] _06044_ vssd1 vssd1 vccd1 vccd1
+ _06048_ sky130_fd_sc_hd__o221a_1
X_14903_ net895 _05980_ net66 vssd1 vssd1 vccd1 vccd1 _01541_ sky130_fd_sc_hd__and3_2
X_10026_ ag2.body\[506\] net1184 vssd1 vssd1 vccd1 vccd1 _04999_ sky130_fd_sc_hd__nand2_1
XANTENNA__11875__B1 net582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18671_ clknet_leaf_27_clk img_gen.tracker.next_frame\[109\] net1339 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[109\] sky130_fd_sc_hd__dfrtp_1
X_15883_ _04539_ net67 vssd1 vssd1 vccd1 vccd1 _01649_ sky130_fd_sc_hd__and2_2
X_17622_ ag2.body\[186\] net724 net697 ag2.body\[190\] _03300_ vssd1 vssd1 vccd1 vccd1
+ _03301_ sky130_fd_sc_hd__o221a_1
XFILLER_0_99_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14834_ _08236_ _08246_ _08378_ _08457_ vssd1 vssd1 vccd1 vccd1 _01505_ sky130_fd_sc_hd__and4_1
XFILLER_0_53_15 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17553_ ag2.body\[357\] net953 vssd1 vssd1 vccd1 vccd1 _03232_ sky130_fd_sc_hd__xor2_1
XANTENNA__11627__B1 net475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14765_ net984 ag2.body\[98\] vssd1 vssd1 vccd1 vccd1 _08926_ sky130_fd_sc_hd__xor2_1
XFILLER_0_15_1304 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_11977_ img_gen.tracker.frame\[553\] net622 net549 img_gen.tracker.frame\[559\] vssd1
+ vssd1 vccd1 vccd1 _06949_ sky130_fd_sc_hd__o22a_1
XFILLER_0_118_1398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16504_ obsg2.obstacleArray\[0\] obsg2.obstacleArray\[1\] net457 vssd1 vssd1 vccd1
+ vccd1 _02183_ sky130_fd_sc_hd__mux2_1
XANTENNA__11225__A net1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15920__A _05921_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13716_ track.highScore\[5\] _08027_ net356 vssd1 vssd1 vccd1 vccd1 track.nextHighScore\[5\]
+ sky130_fd_sc_hd__mux2_1
X_17484_ _03152_ _03153_ _03159_ _03160_ vssd1 vssd1 vccd1 vccd1 _03163_ sky130_fd_sc_hd__a22o_1
X_10928_ net761 control.body\[1036\] control.body\[1038\] net750 vssd1 vssd1 vccd1
+ vccd1 _05901_ sky130_fd_sc_hd__a2bb2o_1
X_14696_ net1033 ag2.body\[325\] vssd1 vssd1 vccd1 vccd1 _08857_ sky130_fd_sc_hd__xnor2_1
X_19223_ clknet_leaf_67_clk _00167_ net1494 vssd1 vssd1 vccd1 vccd1 ag2.body\[86\]
+ sky130_fd_sc_hd__dfrtp_4
X_16435_ net401 _02113_ _02112_ net366 vssd1 vssd1 vccd1 vccd1 _02114_ sky130_fd_sc_hd__a211o_1
X_13647_ _08005_ vssd1 vssd1 vccd1 vccd1 _08006_ sky130_fd_sc_hd__inv_2
XFILLER_0_32_1651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10859_ net1193 control.body\[689\] vssd1 vssd1 vccd1 vccd1 _05832_ sky130_fd_sc_hd__xor2_1
XANTENNA__18008__A net519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13440__A _07575_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19154_ clknet_leaf_50_clk _00098_ net1367 vssd1 vssd1 vccd1 vccd1 ag2.body\[18\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_13_1072 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_920 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_16366_ obsg2.obstacleArray\[13\] net413 _02044_ net419 vssd1 vssd1 vccd1 vccd1 _02045_
+ sky130_fd_sc_hd__o211a_1
X_13578_ control.divider.fsm.current_mode\[2\] control.divider.fsm.current_mode\[0\]
+ vssd1 vssd1 vccd1 vccd1 _07953_ sky130_fd_sc_hd__nor2_2
X_18105_ net38 _03685_ vssd1 vssd1 vccd1 vccd1 _03686_ sky130_fd_sc_hd__and2_1
XFILLER_0_5_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15317_ net2308 net77 _01588_ control.body\[718\] vssd1 vssd1 vccd1 vccd1 _00616_
+ sky130_fd_sc_hd__a22o_1
X_12529_ net1786 net651 _07461_ vssd1 vssd1 vccd1 vccd1 img_gen.tracker.next_frame\[25\]
+ sky130_fd_sc_hd__and3_1
X_19085_ clknet_leaf_29_clk img_gen.tracker.next_frame\[523\] net1334 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[523\] sky130_fd_sc_hd__dfrtp_1
X_16297_ obsg2.obstacleArray\[112\] obsg2.obstacleArray\[113\] net406 vssd1 vssd1
+ vccd1 vccd1 _01976_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_1709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18036_ net39 _03640_ vssd1 vssd1 vccd1 vccd1 _03641_ sky130_fd_sc_hd__and2_1
X_15248_ control.body\[778\] net97 _01579_ net2161 vssd1 vssd1 vccd1 vccd1 _00556_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_111_113 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_1302 vccd1 vssd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11895__A net472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14271__A net1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15179_ control.body\[845\] net101 _01571_ net2331 vssd1 vssd1 vccd1 vccd1 _00495_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_103_1623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_1319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout308 net309 vssd1 vssd1 vccd1 vccd1 net308 sky130_fd_sc_hd__buf_4
Xfanout319 _01817_ vssd1 vssd1 vccd1 vccd1 net319 sky130_fd_sc_hd__clkbuf_4
X_19987_ clknet_leaf_65_clk _00931_ net1477 vssd1 vssd1 vccd1 vccd1 ag2.body\[401\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_96_1409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09740_ ag2.body\[359\] net1065 vssd1 vssd1 vccd1 vccd1 _04713_ sky130_fd_sc_hd__xor2_1
XANTENNA__10304__A net1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18938_ clknet_leaf_139_clk img_gen.tracker.next_frame\[376\] net1288 vssd1 vssd1
+ vccd1 vccd1 img_gen.tracker.frame\[376\] sky130_fd_sc_hd__dfrtp_1
.ends

