module tb_gameState;


endmodule