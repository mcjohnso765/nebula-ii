magic
tech sky130A
magscale 1 2
timestamp 1724863899
<< viali >>
rect 22753 37417 22787 37451
rect 23397 37417 23431 37451
rect 27077 37417 27111 37451
rect 28549 37417 28583 37451
rect 27353 37213 27387 37247
rect 23029 37145 23063 37179
rect 23673 37145 23707 37179
rect 28825 37145 28859 37179
rect 24961 36873 24995 36907
rect 25237 36873 25271 36907
rect 25697 36873 25731 36907
rect 27169 36873 27203 36907
rect 27629 36873 27663 36907
rect 28825 36873 28859 36907
rect 29469 36873 29503 36907
rect 30113 36873 30147 36907
rect 30849 36873 30883 36907
rect 31493 36873 31527 36907
rect 32321 36873 32355 36907
rect 32781 36873 32815 36907
rect 33425 36873 33459 36907
rect 34069 36873 34103 36907
rect 34713 36873 34747 36907
rect 35449 36873 35483 36907
rect 35909 36873 35943 36907
rect 36553 36873 36587 36907
rect 37473 36873 37507 36907
rect 37933 36873 37967 36907
rect 38577 36873 38611 36907
rect 39221 36873 39255 36907
rect 39865 36873 39899 36907
rect 40509 36873 40543 36907
rect 41153 36873 41187 36907
rect 41797 36873 41831 36907
rect 42625 36873 42659 36907
rect 43085 36873 43119 36907
rect 43729 36873 43763 36907
rect 44373 36873 44407 36907
rect 45017 36873 45051 36907
rect 45661 36873 45695 36907
rect 46397 36873 46431 36907
rect 46765 36873 46799 36907
rect 47133 36873 47167 36907
rect 24685 36737 24719 36771
rect 24777 36737 24811 36771
rect 25421 36737 25455 36771
rect 25881 36737 25915 36771
rect 25973 36737 26007 36771
rect 26801 36737 26835 36771
rect 26985 36737 27019 36771
rect 27813 36737 27847 36771
rect 27905 36737 27939 36771
rect 29009 36737 29043 36771
rect 29101 36737 29135 36771
rect 29653 36737 29687 36771
rect 29745 36737 29779 36771
rect 30297 36737 30331 36771
rect 30389 36737 30423 36771
rect 31033 36737 31067 36771
rect 31125 36737 31159 36771
rect 31677 36737 31711 36771
rect 31769 36737 31803 36771
rect 32137 36737 32171 36771
rect 32965 36737 32999 36771
rect 33057 36737 33091 36771
rect 33609 36737 33643 36771
rect 33701 36737 33735 36771
rect 34253 36737 34287 36771
rect 34345 36737 34379 36771
rect 34897 36737 34931 36771
rect 34989 36737 35023 36771
rect 35265 36737 35299 36771
rect 36093 36737 36127 36771
rect 36185 36737 36219 36771
rect 36737 36737 36771 36771
rect 36829 36737 36863 36771
rect 37289 36737 37323 36771
rect 38117 36737 38151 36771
rect 38209 36737 38243 36771
rect 38761 36737 38795 36771
rect 38853 36737 38887 36771
rect 39405 36737 39439 36771
rect 39497 36737 39531 36771
rect 40049 36737 40083 36771
rect 40141 36737 40175 36771
rect 40693 36737 40727 36771
rect 40785 36737 40819 36771
rect 41337 36737 41371 36771
rect 41429 36737 41463 36771
rect 41981 36737 42015 36771
rect 42073 36737 42107 36771
rect 42441 36737 42475 36771
rect 43269 36737 43303 36771
rect 43361 36737 43395 36771
rect 43913 36737 43947 36771
rect 44005 36737 44039 36771
rect 44557 36737 44591 36771
rect 44649 36737 44683 36771
rect 45201 36737 45235 36771
rect 45293 36737 45327 36771
rect 45845 36737 45879 36771
rect 45937 36737 45971 36771
rect 46213 36737 46247 36771
rect 46949 36737 46983 36771
rect 47317 36737 47351 36771
rect 47869 36737 47903 36771
rect 47593 36669 47627 36703
rect 24225 36329 24259 36363
rect 25329 36329 25363 36363
rect 32229 36329 32263 36363
rect 35265 36329 35299 36363
rect 37381 36329 37415 36363
rect 42533 36329 42567 36363
rect 46213 36329 46247 36363
rect 24961 36193 24995 36227
rect 22845 36125 22879 36159
rect 29377 36125 29411 36159
rect 23112 36057 23146 36091
rect 24409 36057 24443 36091
rect 28825 36057 28859 36091
rect 29101 36057 29135 36091
rect 29745 36057 29779 36091
rect 29929 36057 29963 36091
rect 30021 36057 30055 36091
rect 29561 35989 29595 36023
rect 30297 35989 30331 36023
rect 23213 35785 23247 35819
rect 23305 35785 23339 35819
rect 24133 35785 24167 35819
rect 29929 35785 29963 35819
rect 22089 35649 22123 35683
rect 23581 35649 23615 35683
rect 23673 35649 23707 35683
rect 23765 35649 23799 35683
rect 23949 35649 23983 35683
rect 28816 35649 28850 35683
rect 21833 35581 21867 35615
rect 25053 35581 25087 35615
rect 25329 35581 25363 35615
rect 28549 35581 28583 35615
rect 26801 35445 26835 35479
rect 21925 35241 21959 35275
rect 23581 35241 23615 35275
rect 25237 35241 25271 35275
rect 26065 35241 26099 35275
rect 28561 35241 28595 35275
rect 28917 35241 28951 35275
rect 29101 35241 29135 35275
rect 31677 35241 31711 35275
rect 22753 35105 22787 35139
rect 23305 35105 23339 35139
rect 28825 35105 28859 35139
rect 18613 35037 18647 35071
rect 22201 35037 22235 35071
rect 22293 35037 22327 35071
rect 22385 35037 22419 35071
rect 22569 35037 22603 35071
rect 24961 35037 24995 35071
rect 25145 35037 25179 35071
rect 25421 35037 25455 35071
rect 25697 35037 25731 35071
rect 25789 35037 25823 35071
rect 26065 35037 26099 35071
rect 26249 35037 26283 35071
rect 26985 35037 27019 35071
rect 31033 35037 31067 35071
rect 31861 35037 31895 35071
rect 21833 34969 21867 35003
rect 29285 34969 29319 35003
rect 17969 34901 18003 34935
rect 25053 34901 25087 34935
rect 25605 34901 25639 34935
rect 26341 34901 26375 34935
rect 27077 34901 27111 34935
rect 29085 34901 29119 34935
rect 31217 34901 31251 34935
rect 24869 34697 24903 34731
rect 26065 34629 26099 34663
rect 26709 34629 26743 34663
rect 26985 34629 27019 34663
rect 27185 34629 27219 34663
rect 16865 34561 16899 34595
rect 21281 34561 21315 34595
rect 22661 34561 22695 34595
rect 25513 34561 25547 34595
rect 26249 34561 26283 34595
rect 26433 34561 26467 34595
rect 26525 34561 26559 34595
rect 26801 34561 26835 34595
rect 30205 34561 30239 34595
rect 16957 34493 16991 34527
rect 17325 34493 17359 34527
rect 17601 34493 17635 34527
rect 19073 34493 19107 34527
rect 23121 34493 23155 34527
rect 23397 34493 23431 34527
rect 30481 34493 30515 34527
rect 32965 34493 32999 34527
rect 33241 34493 33275 34527
rect 34713 34493 34747 34527
rect 26525 34425 26559 34459
rect 17233 34357 17267 34391
rect 21189 34357 21223 34391
rect 24961 34357 24995 34391
rect 27169 34357 27203 34391
rect 27353 34357 27387 34391
rect 31953 34357 31987 34391
rect 21281 34153 21315 34187
rect 21741 34153 21775 34187
rect 30573 34153 30607 34187
rect 30757 34153 30791 34187
rect 31953 34153 31987 34187
rect 33057 34153 33091 34187
rect 33977 34153 34011 34187
rect 20269 34085 20303 34119
rect 26617 34085 26651 34119
rect 32873 34085 32907 34119
rect 34345 34085 34379 34119
rect 17693 34017 17727 34051
rect 20637 34017 20671 34051
rect 26157 34017 26191 34051
rect 34437 34017 34471 34051
rect 17785 33949 17819 33983
rect 17877 33949 17911 33983
rect 17969 33949 18003 33983
rect 20545 33949 20579 33983
rect 23949 33949 23983 33983
rect 24685 33949 24719 33983
rect 25789 33949 25823 33983
rect 26341 33949 26375 33983
rect 27353 33949 27387 33983
rect 31125 33949 31159 33983
rect 32137 33949 32171 33983
rect 32229 33949 32263 33983
rect 32505 33949 32539 33983
rect 32689 33949 32723 33983
rect 32781 33949 32815 33983
rect 33425 33949 33459 33983
rect 33885 33949 33919 33983
rect 34161 33949 34195 33983
rect 20269 33881 20303 33915
rect 20453 33881 20487 33915
rect 21925 33881 21959 33915
rect 25421 33881 25455 33915
rect 26617 33881 26651 33915
rect 26801 33881 26835 33915
rect 31953 33881 31987 33915
rect 32321 33881 32355 33915
rect 33241 33881 33275 33915
rect 33793 33881 33827 33915
rect 18153 33813 18187 33847
rect 21557 33813 21591 33847
rect 21725 33813 21759 33847
rect 25881 33813 25915 33847
rect 26433 33813 26467 33847
rect 30757 33813 30791 33847
rect 33031 33813 33065 33847
rect 33701 33813 33735 33847
rect 37105 33813 37139 33847
rect 21649 33609 21683 33643
rect 24409 33609 24443 33643
rect 27143 33609 27177 33643
rect 37105 33609 37139 33643
rect 20177 33541 20211 33575
rect 27353 33541 27387 33575
rect 36921 33541 36955 33575
rect 37565 33541 37599 33575
rect 16957 33473 16991 33507
rect 17141 33473 17175 33507
rect 22017 33473 22051 33507
rect 22201 33473 22235 33507
rect 23397 33473 23431 33507
rect 24684 33473 24718 33507
rect 24777 33473 24811 33507
rect 25053 33473 25087 33507
rect 29101 33473 29135 33507
rect 31125 33473 31159 33507
rect 32781 33473 32815 33507
rect 33241 33473 33275 33507
rect 33517 33473 33551 33507
rect 17233 33405 17267 33439
rect 17509 33405 17543 33439
rect 19901 33405 19935 33439
rect 22293 33405 22327 33439
rect 22477 33405 22511 33439
rect 23029 33405 23063 33439
rect 23213 33405 23247 33439
rect 25329 33405 25363 33439
rect 29377 33405 29411 33439
rect 30941 33405 30975 33439
rect 31401 33405 31435 33439
rect 33149 33405 33183 33439
rect 33793 33405 33827 33439
rect 37289 33405 37323 33439
rect 26801 33337 26835 33371
rect 31309 33337 31343 33371
rect 36553 33337 36587 33371
rect 17049 33269 17083 33303
rect 18981 33269 19015 33303
rect 21833 33269 21867 33303
rect 23581 33269 23615 33303
rect 26985 33269 27019 33303
rect 27169 33269 27203 33303
rect 30849 33269 30883 33303
rect 33057 33269 33091 33303
rect 33425 33269 33459 33303
rect 33793 33269 33827 33303
rect 34069 33269 34103 33303
rect 36921 33269 36955 33303
rect 39037 33269 39071 33303
rect 18245 33065 18279 33099
rect 19809 33065 19843 33099
rect 22569 33065 22603 33099
rect 24133 33065 24167 33099
rect 24961 33065 24995 33099
rect 25145 33065 25179 33099
rect 25789 33065 25823 33099
rect 26065 33065 26099 33099
rect 30389 33065 30423 33099
rect 33241 33065 33275 33099
rect 34069 33065 34103 33099
rect 38025 33065 38059 33099
rect 18337 32997 18371 33031
rect 23949 32997 23983 33031
rect 34253 32997 34287 33031
rect 16129 32929 16163 32963
rect 19533 32929 19567 32963
rect 21097 32929 21131 32963
rect 24409 32929 24443 32963
rect 27813 32929 27847 32963
rect 35817 32929 35851 32963
rect 14381 32861 14415 32895
rect 17049 32861 17083 32895
rect 17969 32861 18003 32895
rect 18153 32861 18187 32895
rect 19441 32861 19475 32895
rect 20821 32861 20855 32895
rect 23213 32861 23247 32895
rect 23397 32861 23431 32895
rect 23673 32861 23707 32895
rect 24777 32861 24811 32895
rect 25513 32861 25547 32895
rect 25789 32861 25823 32895
rect 25973 32861 26007 32895
rect 30573 32861 30607 32895
rect 30665 32861 30699 32895
rect 30757 32861 30791 32895
rect 30941 32861 30975 32895
rect 33425 32861 33459 32895
rect 33517 32861 33551 32895
rect 33701 32861 33735 32895
rect 33793 32861 33827 32895
rect 34345 32861 34379 32895
rect 34529 32861 34563 32895
rect 14657 32793 14691 32827
rect 17785 32793 17819 32827
rect 18705 32793 18739 32827
rect 19901 32793 19935 32827
rect 23305 32793 23339 32827
rect 27537 32793 27571 32827
rect 30389 32793 30423 32827
rect 33885 32793 33919 32827
rect 34101 32793 34135 32827
rect 36093 32793 36127 32827
rect 37657 32793 37691 32827
rect 37841 32793 37875 32827
rect 16405 32725 16439 32759
rect 17601 32725 17635 32759
rect 17877 32725 17911 32759
rect 19257 32725 19291 32759
rect 24593 32725 24627 32759
rect 30849 32725 30883 32759
rect 34437 32725 34471 32759
rect 37565 32725 37599 32759
rect 38209 32725 38243 32759
rect 15945 32521 15979 32555
rect 27353 32521 27387 32555
rect 34789 32521 34823 32555
rect 36093 32521 36127 32555
rect 36645 32521 36679 32555
rect 33149 32453 33183 32487
rect 33885 32453 33919 32487
rect 34069 32453 34103 32487
rect 34529 32453 34563 32487
rect 34989 32453 35023 32487
rect 33379 32419 33413 32453
rect 34299 32419 34333 32453
rect 16313 32385 16347 32419
rect 16773 32385 16807 32419
rect 26433 32385 26467 32419
rect 26985 32385 27019 32419
rect 27169 32385 27203 32419
rect 30113 32385 30147 32419
rect 30481 32385 30515 32419
rect 30665 32385 30699 32419
rect 35081 32385 35115 32419
rect 36277 32385 36311 32419
rect 36461 32385 36495 32419
rect 36553 32385 36587 32419
rect 36829 32385 36863 32419
rect 37013 32385 37047 32419
rect 16405 32317 16439 32351
rect 26525 32317 26559 32351
rect 26801 32317 26835 32351
rect 30389 32317 30423 32351
rect 30481 32249 30515 32283
rect 33517 32249 33551 32283
rect 34161 32249 34195 32283
rect 34621 32249 34655 32283
rect 17969 32181 18003 32215
rect 29929 32181 29963 32215
rect 30297 32181 30331 32215
rect 33333 32181 33367 32215
rect 33701 32181 33735 32215
rect 33885 32181 33919 32215
rect 34345 32181 34379 32215
rect 34805 32181 34839 32215
rect 19441 31977 19475 32011
rect 29824 31977 29858 32011
rect 31309 31977 31343 32011
rect 33793 31977 33827 32011
rect 34161 31977 34195 32011
rect 37473 31977 37507 32011
rect 15577 31909 15611 31943
rect 26065 31909 26099 31943
rect 37105 31909 37139 31943
rect 37657 31909 37691 31943
rect 17509 31841 17543 31875
rect 19349 31841 19383 31875
rect 20269 31841 20303 31875
rect 23857 31841 23891 31875
rect 24961 31841 24995 31875
rect 29561 31841 29595 31875
rect 15301 31773 15335 31807
rect 15577 31773 15611 31807
rect 15761 31773 15795 31807
rect 16405 31773 16439 31807
rect 18061 31773 18095 31807
rect 18153 31773 18187 31807
rect 18337 31773 18371 31807
rect 19257 31773 19291 31807
rect 19533 31773 19567 31807
rect 22098 31773 22132 31807
rect 25421 31773 25455 31807
rect 26157 31773 26191 31807
rect 26249 31773 26283 31807
rect 26341 31773 26375 31807
rect 29101 31773 29135 31807
rect 29285 31773 29319 31807
rect 29377 31773 29411 31807
rect 32321 31773 32355 31807
rect 33057 31773 33091 31807
rect 33149 31751 33183 31785
rect 33241 31773 33275 31807
rect 33609 31773 33643 31807
rect 33793 31773 33827 31807
rect 34161 31773 34195 31807
rect 34253 31773 34287 31807
rect 38117 31773 38151 31807
rect 15393 31705 15427 31739
rect 17233 31705 17267 31739
rect 20545 31705 20579 31739
rect 22385 31705 22419 31739
rect 33333 31705 33367 31739
rect 34437 31705 34471 31739
rect 37933 31705 37967 31739
rect 16313 31637 16347 31671
rect 18245 31637 18279 31671
rect 19717 31637 19751 31671
rect 22017 31637 22051 31671
rect 24409 31637 24443 31671
rect 29377 31637 29411 31671
rect 33517 31637 33551 31671
rect 33977 31637 34011 31671
rect 37473 31637 37507 31671
rect 37749 31637 37783 31671
rect 16681 31433 16715 31467
rect 18169 31433 18203 31467
rect 18337 31433 18371 31467
rect 21925 31433 21959 31467
rect 23857 31433 23891 31467
rect 24777 31433 24811 31467
rect 30481 31433 30515 31467
rect 36737 31433 36771 31467
rect 37289 31433 37323 31467
rect 17785 31365 17819 31399
rect 17969 31365 18003 31399
rect 22277 31365 22311 31399
rect 22477 31365 22511 31399
rect 23397 31365 23431 31399
rect 30665 31365 30699 31399
rect 31493 31365 31527 31399
rect 36889 31365 36923 31399
rect 37105 31365 37139 31399
rect 38761 31365 38795 31399
rect 13921 31297 13955 31331
rect 16129 31297 16163 31331
rect 18521 31297 18555 31331
rect 18717 31297 18751 31331
rect 18981 31297 19015 31331
rect 20177 31297 20211 31331
rect 20913 31297 20947 31331
rect 21465 31297 21499 31331
rect 21833 31297 21867 31331
rect 22017 31297 22051 31331
rect 22661 31297 22695 31331
rect 23673 31297 23707 31331
rect 24685 31297 24719 31331
rect 24961 31297 24995 31331
rect 25053 31297 25087 31331
rect 25697 31297 25731 31331
rect 26525 31297 26559 31331
rect 26709 31297 26743 31331
rect 28457 31297 28491 31331
rect 33425 31297 33459 31331
rect 33517 31297 33551 31331
rect 33885 31297 33919 31331
rect 34345 31297 34379 31331
rect 34713 31297 34747 31331
rect 14197 31229 14231 31263
rect 15761 31229 15795 31263
rect 16221 31229 16255 31263
rect 17233 31229 17267 31263
rect 18797 31229 18831 31263
rect 19809 31229 19843 31263
rect 20269 31229 20303 31263
rect 20545 31229 20579 31263
rect 23581 31229 23615 31263
rect 26341 31229 26375 31263
rect 28733 31229 28767 31263
rect 34253 31229 34287 31263
rect 36645 31229 36679 31263
rect 39037 31229 39071 31263
rect 15669 31161 15703 31195
rect 19165 31161 19199 31195
rect 24961 31161 24995 31195
rect 26617 31161 26651 31195
rect 17509 31093 17543 31127
rect 18153 31093 18187 31127
rect 18521 31093 18555 31127
rect 19257 31093 19291 31127
rect 22109 31093 22143 31127
rect 22293 31093 22327 31127
rect 23213 31093 23247 31127
rect 23673 31093 23707 31127
rect 25789 31093 25823 31127
rect 30205 31093 30239 31127
rect 33793 31093 33827 31127
rect 34069 31093 34103 31127
rect 34621 31093 34655 31127
rect 34897 31093 34931 31127
rect 36921 31093 36955 31127
rect 15577 30889 15611 30923
rect 17877 30889 17911 30923
rect 23121 30889 23155 30923
rect 25053 30889 25087 30923
rect 25973 30889 26007 30923
rect 30297 30889 30331 30923
rect 33609 30889 33643 30923
rect 34272 30889 34306 30923
rect 34897 30889 34931 30923
rect 36369 30889 36403 30923
rect 36829 30889 36863 30923
rect 19257 30821 19291 30855
rect 25237 30821 25271 30855
rect 34161 30821 34195 30855
rect 25605 30753 25639 30787
rect 25881 30753 25915 30787
rect 27445 30753 27479 30787
rect 27721 30753 27755 30787
rect 31033 30753 31067 30787
rect 33517 30753 33551 30787
rect 34071 30753 34105 30787
rect 17325 30685 17359 30719
rect 17785 30685 17819 30719
rect 17969 30685 18003 30719
rect 19257 30685 19291 30719
rect 19441 30685 19475 30719
rect 22845 30685 22879 30719
rect 22937 30685 22971 30719
rect 23121 30685 23155 30719
rect 25513 30685 25547 30719
rect 30481 30685 30515 30719
rect 30573 30685 30607 30719
rect 33333 30685 33367 30719
rect 33609 30685 33643 30719
rect 34437 30685 34471 30719
rect 34897 30685 34931 30719
rect 35081 30685 35115 30719
rect 36553 30685 36587 30719
rect 36645 30685 36679 30719
rect 36921 30685 36955 30719
rect 17049 30617 17083 30651
rect 24869 30617 24903 30651
rect 31309 30617 31343 30651
rect 35357 30617 35391 30651
rect 37197 30617 37231 30651
rect 38761 30617 38795 30651
rect 18153 30549 18187 30583
rect 25069 30549 25103 30583
rect 32781 30549 32815 30583
rect 33149 30549 33183 30583
rect 33793 30549 33827 30583
rect 34713 30549 34747 30583
rect 38669 30549 38703 30583
rect 19809 30345 19843 30379
rect 24317 30345 24351 30379
rect 25053 30345 25087 30379
rect 32965 30345 32999 30379
rect 33517 30345 33551 30379
rect 18337 30277 18371 30311
rect 19993 30277 20027 30311
rect 22477 30277 22511 30311
rect 26525 30277 26559 30311
rect 32689 30277 32723 30311
rect 33333 30277 33367 30311
rect 33793 30277 33827 30311
rect 33993 30277 34027 30311
rect 38669 30277 38703 30311
rect 38853 30277 38887 30311
rect 42257 30277 42291 30311
rect 18061 30209 18095 30243
rect 22569 30209 22603 30243
rect 32965 30209 32999 30243
rect 33609 30209 33643 30243
rect 38577 30209 38611 30243
rect 42441 30209 42475 30243
rect 42533 30209 42567 30243
rect 42717 30209 42751 30243
rect 22845 30141 22879 30175
rect 26801 30141 26835 30175
rect 37841 30141 37875 30175
rect 42809 30141 42843 30175
rect 43085 30141 43119 30175
rect 44833 30141 44867 30175
rect 32873 30073 32907 30107
rect 33333 30073 33367 30107
rect 34161 30073 34195 30107
rect 39129 30073 39163 30107
rect 42717 30073 42751 30107
rect 33977 30005 34011 30039
rect 34621 30005 34655 30039
rect 39037 30005 39071 30039
rect 22569 29801 22603 29835
rect 28825 29801 28859 29835
rect 34253 29801 34287 29835
rect 35081 29801 35115 29835
rect 37289 29801 37323 29835
rect 37473 29801 37507 29835
rect 43453 29801 43487 29835
rect 29745 29733 29779 29767
rect 37841 29733 37875 29767
rect 38025 29733 38059 29767
rect 40877 29733 40911 29767
rect 22845 29665 22879 29699
rect 24961 29665 24995 29699
rect 38209 29665 38243 29699
rect 40509 29665 40543 29699
rect 44557 29665 44591 29699
rect 22937 29597 22971 29631
rect 24409 29597 24443 29631
rect 29101 29597 29135 29631
rect 29285 29597 29319 29631
rect 29561 29597 29595 29631
rect 33793 29597 33827 29631
rect 33977 29597 34011 29631
rect 34897 29597 34931 29631
rect 37933 29597 37967 29631
rect 40233 29597 40267 29631
rect 40325 29597 40359 29631
rect 40601 29597 40635 29631
rect 43269 29597 43303 29631
rect 43453 29597 43487 29631
rect 43637 29597 43671 29631
rect 47409 29597 47443 29631
rect 29009 29529 29043 29563
rect 29653 29529 29687 29563
rect 29837 29529 29871 29563
rect 32413 29529 32447 29563
rect 32597 29529 32631 29563
rect 34069 29529 34103 29563
rect 34713 29529 34747 29563
rect 37473 29529 37507 29563
rect 40877 29529 40911 29563
rect 44005 29529 44039 29563
rect 45385 29529 45419 29563
rect 47133 29529 47167 29563
rect 28641 29461 28675 29495
rect 28809 29461 28843 29495
rect 29101 29461 29135 29495
rect 32781 29461 32815 29495
rect 33977 29461 34011 29495
rect 34269 29461 34303 29495
rect 34437 29461 34471 29495
rect 38209 29461 38243 29495
rect 40509 29461 40543 29495
rect 40693 29461 40727 29495
rect 42717 29461 42751 29495
rect 47501 29461 47535 29495
rect 30481 29257 30515 29291
rect 33977 29257 34011 29291
rect 37105 29257 37139 29291
rect 40417 29257 40451 29291
rect 43821 29257 43855 29291
rect 46029 29257 46063 29291
rect 46489 29257 46523 29291
rect 27353 29189 27387 29223
rect 27537 29189 27571 29223
rect 28273 29189 28307 29223
rect 28489 29189 28523 29223
rect 37657 29189 37691 29223
rect 42993 29189 43027 29223
rect 27905 29121 27939 29155
rect 31769 29121 31803 29155
rect 31953 29121 31987 29155
rect 32137 29121 32171 29155
rect 35725 29121 35759 29155
rect 37381 29121 37415 29155
rect 39405 29121 39439 29155
rect 39773 29121 39807 29155
rect 40049 29121 40083 29155
rect 40203 29121 40237 29155
rect 40601 29121 40635 29155
rect 40785 29121 40819 29155
rect 40877 29121 40911 29155
rect 41153 29121 41187 29155
rect 41429 29121 41463 29155
rect 41521 29121 41555 29155
rect 43453 29121 43487 29155
rect 44005 29121 44039 29155
rect 44097 29121 44131 29155
rect 44189 29121 44223 29155
rect 46121 29121 46155 29155
rect 26525 29053 26559 29087
rect 28733 29053 28767 29087
rect 29009 29053 29043 29087
rect 32413 29053 32447 29087
rect 35449 29053 35483 29087
rect 41245 29053 41279 29087
rect 41613 29053 41647 29087
rect 41705 29053 41739 29087
rect 43545 29053 43579 29087
rect 45661 29053 45695 29087
rect 45937 29053 45971 29087
rect 26249 28985 26283 29019
rect 27169 28985 27203 29019
rect 28089 28985 28123 29019
rect 28641 28985 28675 29019
rect 41061 28985 41095 29019
rect 42993 28985 43027 29019
rect 26065 28917 26099 28951
rect 28457 28917 28491 28951
rect 31861 28917 31895 28951
rect 33885 28917 33919 28951
rect 39681 28917 39715 28951
rect 43729 28917 43763 28951
rect 27353 28713 27387 28747
rect 28825 28713 28859 28747
rect 30665 28713 30699 28747
rect 32321 28713 32355 28747
rect 32505 28713 32539 28747
rect 32689 28713 32723 28747
rect 38025 28713 38059 28747
rect 38577 28713 38611 28747
rect 42993 28713 43027 28747
rect 43729 28713 43763 28747
rect 44189 28713 44223 28747
rect 45753 28713 45787 28747
rect 40601 28645 40635 28679
rect 44465 28645 44499 28679
rect 25605 28577 25639 28611
rect 36001 28577 36035 28611
rect 42717 28577 42751 28611
rect 29193 28509 29227 28543
rect 30021 28509 30055 28543
rect 30205 28509 30239 28543
rect 30481 28509 30515 28543
rect 32689 28509 32723 28543
rect 32873 28509 32907 28543
rect 33057 28509 33091 28543
rect 33149 28509 33183 28543
rect 38761 28509 38795 28543
rect 40233 28509 40267 28543
rect 40387 28509 40421 28543
rect 42809 28509 42843 28543
rect 43177 28509 43211 28543
rect 43269 28509 43303 28543
rect 43453 28509 43487 28543
rect 43545 28509 43579 28543
rect 43637 28519 43671 28553
rect 43913 28509 43947 28543
rect 45017 28509 45051 28543
rect 45201 28509 45235 28543
rect 45293 28509 45327 28543
rect 45661 28509 45695 28543
rect 50905 28509 50939 28543
rect 25881 28441 25915 28475
rect 29009 28441 29043 28475
rect 32137 28441 32171 28475
rect 32337 28441 32371 28475
rect 36277 28441 36311 28475
rect 38485 28441 38519 28475
rect 38945 28441 38979 28475
rect 44741 28441 44775 28475
rect 30297 28373 30331 28407
rect 37749 28373 37783 28407
rect 44281 28373 44315 28407
rect 50353 28373 50387 28407
rect 30021 28169 30055 28203
rect 37289 28169 37323 28203
rect 46857 28169 46891 28203
rect 47777 28169 47811 28203
rect 28549 28101 28583 28135
rect 37013 28101 37047 28135
rect 40141 28101 40175 28135
rect 45201 28101 45235 28135
rect 46949 28101 46983 28135
rect 50997 28101 51031 28135
rect 37657 28033 37691 28067
rect 42257 28033 42291 28067
rect 42717 28033 42751 28067
rect 42809 28033 42843 28067
rect 42993 28033 43027 28067
rect 43085 28033 43119 28067
rect 43729 28033 43763 28067
rect 44097 28033 44131 28067
rect 44557 28033 44591 28067
rect 45017 28033 45051 28067
rect 47593 28033 47627 28067
rect 49617 28033 49651 28067
rect 49893 28033 49927 28067
rect 50261 28033 50295 28067
rect 28273 27965 28307 27999
rect 37749 27965 37783 27999
rect 37841 27965 37875 27999
rect 42165 27965 42199 27999
rect 43269 27965 43303 27999
rect 44373 27965 44407 27999
rect 44649 27965 44683 27999
rect 44741 27965 44775 27999
rect 44833 27965 44867 27999
rect 47133 27965 47167 27999
rect 40509 27897 40543 27931
rect 44097 27897 44131 27931
rect 46397 27897 46431 27931
rect 40601 27829 40635 27863
rect 42533 27829 42567 27863
rect 45385 27829 45419 27863
rect 46489 27829 46523 27863
rect 49433 27829 49467 27863
rect 49801 27829 49835 27863
rect 50077 27829 50111 27863
rect 37920 27625 37954 27659
rect 43085 27625 43119 27659
rect 43269 27625 43303 27659
rect 43637 27625 43671 27659
rect 44005 27625 44039 27659
rect 44649 27625 44683 27659
rect 46654 27625 46688 27659
rect 48145 27625 48179 27659
rect 39865 27557 39899 27591
rect 40969 27557 41003 27591
rect 48329 27557 48363 27591
rect 32505 27489 32539 27523
rect 34713 27489 34747 27523
rect 40509 27489 40543 27523
rect 44189 27489 44223 27523
rect 51917 27489 51951 27523
rect 52561 27489 52595 27523
rect 30389 27421 30423 27455
rect 30573 27421 30607 27455
rect 30941 27421 30975 27455
rect 32873 27421 32907 27455
rect 35081 27421 35115 27455
rect 37657 27421 37691 27455
rect 41245 27421 41279 27455
rect 41521 27421 41555 27455
rect 42533 27421 42567 27455
rect 42625 27421 42659 27455
rect 42901 27421 42935 27455
rect 43085 27421 43119 27455
rect 43177 27421 43211 27455
rect 43361 27421 43395 27455
rect 44281 27421 44315 27455
rect 44557 27421 44591 27455
rect 46397 27421 46431 27455
rect 49709 27421 49743 27455
rect 50169 27421 50203 27455
rect 29377 27353 29411 27387
rect 29561 27353 29595 27387
rect 39681 27353 39715 27387
rect 41061 27353 41095 27387
rect 41797 27353 41831 27387
rect 43453 27353 43487 27387
rect 43669 27353 43703 27387
rect 50445 27353 50479 27387
rect 32367 27285 32401 27319
rect 34299 27285 34333 27319
rect 36507 27285 36541 27319
rect 40233 27285 40267 27319
rect 40325 27285 40359 27319
rect 43821 27285 43855 27319
rect 52009 27285 52043 27319
rect 32137 27081 32171 27115
rect 32781 27081 32815 27115
rect 33425 27081 33459 27115
rect 39957 27081 39991 27115
rect 43453 27081 43487 27115
rect 43821 27081 43855 27115
rect 50721 27081 50755 27115
rect 52469 27081 52503 27115
rect 47593 27013 47627 27047
rect 49157 27013 49191 27047
rect 32321 26945 32355 26979
rect 32413 26945 32447 26979
rect 32689 26945 32723 26979
rect 32965 26945 32999 26979
rect 33057 26945 33091 26979
rect 33333 26945 33367 26979
rect 33609 26945 33643 26979
rect 33701 26945 33735 26979
rect 33793 26945 33827 26979
rect 33957 26945 33991 26979
rect 34529 26945 34563 26979
rect 34713 26945 34747 26979
rect 34805 26945 34839 26979
rect 34897 26945 34931 26979
rect 37013 26945 37047 26979
rect 40141 26945 40175 26979
rect 40969 26945 41003 26979
rect 41153 26945 41187 26979
rect 41245 26945 41279 26979
rect 41521 26945 41555 26979
rect 43269 26945 43303 26979
rect 43545 26945 43579 26979
rect 43637 26945 43671 26979
rect 43913 26945 43947 26979
rect 47041 26945 47075 26979
rect 47133 26945 47167 26979
rect 47409 26945 47443 26979
rect 48145 26945 48179 26979
rect 50905 26945 50939 26979
rect 51181 26945 51215 26979
rect 23213 26877 23247 26911
rect 23489 26877 23523 26911
rect 25053 26877 25087 26911
rect 25329 26877 25363 26911
rect 27353 26877 27387 26911
rect 27629 26877 27663 26911
rect 36645 26877 36679 26911
rect 40325 26877 40359 26911
rect 41429 26877 41463 26911
rect 48697 26877 48731 26911
rect 48881 26877 48915 26911
rect 50629 26877 50663 26911
rect 52745 26877 52779 26911
rect 53021 26877 53055 26911
rect 47317 26809 47351 26843
rect 24961 26741 24995 26775
rect 26801 26741 26835 26775
rect 29101 26741 29135 26775
rect 32597 26741 32631 26775
rect 33241 26741 33275 26775
rect 35081 26741 35115 26775
rect 35219 26741 35253 26775
rect 39773 26741 39807 26775
rect 43085 26741 43119 26775
rect 43637 26741 43671 26775
rect 46857 26741 46891 26775
rect 51089 26741 51123 26775
rect 54493 26741 54527 26775
rect 24409 26537 24443 26571
rect 25145 26537 25179 26571
rect 32321 26537 32355 26571
rect 34897 26537 34931 26571
rect 38945 26537 38979 26571
rect 40233 26537 40267 26571
rect 48329 26537 48363 26571
rect 49341 26537 49375 26571
rect 50813 26537 50847 26571
rect 52469 26537 52503 26571
rect 25789 26469 25823 26503
rect 27537 26469 27571 26503
rect 29009 26469 29043 26503
rect 36093 26469 36127 26503
rect 39129 26469 39163 26503
rect 45937 26469 45971 26503
rect 46397 26469 46431 26503
rect 58449 26469 58483 26503
rect 25605 26401 25639 26435
rect 26433 26401 26467 26435
rect 30205 26401 30239 26435
rect 35357 26401 35391 26435
rect 36185 26401 36219 26435
rect 36645 26401 36679 26435
rect 39681 26401 39715 26435
rect 40601 26401 40635 26435
rect 41245 26401 41279 26435
rect 46581 26401 46615 26435
rect 46857 26401 46891 26435
rect 52837 26401 52871 26435
rect 24593 26333 24627 26367
rect 24777 26333 24811 26367
rect 24869 26333 24903 26367
rect 25329 26333 25363 26367
rect 25421 26333 25455 26367
rect 25697 26333 25731 26367
rect 25973 26333 26007 26367
rect 26341 26333 26375 26367
rect 26985 26333 27019 26367
rect 27721 26333 27755 26367
rect 28089 26333 28123 26367
rect 28733 26333 28767 26367
rect 28825 26333 28859 26367
rect 29101 26333 29135 26367
rect 29653 26333 29687 26367
rect 32505 26333 32539 26367
rect 32597 26333 32631 26367
rect 32873 26333 32907 26367
rect 35081 26333 35115 26367
rect 35173 26333 35207 26367
rect 35449 26333 35483 26367
rect 35541 26333 35575 26367
rect 35725 26333 35759 26367
rect 35909 26333 35943 26367
rect 36369 26333 36403 26367
rect 36461 26333 36495 26367
rect 36737 26333 36771 26367
rect 38853 26333 38887 26367
rect 39037 26333 39071 26367
rect 39497 26333 39531 26367
rect 40693 26333 40727 26367
rect 40969 26333 41003 26367
rect 46213 26333 46247 26367
rect 46489 26333 46523 26367
rect 49520 26333 49554 26367
rect 49892 26333 49926 26367
rect 49985 26333 50019 26367
rect 50169 26333 50203 26367
rect 50262 26333 50296 26367
rect 50537 26333 50571 26367
rect 50634 26333 50668 26367
rect 52653 26333 52687 26367
rect 52929 26333 52963 26367
rect 53573 26333 53607 26367
rect 54125 26333 54159 26367
rect 58265 26333 58299 26367
rect 40187 26299 40221 26333
rect 26065 26265 26099 26299
rect 26157 26265 26191 26299
rect 27813 26265 27847 26299
rect 27905 26265 27939 26299
rect 32689 26265 32723 26299
rect 35817 26265 35851 26299
rect 40417 26265 40451 26299
rect 49617 26265 49651 26299
rect 49709 26265 49743 26299
rect 50445 26265 50479 26299
rect 22753 26197 22787 26231
rect 28549 26197 28583 26231
rect 39313 26197 39347 26231
rect 39405 26197 39439 26231
rect 40049 26197 40083 26231
rect 46029 26197 46063 26231
rect 24685 25993 24719 26027
rect 30113 25993 30147 26027
rect 39247 25993 39281 26027
rect 42625 25993 42659 26027
rect 42917 25993 42951 26027
rect 44557 25993 44591 26027
rect 47593 25993 47627 26027
rect 48329 25993 48363 26027
rect 52193 25993 52227 26027
rect 25145 25925 25179 25959
rect 28641 25925 28675 25959
rect 32413 25925 32447 25959
rect 35909 25925 35943 25959
rect 39037 25925 39071 25959
rect 42717 25925 42751 25959
rect 43821 25925 43855 25959
rect 45845 25925 45879 25959
rect 51825 25925 51859 25959
rect 51917 25925 51951 25959
rect 53021 25925 53055 25959
rect 53113 25925 53147 25959
rect 19073 25857 19107 25891
rect 19165 25857 19199 25891
rect 19441 25857 19475 25891
rect 22104 25857 22138 25891
rect 22201 25857 22235 25891
rect 22293 25857 22327 25891
rect 22476 25857 22510 25891
rect 22569 25857 22603 25891
rect 22845 25857 22879 25891
rect 25007 25857 25041 25891
rect 25237 25857 25271 25891
rect 25420 25857 25454 25891
rect 25513 25857 25547 25891
rect 27721 25857 27755 25891
rect 27905 25857 27939 25891
rect 27997 25857 28031 25891
rect 28273 25857 28307 25891
rect 28365 25857 28399 25891
rect 32137 25857 32171 25891
rect 32321 25857 32355 25891
rect 32505 25857 32539 25891
rect 35725 25857 35759 25891
rect 35817 25857 35851 25891
rect 36093 25857 36127 25891
rect 39681 25857 39715 25891
rect 43913 25857 43947 25891
rect 44005 25857 44039 25891
rect 44189 25857 44223 25891
rect 48513 25857 48547 25891
rect 48605 25857 48639 25891
rect 48697 25857 48731 25891
rect 48881 25857 48915 25891
rect 49985 25857 50019 25891
rect 50261 25857 50295 25891
rect 51549 25857 51583 25891
rect 51642 25857 51676 25891
rect 52055 25857 52089 25891
rect 52883 25857 52917 25891
rect 53241 25857 53275 25891
rect 53389 25857 53423 25891
rect 56701 25857 56735 25891
rect 56885 25857 56919 25891
rect 57069 25857 57103 25891
rect 57161 25857 57195 25891
rect 57253 25857 57287 25891
rect 57897 25857 57931 25891
rect 23121 25789 23155 25823
rect 23213 25789 23247 25823
rect 23765 25789 23799 25823
rect 39497 25789 39531 25823
rect 39957 25789 39991 25823
rect 40049 25789 40083 25823
rect 43177 25789 43211 25823
rect 43361 25789 43395 25823
rect 43453 25789 43487 25823
rect 45569 25789 45603 25823
rect 47317 25789 47351 25823
rect 48145 25789 48179 25823
rect 50169 25789 50203 25823
rect 54493 25789 54527 25823
rect 55965 25789 55999 25823
rect 56241 25789 56275 25823
rect 58449 25789 58483 25823
rect 19349 25721 19383 25755
rect 24869 25721 24903 25755
rect 25881 25721 25915 25755
rect 43085 25721 43119 25755
rect 50445 25721 50479 25755
rect 18889 25653 18923 25687
rect 21925 25653 21959 25687
rect 22661 25653 22695 25687
rect 23029 25653 23063 25687
rect 28181 25653 28215 25687
rect 32689 25653 32723 25687
rect 35541 25653 35575 25687
rect 39221 25653 39255 25687
rect 39405 25653 39439 25687
rect 40233 25653 40267 25687
rect 42901 25653 42935 25687
rect 44373 25653 44407 25687
rect 49985 25653 50019 25687
rect 51365 25653 51399 25687
rect 52745 25653 52779 25687
rect 56517 25653 56551 25687
rect 57529 25653 57563 25687
rect 17588 25449 17622 25483
rect 19993 25449 20027 25483
rect 20453 25449 20487 25483
rect 21005 25449 21039 25483
rect 23305 25449 23339 25483
rect 28917 25449 28951 25483
rect 36507 25449 36541 25483
rect 41613 25449 41647 25483
rect 42993 25449 43027 25483
rect 43361 25449 43395 25483
rect 43821 25449 43855 25483
rect 48237 25449 48271 25483
rect 50169 25449 50203 25483
rect 56057 25449 56091 25483
rect 58265 25449 58299 25483
rect 26617 25381 26651 25415
rect 33517 25381 33551 25415
rect 37197 25381 37231 25415
rect 39405 25381 39439 25415
rect 41797 25381 41831 25415
rect 42533 25381 42567 25415
rect 44281 25381 44315 25415
rect 49617 25381 49651 25415
rect 54677 25381 54711 25415
rect 17325 25313 17359 25347
rect 19073 25313 19107 25347
rect 21465 25313 21499 25347
rect 23213 25313 23247 25347
rect 26433 25313 26467 25347
rect 31125 25313 31159 25347
rect 31493 25313 31527 25347
rect 33057 25313 33091 25347
rect 34713 25313 34747 25347
rect 37749 25313 37783 25347
rect 38209 25313 38243 25347
rect 40509 25313 40543 25347
rect 41981 25313 42015 25347
rect 42073 25313 42107 25347
rect 42165 25313 42199 25347
rect 44373 25313 44407 25347
rect 47501 25313 47535 25347
rect 52101 25313 52135 25347
rect 52193 25313 52227 25347
rect 56885 25313 56919 25347
rect 19533 25245 19567 25279
rect 19901 25245 19935 25279
rect 20177 25245 20211 25279
rect 20269 25245 20303 25279
rect 20545 25245 20579 25279
rect 20913 25245 20947 25279
rect 21189 25245 21223 25279
rect 23484 25245 23518 25279
rect 23856 25245 23890 25279
rect 23949 25245 23983 25279
rect 25784 25245 25818 25279
rect 25881 25245 25915 25279
rect 26156 25245 26190 25279
rect 26249 25245 26283 25279
rect 28365 25245 28399 25279
rect 28733 25245 28767 25279
rect 29285 25245 29319 25279
rect 29561 25245 29595 25279
rect 33241 25245 33275 25279
rect 33333 25245 33367 25279
rect 33609 25245 33643 25279
rect 35081 25245 35115 25279
rect 36645 25245 36679 25279
rect 36921 25245 36955 25279
rect 37013 25245 37047 25279
rect 37841 25245 37875 25279
rect 38117 25245 38151 25279
rect 38664 25245 38698 25279
rect 38761 25245 38795 25279
rect 39036 25245 39070 25279
rect 39129 25245 39163 25279
rect 40024 25245 40058 25279
rect 40141 25245 40175 25279
rect 41337 25255 41371 25289
rect 42257 25245 42291 25279
rect 42809 25245 42843 25279
rect 43545 25245 43579 25279
rect 43637 25245 43671 25279
rect 45661 25245 45695 25279
rect 48053 25245 48087 25279
rect 48375 25245 48409 25279
rect 48788 25245 48822 25279
rect 48881 25245 48915 25279
rect 49065 25245 49099 25279
rect 49341 25245 49375 25279
rect 49433 25245 49467 25279
rect 49709 25245 49743 25279
rect 50307 25245 50341 25279
rect 50445 25245 50479 25279
rect 50720 25245 50754 25279
rect 50813 25245 50847 25279
rect 51825 25245 51859 25279
rect 52009 25245 52043 25279
rect 54033 25245 54067 25279
rect 54126 25245 54160 25279
rect 54498 25245 54532 25279
rect 55321 25245 55355 25279
rect 56241 25245 56275 25279
rect 56425 25245 56459 25279
rect 56517 25245 56551 25279
rect 57152 25245 57186 25279
rect 19625 25177 19659 25211
rect 19717 25177 19751 25211
rect 21741 25177 21775 25211
rect 23581 25177 23615 25211
rect 23673 25177 23707 25211
rect 25973 25177 26007 25211
rect 28549 25177 28583 25211
rect 28641 25177 28675 25211
rect 32919 25177 32953 25211
rect 36829 25177 36863 25211
rect 37473 25177 37507 25211
rect 38853 25177 38887 25211
rect 40233 25177 40267 25211
rect 41429 25177 41463 25211
rect 41645 25177 41679 25211
rect 42717 25177 42751 25211
rect 45937 25177 45971 25211
rect 48513 25177 48547 25211
rect 48605 25177 48639 25211
rect 49249 25177 49283 25211
rect 50537 25177 50571 25211
rect 51641 25177 51675 25211
rect 52469 25177 52503 25211
rect 54309 25177 54343 25211
rect 54401 25177 54435 25211
rect 55965 25177 55999 25211
rect 19349 25109 19383 25143
rect 21373 25109 21407 25143
rect 24133 25109 24167 25143
rect 25605 25109 25639 25143
rect 26801 25109 26835 25143
rect 29101 25109 29135 25143
rect 37289 25109 37323 25143
rect 38393 25109 38427 25143
rect 38485 25109 38519 25143
rect 39221 25109 39255 25143
rect 39865 25109 39899 25143
rect 41245 25109 41279 25143
rect 42441 25109 42475 25143
rect 47409 25109 47443 25143
rect 49893 25109 49927 25143
rect 50905 25109 50939 25143
rect 53941 25109 53975 25143
rect 19809 24905 19843 24939
rect 26525 24905 26559 24939
rect 32137 24905 32171 24939
rect 45845 24905 45879 24939
rect 45937 24905 45971 24939
rect 50077 24905 50111 24939
rect 50445 24905 50479 24939
rect 18245 24837 18279 24871
rect 20177 24837 20211 24871
rect 22109 24837 22143 24871
rect 25145 24837 25179 24871
rect 32413 24837 32447 24871
rect 36001 24837 36035 24871
rect 38009 24837 38043 24871
rect 38209 24837 38243 24871
rect 39773 24837 39807 24871
rect 43269 24837 43303 24871
rect 48789 24837 48823 24871
rect 49801 24837 49835 24871
rect 50721 24837 50755 24871
rect 55597 24837 55631 24871
rect 17969 24769 18003 24803
rect 19993 24769 20027 24803
rect 20085 24769 20119 24803
rect 20361 24769 20395 24803
rect 24961 24769 24995 24803
rect 25237 24769 25271 24803
rect 25329 24769 25363 24803
rect 25789 24769 25823 24803
rect 25881 24769 25915 24803
rect 26065 24769 26099 24803
rect 26157 24769 26191 24803
rect 31585 24769 31619 24803
rect 31677 24769 31711 24803
rect 31953 24769 31987 24803
rect 32321 24769 32355 24803
rect 32505 24769 32539 24803
rect 32689 24769 32723 24803
rect 34989 24769 35023 24803
rect 35357 24769 35391 24803
rect 35541 24769 35575 24803
rect 35633 24769 35667 24803
rect 35909 24769 35943 24803
rect 37473 24769 37507 24803
rect 37749 24769 37783 24803
rect 39865 24769 39899 24803
rect 40877 24769 40911 24803
rect 40969 24769 41003 24803
rect 41061 24769 41095 24803
rect 41245 24769 41279 24803
rect 41613 24769 41647 24803
rect 41797 24769 41831 24803
rect 41889 24769 41923 24803
rect 41981 24769 42015 24803
rect 42625 24769 42659 24803
rect 42717 24769 42751 24803
rect 46121 24769 46155 24803
rect 46305 24769 46339 24803
rect 46397 24769 46431 24803
rect 46581 24769 46615 24803
rect 49617 24769 49651 24803
rect 49709 24769 49743 24803
rect 49985 24769 50019 24803
rect 50261 24769 50295 24803
rect 50537 24769 50571 24803
rect 52837 24769 52871 24803
rect 55229 24769 55263 24803
rect 55377 24769 55411 24803
rect 55505 24769 55539 24803
rect 55694 24769 55728 24803
rect 21833 24701 21867 24735
rect 27537 24701 27571 24735
rect 27813 24701 27847 24735
rect 29285 24701 29319 24735
rect 29929 24701 29963 24735
rect 35817 24701 35851 24735
rect 37657 24701 37691 24735
rect 43821 24701 43855 24735
rect 49249 24701 49283 24735
rect 53389 24701 53423 24735
rect 55965 24701 55999 24735
rect 56241 24701 56275 24735
rect 19717 24633 19751 24667
rect 25605 24633 25639 24667
rect 37841 24633 37875 24667
rect 40601 24633 40635 24667
rect 42257 24633 42291 24667
rect 43545 24633 43579 24667
rect 47593 24633 47627 24667
rect 20453 24565 20487 24599
rect 21557 24565 21591 24599
rect 23581 24565 23615 24599
rect 24869 24565 24903 24599
rect 25513 24565 25547 24599
rect 26341 24565 26375 24599
rect 29377 24565 29411 24599
rect 31401 24565 31435 24599
rect 31861 24565 31895 24599
rect 37289 24565 37323 24599
rect 37473 24565 37507 24599
rect 38025 24565 38059 24599
rect 39589 24565 39623 24599
rect 40049 24565 40083 24599
rect 40509 24565 40543 24599
rect 42441 24565 42475 24599
rect 42901 24565 42935 24599
rect 43729 24565 43763 24599
rect 46857 24565 46891 24599
rect 47133 24565 47167 24599
rect 47317 24565 47351 24599
rect 49065 24565 49099 24599
rect 49433 24565 49467 24599
rect 55873 24565 55907 24599
rect 57713 24565 57747 24599
rect 22845 24361 22879 24395
rect 24961 24361 24995 24395
rect 25421 24361 25455 24395
rect 26157 24361 26191 24395
rect 26525 24361 26559 24395
rect 27997 24361 28031 24395
rect 28457 24361 28491 24395
rect 32827 24361 32861 24395
rect 34069 24361 34103 24395
rect 34529 24361 34563 24395
rect 43545 24361 43579 24395
rect 44189 24361 44223 24395
rect 49065 24361 49099 24395
rect 49433 24361 49467 24395
rect 50997 24361 51031 24395
rect 51273 24361 51307 24395
rect 53941 24361 53975 24395
rect 56149 24361 56183 24395
rect 23305 24293 23339 24327
rect 29929 24293 29963 24327
rect 33793 24293 33827 24327
rect 36369 24293 36403 24327
rect 39221 24293 39255 24327
rect 40601 24293 40635 24327
rect 48053 24293 48087 24327
rect 19717 24225 19751 24259
rect 31401 24225 31435 24259
rect 34345 24225 34379 24259
rect 35081 24225 35115 24259
rect 35909 24225 35943 24259
rect 39865 24225 39899 24259
rect 41981 24225 42015 24259
rect 42257 24225 42291 24259
rect 43085 24225 43119 24259
rect 47225 24225 47259 24259
rect 49157 24225 49191 24259
rect 54125 24225 54159 24259
rect 56517 24225 56551 24259
rect 56609 24225 56643 24259
rect 19441 24157 19475 24191
rect 19533 24157 19567 24191
rect 19809 24157 19843 24191
rect 22385 24157 22419 24191
rect 22477 24157 22511 24191
rect 22753 24157 22787 24191
rect 23029 24157 23063 24191
rect 23121 24157 23155 24191
rect 23379 24157 23413 24191
rect 25145 24157 25179 24191
rect 25237 24157 25271 24191
rect 25421 24157 25455 24191
rect 25513 24157 25547 24191
rect 25606 24157 25640 24191
rect 25789 24157 25823 24191
rect 26019 24157 26053 24191
rect 28181 24157 28215 24191
rect 28273 24157 28307 24191
rect 28549 24157 28583 24191
rect 28825 24157 28859 24191
rect 29009 24157 29043 24191
rect 30108 24157 30142 24191
rect 30205 24157 30239 24191
rect 30425 24157 30459 24191
rect 30573 24157 30607 24191
rect 31033 24157 31067 24191
rect 33149 24157 33183 24191
rect 33242 24157 33276 24191
rect 33517 24157 33551 24191
rect 33655 24157 33689 24191
rect 34253 24157 34287 24191
rect 34529 24157 34563 24191
rect 36093 24157 36127 24191
rect 36185 24157 36219 24191
rect 36461 24157 36495 24191
rect 36737 24157 36771 24191
rect 36921 24157 36955 24191
rect 37105 24157 37139 24191
rect 39405 24157 39439 24191
rect 40325 24157 40359 24191
rect 41889 24157 41923 24191
rect 42073 24157 42107 24191
rect 42533 24157 42567 24191
rect 43361 24157 43395 24191
rect 46213 24157 46247 24191
rect 47409 24157 47443 24191
rect 47502 24157 47536 24191
rect 47874 24157 47908 24191
rect 49065 24157 49099 24191
rect 50721 24157 50755 24191
rect 50813 24157 50847 24191
rect 51089 24157 51123 24191
rect 51641 24157 51675 24191
rect 52193 24157 52227 24191
rect 53205 24157 53239 24191
rect 53573 24157 53607 24191
rect 54033 24157 54067 24191
rect 54309 24157 54343 24191
rect 54401 24157 54435 24191
rect 56333 24157 56367 24191
rect 57437 24157 57471 24191
rect 22569 24089 22603 24123
rect 25881 24089 25915 24123
rect 26341 24089 26375 24123
rect 28641 24089 28675 24123
rect 30297 24089 30331 24123
rect 33425 24089 33459 24123
rect 34713 24089 34747 24123
rect 35817 24089 35851 24123
rect 36829 24089 36863 24123
rect 40417 24089 40451 24123
rect 40785 24089 40819 24123
rect 42441 24089 42475 24123
rect 42993 24089 43027 24123
rect 43269 24089 43303 24123
rect 46397 24089 46431 24123
rect 47685 24089 47719 24123
rect 47777 24089 47811 24123
rect 53389 24089 53423 24123
rect 53481 24089 53515 24123
rect 19257 24021 19291 24055
rect 22201 24021 22235 24055
rect 26709 24021 26743 24055
rect 30665 24021 30699 24055
rect 30849 24021 30883 24055
rect 33977 24021 34011 24055
rect 36553 24021 36587 24055
rect 38761 24021 38795 24055
rect 43913 24021 43947 24055
rect 44833 24021 44867 24055
rect 48145 24021 48179 24055
rect 48421 24021 48455 24055
rect 50537 24021 50571 24055
rect 53757 24021 53791 24055
rect 54585 24021 54619 24055
rect 55781 24021 55815 24055
rect 57621 24021 57655 24055
rect 20085 23817 20119 23851
rect 23489 23817 23523 23851
rect 25053 23817 25087 23851
rect 25513 23817 25547 23851
rect 27261 23817 27295 23851
rect 33425 23817 33459 23851
rect 34805 23817 34839 23851
rect 34989 23817 35023 23851
rect 37013 23817 37047 23851
rect 45125 23817 45159 23851
rect 45293 23817 45327 23851
rect 46397 23817 46431 23851
rect 48789 23817 48823 23851
rect 49341 23817 49375 23851
rect 52193 23817 52227 23851
rect 55873 23817 55907 23851
rect 18521 23749 18555 23783
rect 20361 23749 20395 23783
rect 20453 23749 20487 23783
rect 22845 23749 22879 23783
rect 24777 23749 24811 23783
rect 26433 23749 26467 23783
rect 26525 23749 26559 23783
rect 27077 23749 27111 23783
rect 32413 23749 32447 23783
rect 33593 23749 33627 23783
rect 33793 23749 33827 23783
rect 34437 23749 34471 23783
rect 34529 23749 34563 23783
rect 36645 23749 36679 23783
rect 36829 23749 36863 23783
rect 38945 23749 38979 23783
rect 39497 23749 39531 23783
rect 39773 23749 39807 23783
rect 40509 23749 40543 23783
rect 42625 23749 42659 23783
rect 43177 23749 43211 23783
rect 43913 23749 43947 23783
rect 44925 23749 44959 23783
rect 45569 23749 45603 23783
rect 46673 23749 46707 23783
rect 48513 23749 48547 23783
rect 49985 23749 50019 23783
rect 50077 23749 50111 23783
rect 50721 23749 50755 23783
rect 53849 23749 53883 23783
rect 20269 23681 20303 23715
rect 20637 23681 20671 23715
rect 21557 23681 21591 23715
rect 22017 23681 22051 23715
rect 23029 23681 23063 23715
rect 23673 23681 23707 23715
rect 23765 23681 23799 23715
rect 23857 23681 23891 23715
rect 24041 23681 24075 23715
rect 24501 23681 24535 23715
rect 24685 23681 24719 23715
rect 24869 23681 24903 23715
rect 25237 23681 25271 23715
rect 25697 23681 25731 23715
rect 25789 23681 25823 23715
rect 25973 23681 26007 23715
rect 26065 23681 26099 23715
rect 26341 23681 26375 23715
rect 26709 23681 26743 23715
rect 27537 23681 27571 23715
rect 27721 23681 27755 23715
rect 27813 23681 27847 23715
rect 27905 23681 27939 23715
rect 28365 23681 28399 23715
rect 28457 23681 28491 23715
rect 28549 23681 28583 23715
rect 28733 23681 28767 23715
rect 32137 23681 32171 23715
rect 32321 23681 32355 23715
rect 32505 23681 32539 23715
rect 34253 23681 34287 23715
rect 34621 23681 34655 23715
rect 35168 23681 35202 23715
rect 35265 23681 35299 23715
rect 35357 23681 35391 23715
rect 35540 23681 35574 23715
rect 35633 23681 35667 23715
rect 38117 23681 38151 23715
rect 38209 23681 38243 23715
rect 39037 23681 39071 23715
rect 39865 23681 39899 23715
rect 42717 23681 42751 23715
rect 43361 23681 43395 23715
rect 44557 23681 44591 23715
rect 46535 23681 46569 23715
rect 46765 23681 46799 23715
rect 46948 23681 46982 23715
rect 47041 23681 47075 23715
rect 47593 23681 47627 23715
rect 47777 23681 47811 23715
rect 47869 23681 47903 23715
rect 47961 23681 47995 23715
rect 48237 23681 48271 23715
rect 48421 23681 48455 23715
rect 48605 23681 48639 23715
rect 49709 23681 49743 23715
rect 49857 23681 49891 23715
rect 50174 23681 50208 23715
rect 52745 23681 52779 23715
rect 52929 23681 52963 23715
rect 56241 23681 56275 23715
rect 56333 23681 56367 23715
rect 56977 23681 57011 23715
rect 58265 23681 58299 23715
rect 18245 23613 18279 23647
rect 36277 23613 36311 23647
rect 36553 23613 36587 23647
rect 42441 23613 42475 23647
rect 43269 23613 43303 23647
rect 44373 23613 44407 23647
rect 45753 23613 45787 23647
rect 48973 23613 49007 23647
rect 50445 23613 50479 23647
rect 54033 23613 54067 23647
rect 54309 23613 54343 23647
rect 56701 23613 56735 23647
rect 57529 23613 57563 23647
rect 26157 23545 26191 23579
rect 28089 23545 28123 23579
rect 28917 23545 28951 23579
rect 34069 23545 34103 23579
rect 40601 23545 40635 23579
rect 44097 23545 44131 23579
rect 45477 23545 45511 23579
rect 49525 23545 49559 23579
rect 50353 23545 50387 23579
rect 19993 23477 20027 23511
rect 25421 23477 25455 23511
rect 28181 23477 28215 23511
rect 29009 23477 29043 23511
rect 32689 23477 32723 23511
rect 33609 23477 33643 23511
rect 38393 23477 38427 23511
rect 38761 23477 38795 23511
rect 39589 23477 39623 23511
rect 40049 23477 40083 23511
rect 43545 23477 43579 23511
rect 44741 23477 44775 23511
rect 45109 23477 45143 23511
rect 47225 23477 47259 23511
rect 48145 23477 48179 23511
rect 53113 23477 53147 23511
rect 55781 23477 55815 23511
rect 56057 23477 56091 23511
rect 58449 23477 58483 23511
rect 21005 23273 21039 23307
rect 23857 23273 23891 23307
rect 29285 23273 29319 23307
rect 34943 23273 34977 23307
rect 39221 23273 39255 23307
rect 39681 23273 39715 23307
rect 40141 23273 40175 23307
rect 40509 23273 40543 23307
rect 41153 23273 41187 23307
rect 41705 23273 41739 23307
rect 43821 23273 43855 23307
rect 44281 23273 44315 23307
rect 44741 23273 44775 23307
rect 46673 23273 46707 23307
rect 49341 23273 49375 23307
rect 50905 23273 50939 23307
rect 54033 23273 54067 23307
rect 57437 23273 57471 23307
rect 38853 23205 38887 23239
rect 41797 23205 41831 23239
rect 43637 23205 43671 23239
rect 19257 23137 19291 23171
rect 21557 23137 21591 23171
rect 22109 23137 22143 23171
rect 22385 23137 22419 23171
rect 32321 23137 32355 23171
rect 32873 23137 32907 23171
rect 36737 23137 36771 23171
rect 38301 23137 38335 23171
rect 39865 23137 39899 23171
rect 42533 23137 42567 23171
rect 44833 23137 44867 23171
rect 45753 23137 45787 23171
rect 48421 23137 48455 23171
rect 55965 23137 55999 23171
rect 18153 23069 18187 23103
rect 21465 23069 21499 23103
rect 21741 23069 21775 23103
rect 21833 23069 21867 23103
rect 25789 23069 25823 23103
rect 26065 23069 26099 23103
rect 26157 23069 26191 23103
rect 27537 23069 27571 23103
rect 31953 23069 31987 23103
rect 32413 23069 32447 23103
rect 32597 23069 32631 23103
rect 32689 23069 32723 23103
rect 32965 23069 32999 23103
rect 36369 23069 36403 23103
rect 38485 23069 38519 23103
rect 39497 23069 39531 23103
rect 39681 23069 39715 23103
rect 39957 23069 39991 23103
rect 41429 23069 41463 23103
rect 41613 23069 41647 23103
rect 41889 23069 41923 23103
rect 42625 23069 42659 23103
rect 43177 23069 43211 23103
rect 43453 23069 43487 23103
rect 44557 23069 44591 23103
rect 45196 23069 45230 23103
rect 45568 23069 45602 23103
rect 45661 23069 45695 23103
rect 46305 23069 46339 23103
rect 48789 23069 48823 23103
rect 49157 23069 49191 23103
rect 49433 23069 49467 23103
rect 50353 23069 50387 23103
rect 50629 23069 50663 23103
rect 50721 23069 50755 23103
rect 53665 23069 53699 23103
rect 54217 23069 54251 23103
rect 55689 23069 55723 23103
rect 19533 23001 19567 23035
rect 25973 23001 26007 23035
rect 27813 23001 27847 23035
rect 39221 23001 39255 23035
rect 42165 23001 42199 23035
rect 43085 23001 43119 23035
rect 45293 23001 45327 23035
rect 45385 23001 45419 23035
rect 48145 23001 48179 23035
rect 48973 23001 49007 23035
rect 49065 23001 49099 23035
rect 50537 23001 50571 23035
rect 53389 23001 53423 23035
rect 54953 23001 54987 23035
rect 22017 22933 22051 22967
rect 26341 22933 26375 22967
rect 30527 22933 30561 22967
rect 38669 22933 38703 22967
rect 39405 22933 39439 22967
rect 41245 22933 41279 22967
rect 43269 22933 43303 22967
rect 43913 22933 43947 22967
rect 44373 22933 44407 22967
rect 45017 22933 45051 22967
rect 48605 22933 48639 22967
rect 51917 22933 51951 22967
rect 19441 22729 19475 22763
rect 23581 22729 23615 22763
rect 28089 22729 28123 22763
rect 36185 22729 36219 22763
rect 37841 22729 37875 22763
rect 38853 22729 38887 22763
rect 39405 22729 39439 22763
rect 42441 22729 42475 22763
rect 48881 22729 48915 22763
rect 49065 22729 49099 22763
rect 49617 22729 49651 22763
rect 54033 22729 54067 22763
rect 19073 22661 19107 22695
rect 28733 22661 28767 22695
rect 35817 22661 35851 22695
rect 35909 22661 35943 22695
rect 38301 22661 38335 22695
rect 42809 22661 42843 22695
rect 44373 22661 44407 22695
rect 18337 22593 18371 22627
rect 19804 22593 19838 22627
rect 19901 22593 19935 22627
rect 19993 22593 20027 22627
rect 20121 22593 20155 22627
rect 20269 22593 20303 22627
rect 21833 22593 21867 22627
rect 25789 22593 25823 22627
rect 26065 22593 26099 22627
rect 26157 22593 26191 22627
rect 28273 22593 28307 22627
rect 28365 22593 28399 22627
rect 28641 22593 28675 22627
rect 32321 22593 32355 22627
rect 32413 22593 32447 22627
rect 32689 22593 32723 22627
rect 32781 22593 32815 22627
rect 35173 22593 35207 22627
rect 35541 22593 35575 22627
rect 35633 22593 35667 22627
rect 36001 22593 36035 22627
rect 36277 22593 36311 22627
rect 36553 22593 36587 22627
rect 36645 22593 36679 22627
rect 38117 22593 38151 22627
rect 38393 22593 38427 22627
rect 39313 22593 39347 22627
rect 39589 22593 39623 22627
rect 41337 22593 41371 22627
rect 41429 22593 41463 22627
rect 41705 22593 41739 22627
rect 41797 22593 41831 22627
rect 42625 22593 42659 22627
rect 42717 22593 42751 22627
rect 42993 22593 43027 22627
rect 47593 22593 47627 22627
rect 48237 22593 48271 22627
rect 48329 22593 48363 22627
rect 48605 22593 48639 22627
rect 48697 22593 48731 22627
rect 49249 22593 49283 22627
rect 49341 22593 49375 22627
rect 52745 22593 52779 22627
rect 53389 22593 53423 22627
rect 53481 22593 53515 22627
rect 53757 22593 53791 22627
rect 53849 22593 53883 22627
rect 56149 22593 56183 22627
rect 58265 22593 58299 22627
rect 22109 22525 22143 22559
rect 34989 22525 35023 22559
rect 36369 22525 36403 22559
rect 44097 22525 44131 22559
rect 47409 22525 47443 22559
rect 54125 22525 54159 22559
rect 55873 22525 55907 22559
rect 25881 22457 25915 22491
rect 28549 22457 28583 22491
rect 41061 22457 41095 22491
rect 43177 22457 43211 22491
rect 58449 22457 58483 22491
rect 19625 22389 19659 22423
rect 20453 22389 20487 22423
rect 26341 22389 26375 22423
rect 32137 22389 32171 22423
rect 32597 22389 32631 22423
rect 32965 22389 32999 22423
rect 36829 22389 36863 22423
rect 37933 22389 37967 22423
rect 39773 22389 39807 22423
rect 39865 22389 39899 22423
rect 41153 22389 41187 22423
rect 41613 22389 41647 22423
rect 45845 22389 45879 22423
rect 48421 22389 48455 22423
rect 53573 22389 53607 22423
rect 54401 22389 54435 22423
rect 18613 22185 18647 22219
rect 25605 22185 25639 22219
rect 27089 22185 27123 22219
rect 33011 22185 33045 22219
rect 35633 22185 35667 22219
rect 36231 22185 36265 22219
rect 40680 22185 40714 22219
rect 49709 22185 49743 22219
rect 33149 22117 33183 22151
rect 47777 22117 47811 22151
rect 27353 22049 27387 22083
rect 31585 22049 31619 22083
rect 38025 22049 38059 22083
rect 50261 22049 50295 22083
rect 53113 22049 53147 22083
rect 18797 21981 18831 22015
rect 18981 21981 19015 22015
rect 19073 21981 19107 22015
rect 19901 21981 19935 22015
rect 23581 21981 23615 22015
rect 27905 21981 27939 22015
rect 29561 21981 29595 22015
rect 31217 21981 31251 22015
rect 33333 21981 33367 22015
rect 33517 21981 33551 22015
rect 33609 21981 33643 22015
rect 35357 21981 35391 22015
rect 35449 21981 35483 22015
rect 35725 21981 35759 22015
rect 35817 21981 35851 22015
rect 37657 21981 37691 22015
rect 40417 21981 40451 22015
rect 45017 21981 45051 22015
rect 45201 21981 45235 22015
rect 47409 21981 47443 22015
rect 47593 21981 47627 22015
rect 48145 21981 48179 22015
rect 48329 21981 48363 22015
rect 48513 21981 48547 22015
rect 48973 21981 49007 22015
rect 49157 21981 49191 22015
rect 49525 21981 49559 22015
rect 52377 21981 52411 22015
rect 54033 21981 54067 22015
rect 56885 21981 56919 22015
rect 19809 21913 19843 21947
rect 27537 21913 27571 21947
rect 27997 21913 28031 21947
rect 48237 21913 48271 21947
rect 52561 21913 52595 21947
rect 52837 21913 52871 21947
rect 55413 21913 55447 21947
rect 55689 21913 55723 21947
rect 57152 21913 57186 21947
rect 20085 21845 20119 21879
rect 20361 21845 20395 21879
rect 23765 21845 23799 21879
rect 29745 21845 29779 21879
rect 35081 21845 35115 21879
rect 35173 21845 35207 21879
rect 36001 21845 36035 21879
rect 42165 21845 42199 21879
rect 42349 21845 42383 21879
rect 45385 21845 45419 21879
rect 47961 21845 47995 21879
rect 48881 21845 48915 21879
rect 49341 21845 49375 21879
rect 50905 21845 50939 21879
rect 52193 21845 52227 21879
rect 52653 21845 52687 21879
rect 53389 21845 53423 21879
rect 55505 21845 55539 21879
rect 58265 21845 58299 21879
rect 19441 21641 19475 21675
rect 20177 21641 20211 21675
rect 20913 21641 20947 21675
rect 26065 21641 26099 21675
rect 30665 21641 30699 21675
rect 31033 21641 31067 21675
rect 32689 21641 32723 21675
rect 32965 21641 32999 21675
rect 34713 21641 34747 21675
rect 46029 21641 46063 21675
rect 55781 21641 55815 21675
rect 57529 21641 57563 21675
rect 19809 21573 19843 21607
rect 20545 21573 20579 21607
rect 23673 21573 23707 21607
rect 32413 21573 32447 21607
rect 47409 21573 47443 21607
rect 52561 21573 52595 21607
rect 53021 21573 53055 21607
rect 54769 21573 54803 21607
rect 55965 21573 55999 21607
rect 56701 21573 56735 21607
rect 19073 21505 19107 21539
rect 19620 21505 19654 21539
rect 19717 21505 19751 21539
rect 19992 21505 20026 21539
rect 20085 21505 20119 21539
rect 20361 21505 20395 21539
rect 20453 21505 20487 21539
rect 20729 21505 20763 21539
rect 23576 21505 23610 21539
rect 23765 21505 23799 21539
rect 23948 21505 23982 21539
rect 24041 21505 24075 21539
rect 24133 21505 24167 21539
rect 24501 21505 24535 21539
rect 24869 21505 24903 21539
rect 26249 21505 26283 21539
rect 26341 21505 26375 21539
rect 26617 21505 26651 21539
rect 26985 21505 27019 21539
rect 29469 21505 29503 21539
rect 29561 21505 29595 21539
rect 29837 21505 29871 21539
rect 29929 21505 29963 21539
rect 30481 21505 30515 21539
rect 30849 21505 30883 21539
rect 31585 21505 31619 21539
rect 31677 21505 31711 21539
rect 31953 21505 31987 21539
rect 32137 21505 32171 21539
rect 32321 21505 32355 21539
rect 32505 21505 32539 21539
rect 32781 21505 32815 21539
rect 34069 21505 34103 21539
rect 34162 21505 34196 21539
rect 34345 21505 34379 21539
rect 34437 21505 34471 21539
rect 34534 21505 34568 21539
rect 35173 21505 35207 21539
rect 41889 21505 41923 21539
rect 41981 21505 42015 21539
rect 42257 21505 42291 21539
rect 46765 21505 46799 21539
rect 47593 21505 47627 21539
rect 52101 21505 52135 21539
rect 52377 21505 52411 21539
rect 54585 21505 54619 21539
rect 54861 21505 54895 21539
rect 54953 21505 54987 21539
rect 55229 21505 55263 21539
rect 55505 21505 55539 21539
rect 55597 21505 55631 21539
rect 56149 21505 56183 21539
rect 56885 21505 56919 21539
rect 57069 21505 57103 21539
rect 57161 21505 57195 21539
rect 57253 21505 57287 21539
rect 57897 21505 57931 21539
rect 58449 21505 58483 21539
rect 19349 21437 19383 21471
rect 26801 21437 26835 21471
rect 27261 21437 27295 21471
rect 28825 21437 28859 21471
rect 34805 21437 34839 21471
rect 44281 21437 44315 21471
rect 44557 21437 44591 21471
rect 47869 21437 47903 21471
rect 49985 21437 50019 21471
rect 50261 21437 50295 21471
rect 51733 21437 51767 21471
rect 52009 21437 52043 21471
rect 52745 21437 52779 21471
rect 26433 21369 26467 21403
rect 41613 21369 41647 21403
rect 42165 21369 42199 21403
rect 55137 21369 55171 21403
rect 18889 21301 18923 21335
rect 19257 21301 19291 21335
rect 23397 21301 23431 21335
rect 24317 21301 24351 21335
rect 24685 21301 24719 21335
rect 25881 21301 25915 21335
rect 28733 21301 28767 21335
rect 29653 21301 29687 21335
rect 30113 21301 30147 21335
rect 31401 21301 31435 21335
rect 31861 21301 31895 21335
rect 36599 21301 36633 21335
rect 41705 21301 41739 21335
rect 46121 21301 46155 21335
rect 49341 21301 49375 21335
rect 49433 21301 49467 21335
rect 52193 21301 52227 21335
rect 54493 21301 54527 21335
rect 55321 21301 55355 21335
rect 56333 21301 56367 21335
rect 25145 21097 25179 21131
rect 25881 21097 25915 21131
rect 26065 21097 26099 21131
rect 29119 21097 29153 21131
rect 33011 21097 33045 21131
rect 35633 21097 35667 21131
rect 36277 21097 36311 21131
rect 36645 21097 36679 21131
rect 43177 21097 43211 21131
rect 45017 21097 45051 21131
rect 45477 21097 45511 21131
rect 45661 21097 45695 21131
rect 47501 21097 47535 21131
rect 47961 21097 47995 21131
rect 49801 21097 49835 21131
rect 50905 21097 50939 21131
rect 51273 21097 51307 21131
rect 52469 21097 52503 21131
rect 18981 21029 19015 21063
rect 26893 21029 26927 21063
rect 44005 21029 44039 21063
rect 44741 21029 44775 21063
rect 50169 21029 50203 21063
rect 19257 20961 19291 20995
rect 22293 20961 22327 20995
rect 22477 20961 22511 20995
rect 24225 20961 24259 20995
rect 24961 20961 24995 20995
rect 30021 20961 30055 20995
rect 31585 20961 31619 20995
rect 39681 20961 39715 20995
rect 40417 20961 40451 20995
rect 41153 20961 41187 20995
rect 46765 20961 46799 20995
rect 51365 20961 51399 20995
rect 58081 20961 58115 20995
rect 18705 20893 18739 20927
rect 18797 20893 18831 20927
rect 19073 20893 19107 20927
rect 22017 20893 22051 20927
rect 22109 20893 22143 20927
rect 22385 20893 22419 20927
rect 25329 20893 25363 20927
rect 25697 20893 25731 20927
rect 26203 20893 26237 20927
rect 26433 20893 26467 20927
rect 26616 20893 26650 20927
rect 26709 20893 26743 20927
rect 27077 20893 27111 20927
rect 29377 20893 29411 20927
rect 29745 20893 29779 20927
rect 29837 20893 29871 20927
rect 30113 20893 30147 20927
rect 30481 20893 30515 20927
rect 31033 20893 31067 20927
rect 31217 20893 31251 20927
rect 35081 20893 35115 20927
rect 35357 20893 35391 20927
rect 35449 20893 35483 20927
rect 37933 20893 37967 20927
rect 40877 20893 40911 20927
rect 42901 20893 42935 20927
rect 44097 20893 44131 20927
rect 44245 20893 44279 20927
rect 44465 20893 44499 20927
rect 44603 20893 44637 20927
rect 45201 20893 45235 20927
rect 45293 20893 45327 20927
rect 45569 20893 45603 20927
rect 46857 20893 46891 20927
rect 47133 20893 47167 20927
rect 47225 20893 47259 20927
rect 47685 20893 47719 20927
rect 47777 20893 47811 20927
rect 48053 20893 48087 20927
rect 48600 20893 48634 20927
rect 48697 20893 48731 20927
rect 48789 20893 48823 20927
rect 48972 20893 49006 20927
rect 49065 20893 49099 20927
rect 49157 20893 49191 20927
rect 49305 20893 49339 20927
rect 49433 20893 49467 20927
rect 49525 20893 49559 20927
rect 49663 20893 49697 20927
rect 50307 20893 50341 20927
rect 50537 20893 50571 20927
rect 50665 20893 50699 20927
rect 50813 20893 50847 20927
rect 51089 20893 51123 20927
rect 51825 20893 51859 20927
rect 51918 20893 51952 20927
rect 52101 20893 52135 20927
rect 52193 20893 52227 20927
rect 52331 20893 52365 20927
rect 55689 20893 55723 20927
rect 56057 20893 56091 20927
rect 18521 20825 18555 20859
rect 19533 20825 19567 20859
rect 22753 20825 22787 20859
rect 24409 20825 24443 20859
rect 25421 20825 25455 20859
rect 25513 20825 25547 20859
rect 26341 20825 26375 20859
rect 35265 20825 35299 20859
rect 36369 20825 36403 20859
rect 36829 20825 36863 20859
rect 38209 20825 38243 20859
rect 42717 20825 42751 20859
rect 44373 20825 44407 20859
rect 47041 20825 47075 20859
rect 50445 20825 50479 20859
rect 55873 20825 55907 20859
rect 55965 20825 55999 20859
rect 57805 20825 57839 20859
rect 21005 20757 21039 20791
rect 21833 20757 21867 20791
rect 27629 20757 27663 20791
rect 29561 20757 29595 20791
rect 34805 20757 34839 20791
rect 39865 20757 39899 20791
rect 42625 20757 42659 20791
rect 45937 20757 45971 20791
rect 46581 20757 46615 20791
rect 47409 20757 47443 20791
rect 48145 20757 48179 20791
rect 48421 20757 48455 20791
rect 49893 20757 49927 20791
rect 55045 20757 55079 20791
rect 56241 20757 56275 20791
rect 56333 20757 56367 20791
rect 20453 20553 20487 20587
rect 23673 20553 23707 20587
rect 25145 20553 25179 20587
rect 26433 20553 26467 20587
rect 28825 20553 28859 20587
rect 36645 20553 36679 20587
rect 38485 20553 38519 20587
rect 43085 20553 43119 20587
rect 45385 20553 45419 20587
rect 47133 20553 47167 20587
rect 47317 20553 47351 20587
rect 49617 20553 49651 20587
rect 56793 20553 56827 20587
rect 20729 20485 20763 20519
rect 20913 20485 20947 20519
rect 24501 20485 24535 20519
rect 25697 20485 25731 20519
rect 28457 20485 28491 20519
rect 28549 20485 28583 20519
rect 29285 20485 29319 20519
rect 29929 20485 29963 20519
rect 39129 20485 39163 20519
rect 42809 20485 42843 20519
rect 44925 20485 44959 20519
rect 45017 20485 45051 20519
rect 47961 20485 47995 20519
rect 48605 20485 48639 20519
rect 49893 20485 49927 20519
rect 50169 20485 50203 20519
rect 18521 20417 18555 20451
rect 21833 20417 21867 20451
rect 23857 20417 23891 20451
rect 24041 20417 24075 20451
rect 24133 20417 24167 20451
rect 24225 20417 24259 20451
rect 24409 20417 24443 20451
rect 24593 20417 24627 20451
rect 25421 20417 25455 20451
rect 25514 20417 25548 20451
rect 25789 20417 25823 20451
rect 25927 20417 25961 20451
rect 26157 20417 26191 20451
rect 28273 20417 28307 20451
rect 28641 20417 28675 20451
rect 29101 20417 29135 20451
rect 29377 20417 29411 20451
rect 35817 20417 35851 20451
rect 36461 20417 36495 20451
rect 38669 20417 38703 20451
rect 38761 20417 38795 20451
rect 39037 20417 39071 20451
rect 39313 20417 39347 20451
rect 42625 20417 42659 20451
rect 42717 20417 42751 20451
rect 42993 20417 43027 20451
rect 43269 20417 43303 20451
rect 43361 20417 43395 20451
rect 43453 20417 43487 20451
rect 43637 20417 43671 20451
rect 44787 20417 44821 20451
rect 45200 20417 45234 20451
rect 45293 20417 45327 20451
rect 47593 20417 47627 20451
rect 47741 20417 47775 20451
rect 47869 20417 47903 20451
rect 48058 20417 48092 20451
rect 48329 20417 48363 20451
rect 48422 20417 48456 20451
rect 48697 20417 48731 20451
rect 48813 20417 48847 20451
rect 49065 20417 49099 20451
rect 49341 20417 49375 20451
rect 50077 20417 50111 20451
rect 53665 20417 53699 20451
rect 55413 20417 55447 20451
rect 56241 20417 56275 20451
rect 56517 20417 56551 20451
rect 56609 20417 56643 20451
rect 18797 20349 18831 20383
rect 20269 20349 20303 20383
rect 22109 20349 22143 20383
rect 23581 20349 23615 20383
rect 28917 20349 28951 20383
rect 29653 20349 29687 20383
rect 31401 20349 31435 20383
rect 33609 20349 33643 20383
rect 33977 20349 34011 20383
rect 35403 20349 35437 20383
rect 35541 20349 35575 20383
rect 39497 20349 39531 20383
rect 40509 20349 40543 20383
rect 40785 20349 40819 20383
rect 49249 20349 49283 20383
rect 53941 20349 53975 20383
rect 55137 20349 55171 20383
rect 42257 20281 42291 20315
rect 44557 20281 44591 20315
rect 48237 20281 48271 20315
rect 49525 20281 49559 20315
rect 56333 20281 56367 20315
rect 24777 20213 24811 20247
rect 24961 20213 24995 20247
rect 26065 20213 26099 20247
rect 36829 20213 36863 20247
rect 38945 20213 38979 20247
rect 39681 20213 39715 20247
rect 42441 20213 42475 20247
rect 44649 20213 44683 20247
rect 45569 20213 45603 20247
rect 48973 20213 49007 20247
rect 49065 20213 49099 20247
rect 53113 20213 53147 20247
rect 53481 20213 53515 20247
rect 53849 20213 53883 20247
rect 55229 20213 55263 20247
rect 55597 20213 55631 20247
rect 56057 20213 56091 20247
rect 25421 20009 25455 20043
rect 25605 20009 25639 20043
rect 26617 20009 26651 20043
rect 27353 20009 27387 20043
rect 33977 20009 34011 20043
rect 34713 20009 34747 20043
rect 35173 20009 35207 20043
rect 36737 20009 36771 20043
rect 41245 20009 41279 20043
rect 41337 20009 41371 20043
rect 47961 20009 47995 20043
rect 48881 20009 48915 20043
rect 50537 20009 50571 20043
rect 53941 20009 53975 20043
rect 55137 20009 55171 20043
rect 57069 20009 57103 20043
rect 26525 19941 26559 19975
rect 33793 19941 33827 19975
rect 35357 19941 35391 19975
rect 41797 19941 41831 19975
rect 25697 19873 25731 19907
rect 26709 19873 26743 19907
rect 30849 19873 30883 19907
rect 31861 19873 31895 19907
rect 37105 19873 37139 19907
rect 44833 19873 44867 19907
rect 48697 19873 48731 19907
rect 51457 19873 51491 19907
rect 55321 19873 55355 19907
rect 1685 19805 1719 19839
rect 24869 19805 24903 19839
rect 25053 19805 25087 19839
rect 25237 19805 25271 19839
rect 25881 19805 25915 19839
rect 26029 19805 26063 19839
rect 26157 19805 26191 19839
rect 26346 19805 26380 19839
rect 26893 19805 26927 19839
rect 31265 19805 31299 19839
rect 31401 19805 31435 19839
rect 31621 19805 31655 19839
rect 31769 19805 31803 19839
rect 34161 19805 34195 19839
rect 34345 19805 34379 19839
rect 34529 19805 34563 19839
rect 34897 19805 34931 19839
rect 34989 19805 35023 19839
rect 35265 19805 35299 19839
rect 35541 19805 35575 19839
rect 35725 19805 35759 19839
rect 35909 19805 35943 19839
rect 36185 19805 36219 19839
rect 36553 19805 36587 19839
rect 36921 19805 36955 19839
rect 39497 19805 39531 19839
rect 41521 19805 41555 19839
rect 41613 19805 41647 19839
rect 41889 19805 41923 19839
rect 45201 19805 45235 19839
rect 45385 19805 45419 19839
rect 45477 19805 45511 19839
rect 47409 19805 47443 19839
rect 47777 19805 47811 19839
rect 48053 19805 48087 19839
rect 48329 19805 48363 19839
rect 48421 19805 48455 19839
rect 49065 19805 49099 19839
rect 49157 19805 49191 19839
rect 49433 19805 49467 19839
rect 50721 19805 50755 19839
rect 50814 19805 50848 19839
rect 50997 19805 51031 19839
rect 51186 19805 51220 19839
rect 53297 19805 53331 19839
rect 53390 19805 53424 19839
rect 53665 19805 53699 19839
rect 53762 19805 53796 19839
rect 54493 19805 54527 19839
rect 54586 19805 54620 19839
rect 54958 19805 54992 19839
rect 57897 19805 57931 19839
rect 58265 19805 58299 19839
rect 25145 19737 25179 19771
rect 26249 19737 26283 19771
rect 26617 19737 26651 19771
rect 30021 19737 30055 19771
rect 31493 19737 31527 19771
rect 34253 19737 34287 19771
rect 35633 19737 35667 19771
rect 36277 19737 36311 19771
rect 36369 19737 36403 19771
rect 37381 19737 37415 19771
rect 44557 19737 44591 19771
rect 45017 19737 45051 19771
rect 45569 19737 45603 19771
rect 47593 19737 47627 19771
rect 47685 19737 47719 19771
rect 48237 19737 48271 19771
rect 49249 19737 49283 19771
rect 51089 19737 51123 19771
rect 51733 19737 51767 19771
rect 53573 19737 53607 19771
rect 54769 19737 54803 19771
rect 54861 19737 54895 19771
rect 55597 19737 55631 19771
rect 1501 19669 1535 19703
rect 27077 19669 27111 19703
rect 27169 19669 27203 19703
rect 29837 19669 29871 19703
rect 31125 19669 31159 19703
rect 32137 19669 32171 19703
rect 36001 19669 36035 19703
rect 38853 19669 38887 19703
rect 38945 19669 38979 19703
rect 43085 19669 43119 19703
rect 46857 19669 46891 19703
rect 48605 19669 48639 19703
rect 49525 19669 49559 19703
rect 49801 19669 49835 19703
rect 51365 19669 51399 19703
rect 53205 19669 53239 19703
rect 58081 19669 58115 19703
rect 58449 19669 58483 19703
rect 15025 19465 15059 19499
rect 19441 19465 19475 19499
rect 22477 19465 22511 19499
rect 26617 19465 26651 19499
rect 28641 19465 28675 19499
rect 28917 19465 28951 19499
rect 38945 19465 38979 19499
rect 44925 19465 44959 19499
rect 46397 19465 46431 19499
rect 52929 19465 52963 19499
rect 55137 19465 55171 19499
rect 56701 19465 56735 19499
rect 19717 19397 19751 19431
rect 28273 19397 28307 19431
rect 28365 19397 28399 19431
rect 40785 19397 40819 19431
rect 46673 19397 46707 19431
rect 46765 19397 46799 19431
rect 52837 19397 52871 19431
rect 16138 19329 16172 19363
rect 16405 19329 16439 19363
rect 18981 19329 19015 19363
rect 19073 19329 19107 19363
rect 19349 19329 19383 19363
rect 19625 19329 19659 19363
rect 19809 19329 19843 19363
rect 19993 19329 20027 19363
rect 22000 19329 22034 19363
rect 22169 19329 22203 19363
rect 22385 19329 22419 19363
rect 23029 19329 23063 19363
rect 23121 19329 23155 19363
rect 23397 19329 23431 19363
rect 26341 19329 26375 19363
rect 26525 19329 26559 19363
rect 27997 19329 28031 19363
rect 28145 19329 28179 19363
rect 28503 19329 28537 19363
rect 28733 19329 28767 19363
rect 31125 19329 31159 19363
rect 31217 19329 31251 19363
rect 31493 19329 31527 19363
rect 34161 19329 34195 19363
rect 35955 19329 35989 19363
rect 38117 19329 38151 19363
rect 38209 19329 38243 19363
rect 38485 19329 38519 19363
rect 39129 19329 39163 19363
rect 39221 19329 39255 19363
rect 39313 19329 39347 19363
rect 39497 19329 39531 19363
rect 40417 19329 40451 19363
rect 45201 19329 45235 19363
rect 45385 19329 45419 19363
rect 46213 19329 46247 19363
rect 46576 19329 46610 19363
rect 46948 19329 46982 19363
rect 47041 19329 47075 19363
rect 48605 19329 48639 19363
rect 48697 19329 48731 19363
rect 48973 19329 49007 19363
rect 49065 19329 49099 19363
rect 53389 19329 53423 19363
rect 56793 19329 56827 19363
rect 56977 19329 57011 19363
rect 57069 19329 57103 19363
rect 57161 19329 57195 19363
rect 57897 19329 57931 19363
rect 24593 19261 24627 19295
rect 34529 19261 34563 19295
rect 37933 19261 37967 19295
rect 41521 19261 41555 19295
rect 44373 19261 44407 19295
rect 45477 19261 45511 19295
rect 48053 19261 48087 19295
rect 49709 19261 49743 19295
rect 49985 19261 50019 19295
rect 51457 19261 51491 19295
rect 52101 19261 52135 19295
rect 53665 19261 53699 19295
rect 58449 19261 58483 19295
rect 20085 19193 20119 19227
rect 23305 19193 23339 19227
rect 23581 19193 23615 19227
rect 41889 19193 41923 19227
rect 47317 19193 47351 19227
rect 47777 19193 47811 19227
rect 48789 19193 48823 19227
rect 18797 19125 18831 19159
rect 19257 19125 19291 19159
rect 21833 19125 21867 19159
rect 22293 19125 22327 19159
rect 22845 19125 22879 19159
rect 26985 19125 27019 19159
rect 30941 19125 30975 19159
rect 31401 19125 31435 19159
rect 38393 19125 38427 19159
rect 45017 19125 45051 19159
rect 47133 19125 47167 19159
rect 47593 19125 47627 19159
rect 49249 19125 49283 19159
rect 51549 19125 51583 19159
rect 57437 19125 57471 19159
rect 16129 18921 16163 18955
rect 16865 18921 16899 18955
rect 25053 18921 25087 18955
rect 25881 18921 25915 18955
rect 30573 18921 30607 18955
rect 34529 18921 34563 18955
rect 34897 18921 34931 18955
rect 39681 18921 39715 18955
rect 46765 18921 46799 18955
rect 47133 18921 47167 18955
rect 50169 18921 50203 18955
rect 51641 18921 51675 18955
rect 53205 18921 53239 18955
rect 58265 18921 58299 18955
rect 49525 18853 49559 18887
rect 50629 18853 50663 18887
rect 15393 18785 15427 18819
rect 17601 18785 17635 18819
rect 19073 18785 19107 18819
rect 21925 18785 21959 18819
rect 22569 18785 22603 18819
rect 24041 18785 24075 18819
rect 27629 18785 27663 18819
rect 32413 18785 32447 18819
rect 34069 18785 34103 18819
rect 37933 18785 37967 18819
rect 45293 18785 45327 18819
rect 48605 18785 48639 18819
rect 48881 18785 48915 18819
rect 52009 18785 52043 18819
rect 16037 18717 16071 18751
rect 16405 18717 16439 18751
rect 16497 18717 16531 18751
rect 16589 18717 16623 18751
rect 16773 18717 16807 18751
rect 17325 18717 17359 18751
rect 19625 18717 19659 18751
rect 19718 18717 19752 18751
rect 20090 18717 20124 18751
rect 22201 18717 22235 18751
rect 22293 18717 22327 18751
rect 24501 18717 24535 18751
rect 24685 18717 24719 18751
rect 24869 18717 24903 18751
rect 25237 18717 25271 18751
rect 25330 18717 25364 18751
rect 25513 18717 25547 18751
rect 25702 18717 25736 18751
rect 25973 18717 26007 18751
rect 26111 18717 26145 18751
rect 26438 18717 26472 18751
rect 26985 18717 27019 18751
rect 27261 18717 27295 18751
rect 27353 18717 27387 18751
rect 30021 18717 30055 18751
rect 30205 18717 30239 18751
rect 30297 18717 30331 18751
rect 30389 18717 30423 18751
rect 33977 18717 34011 18751
rect 34253 18717 34287 18751
rect 34345 18717 34379 18751
rect 35173 18717 35207 18751
rect 37105 18717 37139 18751
rect 40417 18717 40451 18751
rect 45017 18717 45051 18751
rect 48973 18717 49007 18751
rect 49341 18717 49375 18751
rect 50353 18717 50387 18751
rect 50445 18717 50479 18751
rect 50721 18717 50755 18751
rect 51825 18717 51859 18751
rect 52101 18717 52135 18751
rect 56885 18717 56919 18751
rect 57152 18717 57186 18751
rect 19901 18649 19935 18683
rect 19993 18649 20027 18683
rect 24777 18649 24811 18683
rect 25605 18649 25639 18683
rect 26249 18649 26283 18683
rect 26341 18649 26375 18683
rect 27169 18649 27203 18683
rect 27905 18649 27939 18683
rect 32137 18649 32171 18683
rect 36737 18649 36771 18683
rect 38209 18649 38243 18683
rect 39865 18649 39899 18683
rect 49157 18649 49191 18683
rect 49249 18649 49283 18683
rect 20269 18581 20303 18615
rect 20453 18581 20487 18615
rect 26617 18581 26651 18615
rect 26801 18581 26835 18615
rect 27537 18581 27571 18615
rect 29377 18581 29411 18615
rect 30665 18581 30699 18615
rect 36829 18581 36863 18615
rect 19993 18377 20027 18411
rect 21925 18377 21959 18411
rect 23213 18377 23247 18411
rect 24961 18377 24995 18411
rect 30941 18377 30975 18411
rect 32137 18377 32171 18411
rect 37105 18377 37139 18411
rect 38301 18377 38335 18411
rect 40417 18377 40451 18411
rect 41153 18377 41187 18411
rect 42993 18377 43027 18411
rect 45569 18377 45603 18411
rect 56701 18377 56735 18411
rect 37933 18309 37967 18343
rect 39037 18309 39071 18343
rect 39957 18309 39991 18343
rect 40785 18309 40819 18343
rect 50169 18309 50203 18343
rect 16681 18241 16715 18275
rect 17693 18241 17727 18275
rect 20269 18241 20303 18275
rect 20545 18241 20579 18275
rect 22085 18241 22119 18275
rect 22201 18241 22235 18275
rect 22293 18241 22327 18275
rect 22477 18241 22511 18275
rect 23397 18241 23431 18275
rect 23489 18241 23523 18275
rect 23581 18241 23615 18275
rect 23765 18241 23799 18275
rect 27997 18241 28031 18275
rect 28181 18241 28215 18275
rect 28273 18241 28307 18275
rect 28549 18241 28583 18275
rect 28825 18241 28859 18275
rect 30297 18241 30331 18275
rect 30390 18241 30424 18275
rect 30573 18241 30607 18275
rect 30665 18241 30699 18275
rect 30762 18241 30796 18275
rect 32321 18241 32355 18275
rect 32505 18241 32539 18275
rect 37749 18241 37783 18275
rect 38025 18241 38059 18275
rect 38117 18241 38151 18275
rect 38393 18241 38427 18275
rect 38577 18241 38611 18275
rect 38669 18241 38703 18275
rect 38761 18241 38795 18275
rect 39221 18241 39255 18275
rect 39313 18241 39347 18275
rect 39589 18241 39623 18275
rect 39681 18241 39715 18275
rect 39774 18241 39808 18275
rect 40049 18241 40083 18275
rect 40146 18241 40180 18275
rect 40601 18241 40635 18275
rect 40877 18241 40911 18275
rect 40969 18241 41003 18275
rect 41245 18241 41279 18275
rect 41521 18241 41555 18275
rect 41613 18241 41647 18275
rect 46213 18241 46247 18275
rect 49985 18241 50019 18275
rect 50261 18241 50295 18275
rect 50353 18241 50387 18275
rect 52929 18241 52963 18275
rect 53021 18241 53055 18275
rect 53297 18241 53331 18275
rect 53757 18241 53791 18275
rect 56793 18241 56827 18275
rect 56977 18241 57011 18275
rect 57069 18241 57103 18275
rect 57161 18241 57195 18275
rect 57897 18241 57931 18275
rect 58449 18241 58483 18275
rect 17417 18173 17451 18207
rect 18245 18173 18279 18207
rect 18521 18173 18555 18207
rect 20085 18173 20119 18207
rect 25053 18173 25087 18207
rect 26525 18173 26559 18207
rect 26801 18173 26835 18207
rect 28641 18173 28675 18207
rect 29009 18173 29043 18207
rect 29193 18173 29227 18207
rect 31125 18173 31159 18207
rect 31677 18173 31711 18207
rect 32597 18173 32631 18207
rect 35357 18173 35391 18207
rect 35633 18173 35667 18207
rect 39497 18173 39531 18207
rect 54309 18173 54343 18207
rect 20453 18105 20487 18139
rect 24685 18105 24719 18139
rect 28457 18105 28491 18139
rect 38945 18105 38979 18139
rect 40325 18105 40359 18139
rect 53205 18105 53239 18139
rect 26985 18037 27019 18071
rect 31769 18037 31803 18071
rect 41337 18037 41371 18071
rect 41797 18037 41831 18071
rect 50537 18037 50571 18071
rect 52745 18037 52779 18071
rect 53389 18037 53423 18071
rect 56057 18037 56091 18071
rect 57437 18037 57471 18071
rect 24685 17833 24719 17867
rect 25789 17833 25823 17867
rect 25973 17833 26007 17867
rect 35173 17833 35207 17867
rect 36001 17833 36035 17867
rect 38393 17833 38427 17867
rect 38669 17833 38703 17867
rect 39957 17833 39991 17867
rect 40693 17833 40727 17867
rect 43729 17833 43763 17867
rect 43821 17833 43855 17867
rect 49065 17833 49099 17867
rect 49525 17833 49559 17867
rect 49893 17833 49927 17867
rect 58265 17833 58299 17867
rect 36461 17765 36495 17799
rect 36645 17765 36679 17799
rect 54953 17765 54987 17799
rect 56057 17765 56091 17799
rect 30757 17697 30791 17731
rect 40049 17697 40083 17731
rect 41521 17697 41555 17731
rect 42993 17697 43027 17731
rect 46489 17697 46523 17731
rect 48237 17697 48271 17731
rect 49525 17697 49559 17731
rect 50629 17697 50663 17731
rect 52469 17697 52503 17731
rect 54769 17697 54803 17731
rect 56701 17697 56735 17731
rect 16681 17629 16715 17663
rect 26157 17629 26191 17663
rect 26341 17629 26375 17663
rect 26433 17629 26467 17663
rect 30297 17629 30331 17663
rect 34897 17629 34931 17663
rect 34989 17629 35023 17663
rect 35247 17629 35281 17663
rect 36185 17629 36219 17663
rect 36277 17629 36311 17663
rect 36553 17629 36587 17663
rect 36829 17629 36863 17663
rect 36921 17629 36955 17663
rect 37197 17629 37231 17663
rect 40141 17629 40175 17663
rect 40417 17629 40451 17663
rect 40877 17629 40911 17663
rect 40969 17629 41003 17663
rect 41245 17629 41279 17663
rect 43085 17629 43119 17663
rect 43178 17629 43212 17663
rect 43361 17629 43395 17663
rect 43453 17629 43487 17663
rect 43591 17629 43625 17663
rect 48881 17629 48915 17663
rect 49709 17629 49743 17663
rect 54493 17629 54527 17663
rect 54585 17629 54619 17663
rect 54861 17629 54895 17663
rect 55873 17629 55907 17663
rect 56425 17629 56459 17663
rect 56517 17629 56551 17663
rect 56793 17629 56827 17663
rect 56885 17629 56919 17663
rect 57152 17629 57186 17663
rect 31033 17561 31067 17595
rect 37013 17561 37047 17595
rect 39865 17561 39899 17595
rect 40693 17561 40727 17595
rect 46765 17561 46799 17595
rect 49433 17561 49467 17595
rect 50905 17561 50939 17595
rect 52745 17561 52779 17595
rect 30481 17493 30515 17527
rect 32505 17493 32539 17527
rect 34713 17493 34747 17527
rect 39589 17493 39623 17527
rect 40325 17493 40359 17527
rect 41153 17493 41187 17527
rect 48329 17493 48363 17527
rect 52377 17493 52411 17527
rect 54217 17493 54251 17527
rect 54309 17493 54343 17527
rect 55689 17493 55723 17527
rect 56241 17493 56275 17527
rect 24869 17289 24903 17323
rect 26525 17289 26559 17323
rect 29193 17289 29227 17323
rect 32229 17289 32263 17323
rect 32413 17289 32447 17323
rect 32505 17289 32539 17323
rect 35725 17289 35759 17323
rect 37289 17289 37323 17323
rect 37657 17289 37691 17323
rect 38117 17289 38151 17323
rect 39221 17289 39255 17323
rect 39773 17289 39807 17323
rect 40601 17289 40635 17323
rect 41245 17289 41279 17323
rect 41521 17289 41555 17323
rect 42993 17289 43027 17323
rect 43361 17289 43395 17323
rect 47593 17289 47627 17323
rect 49525 17289 49559 17323
rect 49709 17289 49743 17323
rect 50445 17289 50479 17323
rect 50629 17289 50663 17323
rect 53297 17289 53331 17323
rect 54033 17289 54067 17323
rect 55873 17289 55907 17323
rect 19717 17221 19751 17255
rect 24317 17221 24351 17255
rect 24685 17221 24719 17255
rect 26985 17221 27019 17255
rect 30757 17221 30791 17255
rect 31493 17221 31527 17255
rect 33793 17221 33827 17255
rect 40233 17221 40267 17255
rect 41153 17221 41187 17255
rect 42625 17221 42659 17255
rect 42717 17221 42751 17255
rect 48697 17221 48731 17255
rect 49157 17221 49191 17255
rect 49249 17221 49283 17255
rect 50077 17221 50111 17255
rect 53665 17221 53699 17255
rect 54401 17221 54435 17255
rect 56241 17221 56275 17255
rect 19073 17153 19107 17187
rect 19620 17153 19654 17187
rect 19809 17153 19843 17187
rect 19992 17153 20026 17187
rect 20085 17153 20119 17187
rect 23121 17153 23155 17187
rect 24041 17153 24075 17187
rect 24225 17153 24259 17187
rect 24409 17153 24443 17187
rect 25053 17153 25087 17187
rect 25329 17153 25363 17187
rect 25421 17153 25455 17187
rect 25973 17153 26007 17187
rect 26157 17153 26191 17187
rect 27537 17153 27571 17187
rect 29653 17153 29687 17187
rect 29929 17153 29963 17187
rect 30568 17153 30602 17187
rect 30665 17153 30699 17187
rect 30940 17153 30974 17187
rect 31033 17153 31067 17187
rect 31125 17153 31159 17187
rect 31218 17153 31252 17187
rect 31401 17153 31435 17187
rect 31631 17153 31665 17187
rect 33517 17153 33551 17187
rect 35633 17153 35667 17187
rect 35909 17153 35943 17187
rect 36001 17153 36035 17187
rect 36093 17153 36127 17187
rect 36277 17153 36311 17187
rect 38301 17153 38335 17187
rect 38761 17153 38795 17187
rect 38945 17153 38979 17187
rect 39037 17153 39071 17187
rect 39497 17153 39531 17187
rect 39681 17153 39715 17187
rect 39957 17153 39991 17187
rect 40105 17153 40139 17187
rect 40325 17153 40359 17187
rect 40463 17153 40497 17187
rect 40877 17153 40911 17187
rect 42441 17153 42475 17187
rect 42809 17153 42843 17187
rect 46029 17153 46063 17187
rect 46177 17153 46211 17187
rect 46305 17153 46339 17187
rect 46397 17153 46431 17187
rect 46494 17153 46528 17187
rect 47041 17153 47075 17187
rect 47777 17153 47811 17187
rect 47869 17153 47903 17187
rect 48145 17153 48179 17187
rect 48881 17153 48915 17187
rect 49029 17153 49063 17187
rect 49346 17153 49380 17187
rect 49888 17153 49922 17187
rect 49985 17153 50019 17187
rect 50260 17153 50294 17187
rect 50353 17153 50387 17187
rect 50813 17153 50847 17187
rect 50905 17153 50939 17187
rect 51181 17153 51215 17187
rect 51549 17153 51583 17187
rect 52101 17153 52135 17187
rect 52745 17153 52779 17187
rect 52929 17153 52963 17187
rect 53021 17153 53055 17187
rect 53113 17153 53147 17187
rect 53481 17153 53515 17187
rect 53749 17153 53783 17187
rect 53849 17153 53883 17187
rect 17049 17085 17083 17119
rect 17325 17085 17359 17119
rect 18889 17085 18923 17119
rect 19349 17085 19383 17119
rect 23397 17085 23431 17119
rect 25237 17085 25271 17119
rect 25697 17085 25731 17119
rect 26341 17085 26375 17119
rect 27721 17085 27755 17119
rect 27813 17085 27847 17119
rect 29377 17085 29411 17119
rect 35265 17085 35299 17119
rect 37473 17085 37507 17119
rect 43453 17085 43487 17119
rect 43729 17085 43763 17119
rect 45845 17085 45879 17119
rect 46857 17085 46891 17119
rect 47225 17085 47259 17119
rect 48053 17085 48087 17119
rect 54125 17085 54159 17119
rect 55965 17085 55999 17119
rect 57713 17085 57747 17119
rect 18797 17017 18831 17051
rect 19441 17017 19475 17051
rect 25789 17017 25823 17051
rect 30389 17017 30423 17051
rect 35449 17017 35483 17051
rect 36737 17017 36771 17051
rect 40693 17017 40727 17051
rect 43085 17017 43119 17051
rect 19257 16949 19291 16983
rect 22937 16949 22971 16983
rect 23305 16949 23339 16983
rect 24593 16949 24627 16983
rect 25329 16949 25363 16983
rect 25881 16949 25915 16983
rect 27353 16949 27387 16983
rect 29469 16949 29503 16983
rect 29837 16949 29871 16983
rect 30113 16949 30147 16983
rect 31769 16949 31803 16983
rect 31861 16949 31895 16983
rect 36645 16949 36679 16983
rect 38485 16949 38519 16983
rect 45201 16949 45235 16983
rect 45293 16949 45327 16983
rect 46673 16949 46707 16983
rect 48329 16949 48363 16983
rect 48513 16949 48547 16983
rect 51089 16949 51123 16983
rect 22648 16745 22682 16779
rect 24133 16745 24167 16779
rect 25145 16745 25179 16779
rect 25881 16745 25915 16779
rect 26065 16745 26099 16779
rect 28733 16745 28767 16779
rect 30205 16745 30239 16779
rect 37197 16745 37231 16779
rect 38025 16745 38059 16779
rect 39129 16745 39163 16779
rect 43269 16745 43303 16779
rect 43637 16745 43671 16779
rect 44281 16745 44315 16779
rect 45937 16745 45971 16779
rect 48329 16745 48363 16779
rect 48421 16745 48455 16779
rect 56885 16745 56919 16779
rect 19257 16677 19291 16711
rect 26341 16677 26375 16711
rect 37565 16677 37599 16711
rect 38485 16677 38519 16711
rect 39681 16677 39715 16711
rect 49985 16677 50019 16711
rect 16681 16609 16715 16643
rect 16957 16609 16991 16643
rect 18521 16609 18555 16643
rect 20545 16609 20579 16643
rect 22385 16609 22419 16643
rect 26985 16609 27019 16643
rect 27261 16609 27295 16643
rect 30665 16609 30699 16643
rect 31309 16609 31343 16643
rect 33057 16609 33091 16643
rect 35357 16609 35391 16643
rect 40969 16609 41003 16643
rect 45661 16609 45695 16643
rect 47409 16609 47443 16643
rect 18705 16541 18739 16575
rect 18889 16541 18923 16575
rect 18981 16541 19015 16575
rect 19436 16541 19470 16575
rect 19808 16541 19842 16575
rect 19901 16541 19935 16575
rect 24409 16541 24443 16575
rect 24502 16541 24536 16575
rect 24685 16541 24719 16575
rect 24915 16541 24949 16575
rect 25329 16541 25363 16575
rect 25605 16541 25639 16575
rect 25697 16541 25731 16575
rect 26157 16541 26191 16575
rect 26525 16541 26559 16575
rect 26617 16541 26651 16575
rect 26801 16541 26835 16575
rect 26893 16541 26927 16575
rect 29009 16541 29043 16575
rect 29193 16541 29227 16575
rect 29377 16541 29411 16575
rect 29561 16541 29595 16575
rect 29654 16541 29688 16575
rect 29837 16541 29871 16575
rect 30067 16541 30101 16575
rect 35081 16541 35115 16575
rect 35173 16541 35207 16575
rect 35449 16541 35483 16575
rect 35725 16541 35759 16575
rect 35909 16541 35943 16575
rect 36093 16541 36127 16575
rect 36737 16541 36771 16575
rect 37749 16541 37783 16575
rect 38577 16541 38611 16575
rect 38945 16541 38979 16575
rect 39313 16541 39347 16575
rect 40049 16541 40083 16575
rect 40417 16541 40451 16575
rect 40693 16541 40727 16575
rect 40785 16541 40819 16575
rect 41061 16541 41095 16575
rect 41429 16541 41463 16575
rect 41981 16541 42015 16575
rect 42809 16541 42843 16575
rect 42993 16541 43027 16575
rect 43085 16541 43119 16575
rect 43315 16541 43349 16575
rect 44005 16541 44039 16575
rect 44097 16541 44131 16575
rect 44373 16541 44407 16575
rect 46397 16541 46431 16575
rect 47685 16541 47719 16575
rect 47778 16541 47812 16575
rect 48169 16541 48203 16575
rect 48605 16541 48639 16575
rect 48973 16541 49007 16575
rect 49433 16541 49467 16575
rect 49617 16541 49651 16575
rect 49801 16541 49835 16575
rect 56057 16541 56091 16575
rect 56333 16541 56367 16575
rect 56701 16541 56735 16575
rect 57161 16541 57195 16575
rect 57529 16541 57563 16575
rect 19533 16473 19567 16507
rect 19625 16473 19659 16507
rect 20821 16473 20855 16507
rect 24777 16473 24811 16507
rect 25513 16473 25547 16507
rect 29101 16473 29135 16507
rect 29929 16473 29963 16507
rect 32781 16473 32815 16507
rect 35817 16473 35851 16507
rect 36553 16473 36587 16507
rect 37289 16473 37323 16507
rect 37933 16473 37967 16507
rect 38301 16473 38335 16507
rect 38761 16473 38795 16507
rect 38853 16473 38887 16507
rect 40141 16473 40175 16507
rect 40233 16473 40267 16507
rect 43545 16473 43579 16507
rect 46581 16473 46615 16507
rect 47961 16473 47995 16507
rect 48053 16473 48087 16507
rect 48697 16473 48731 16507
rect 48789 16473 48823 16507
rect 49065 16473 49099 16507
rect 49525 16473 49559 16507
rect 54217 16473 54251 16507
rect 55321 16473 55355 16507
rect 56517 16473 56551 16507
rect 56609 16473 56643 16507
rect 57253 16473 57287 16507
rect 57345 16473 57379 16507
rect 18429 16405 18463 16439
rect 22293 16405 22327 16439
rect 25053 16405 25087 16439
rect 28825 16405 28859 16439
rect 30297 16405 30331 16439
rect 31217 16405 31251 16439
rect 34897 16405 34931 16439
rect 35541 16405 35575 16439
rect 36461 16405 36495 16439
rect 36921 16405 36955 16439
rect 39405 16405 39439 16439
rect 39865 16405 39899 16439
rect 40509 16405 40543 16439
rect 41153 16405 41187 16439
rect 42625 16405 42659 16439
rect 43821 16405 43855 16439
rect 49249 16405 49283 16439
rect 56977 16405 57011 16439
rect 19901 16201 19935 16235
rect 21189 16201 21223 16235
rect 23121 16201 23155 16235
rect 24961 16201 24995 16235
rect 25329 16201 25363 16235
rect 27905 16201 27939 16235
rect 29193 16201 29227 16235
rect 31125 16201 31159 16235
rect 31677 16201 31711 16235
rect 36461 16201 36495 16235
rect 39865 16201 39899 16235
rect 44465 16201 44499 16235
rect 47409 16201 47443 16235
rect 49341 16201 49375 16235
rect 49709 16201 49743 16235
rect 49801 16201 49835 16235
rect 50445 16201 50479 16235
rect 53297 16201 53331 16235
rect 22109 16133 22143 16167
rect 23397 16133 23431 16167
rect 24685 16133 24719 16167
rect 27353 16133 27387 16167
rect 27445 16133 27479 16167
rect 29653 16133 29687 16167
rect 33241 16133 33275 16167
rect 36737 16133 36771 16167
rect 39497 16133 39531 16167
rect 40325 16133 40359 16167
rect 42901 16133 42935 16167
rect 50169 16133 50203 16167
rect 52837 16133 52871 16167
rect 55229 16133 55263 16167
rect 55321 16133 55355 16167
rect 19257 16065 19291 16099
rect 19405 16065 19439 16099
rect 19533 16065 19567 16099
rect 19625 16065 19659 16099
rect 19763 16065 19797 16099
rect 21373 16065 21407 16099
rect 22012 16065 22046 16099
rect 22201 16065 22235 16099
rect 22329 16065 22363 16099
rect 22477 16065 22511 16099
rect 23300 16065 23334 16099
rect 23489 16065 23523 16099
rect 23672 16065 23706 16099
rect 23765 16065 23799 16099
rect 24409 16065 24443 16099
rect 24593 16065 24627 16099
rect 24777 16065 24811 16099
rect 25237 16065 25271 16099
rect 26249 16065 26283 16099
rect 26433 16065 26467 16099
rect 26525 16065 26559 16099
rect 26617 16065 26651 16099
rect 27077 16065 27111 16099
rect 27170 16065 27204 16099
rect 27542 16065 27576 16099
rect 28089 16065 28123 16099
rect 29377 16065 29411 16099
rect 31217 16065 31251 16099
rect 31493 16065 31527 16099
rect 32413 16065 32447 16099
rect 33609 16065 33643 16099
rect 35909 16065 35943 16099
rect 36001 16065 36035 16099
rect 36277 16065 36311 16099
rect 36645 16065 36679 16099
rect 36829 16065 36863 16099
rect 37013 16065 37047 16099
rect 37933 16065 37967 16099
rect 38301 16065 38335 16099
rect 38393 16065 38427 16099
rect 38485 16065 38519 16099
rect 38669 16065 38703 16099
rect 39129 16065 39163 16099
rect 39313 16065 39347 16099
rect 39589 16065 39623 16099
rect 39681 16065 39715 16099
rect 40049 16065 40083 16099
rect 44649 16065 44683 16099
rect 44741 16065 44775 16099
rect 44833 16065 44867 16099
rect 45017 16065 45051 16099
rect 46581 16065 46615 16099
rect 48145 16065 48179 16099
rect 48329 16065 48363 16099
rect 48422 16065 48456 16099
rect 48605 16065 48639 16099
rect 48697 16065 48731 16099
rect 48794 16065 48828 16099
rect 49065 16065 49099 16099
rect 49433 16065 49467 16099
rect 49985 16065 50019 16099
rect 50077 16065 50111 16099
rect 50353 16065 50387 16099
rect 54309 16065 54343 16099
rect 54585 16065 54619 16099
rect 54769 16065 54803 16099
rect 55045 16065 55079 16099
rect 55505 16065 55539 16099
rect 21649 15997 21683 16031
rect 28181 15997 28215 16031
rect 33885 15997 33919 16031
rect 35357 15997 35391 16031
rect 37381 15997 37415 16031
rect 42625 15997 42659 16031
rect 44373 15997 44407 16031
rect 46765 15997 46799 16031
rect 46857 15997 46891 16031
rect 47593 15997 47627 16031
rect 55965 15997 55999 16031
rect 56241 15997 56275 16031
rect 21557 15929 21591 15963
rect 21833 15929 21867 15963
rect 26801 15929 26835 15963
rect 32229 15929 32263 15963
rect 48973 15929 49007 15963
rect 54493 15929 54527 15963
rect 25513 15861 25547 15895
rect 27721 15861 27755 15895
rect 31309 15861 31343 15895
rect 35725 15861 35759 15895
rect 36185 15861 36219 15895
rect 37841 15861 37875 15895
rect 38117 15861 38151 15895
rect 38853 15861 38887 15895
rect 41797 15861 41831 15895
rect 46397 15861 46431 15895
rect 53113 15861 53147 15895
rect 57713 15861 57747 15895
rect 13277 15657 13311 15691
rect 19625 15657 19659 15691
rect 19901 15657 19935 15691
rect 24869 15657 24903 15691
rect 27077 15657 27111 15691
rect 36645 15657 36679 15691
rect 39037 15657 39071 15691
rect 39405 15657 39439 15691
rect 40509 15657 40543 15691
rect 42993 15657 43027 15691
rect 48145 15657 48179 15691
rect 48973 15657 49007 15691
rect 55873 15657 55907 15691
rect 56609 15657 56643 15691
rect 25513 15589 25547 15623
rect 26985 15589 27019 15623
rect 30573 15589 30607 15623
rect 31033 15589 31067 15623
rect 48053 15589 48087 15623
rect 51917 15589 51951 15623
rect 52469 15589 52503 15623
rect 53389 15589 53423 15623
rect 12449 15521 12483 15555
rect 12909 15521 12943 15555
rect 19717 15521 19751 15555
rect 22477 15521 22511 15555
rect 25421 15521 25455 15555
rect 31125 15521 31159 15555
rect 31585 15521 31619 15555
rect 32137 15521 32171 15555
rect 34897 15521 34931 15555
rect 35173 15521 35207 15555
rect 40877 15521 40911 15555
rect 45661 15521 45695 15555
rect 50721 15521 50755 15555
rect 53941 15521 53975 15555
rect 55045 15521 55079 15555
rect 56057 15521 56091 15555
rect 57069 15521 57103 15555
rect 12541 15453 12575 15487
rect 14105 15453 14139 15487
rect 14749 15453 14783 15487
rect 19441 15453 19475 15487
rect 19809 15453 19843 15487
rect 20085 15453 20119 15487
rect 22201 15453 22235 15487
rect 22385 15453 22419 15487
rect 22937 15453 22971 15487
rect 23121 15453 23155 15487
rect 23213 15453 23247 15487
rect 24685 15453 24719 15487
rect 25697 15453 25731 15487
rect 29929 15453 29963 15487
rect 30077 15453 30111 15487
rect 30297 15453 30331 15487
rect 30435 15453 30469 15487
rect 30849 15453 30883 15487
rect 33057 15453 33091 15487
rect 37289 15453 37323 15487
rect 39957 15453 39991 15487
rect 40141 15453 40175 15487
rect 40233 15453 40267 15487
rect 40325 15453 40359 15487
rect 42441 15453 42475 15487
rect 42809 15453 42843 15487
rect 43545 15453 43579 15487
rect 43729 15453 43763 15487
rect 43913 15453 43947 15487
rect 48697 15453 48731 15487
rect 48789 15453 48823 15487
rect 49065 15453 49099 15487
rect 50169 15453 50203 15487
rect 51365 15453 51399 15487
rect 51549 15453 51583 15487
rect 51733 15453 51767 15487
rect 52193 15453 52227 15487
rect 52285 15453 52319 15487
rect 52561 15453 52595 15487
rect 52837 15453 52871 15487
rect 53113 15453 53147 15487
rect 53205 15453 53239 15487
rect 53665 15453 53699 15487
rect 53757 15453 53791 15487
rect 54033 15453 54067 15487
rect 54401 15453 54435 15487
rect 55321 15453 55355 15487
rect 55597 15453 55631 15487
rect 55689 15453 55723 15487
rect 55965 15453 55999 15487
rect 56241 15453 56275 15487
rect 56333 15453 56367 15487
rect 56793 15453 56827 15487
rect 56885 15453 56919 15487
rect 57161 15453 57195 15487
rect 13461 15385 13495 15419
rect 23305 15385 23339 15419
rect 24133 15385 24167 15419
rect 30205 15385 30239 15419
rect 31309 15385 31343 15419
rect 36829 15385 36863 15419
rect 37565 15385 37599 15419
rect 39497 15385 39531 15419
rect 42625 15385 42659 15419
rect 42717 15385 42751 15419
rect 43821 15385 43855 15419
rect 45937 15385 45971 15419
rect 51641 15385 51675 15419
rect 53021 15385 53055 15419
rect 53481 15385 53515 15419
rect 55505 15385 55539 15419
rect 13093 15317 13127 15351
rect 13261 15317 13295 15351
rect 19257 15317 19291 15351
rect 20269 15317 20303 15351
rect 22017 15317 22051 15351
rect 22753 15317 22787 15351
rect 24501 15317 24535 15351
rect 25881 15317 25915 15351
rect 30665 15317 30699 15351
rect 37105 15317 37139 15351
rect 40693 15317 40727 15351
rect 44097 15317 44131 15351
rect 47409 15317 47443 15351
rect 48513 15317 48547 15351
rect 52009 15317 52043 15351
rect 52745 15317 52779 15351
rect 56517 15317 56551 15351
rect 19625 15113 19659 15147
rect 19717 15113 19751 15147
rect 22201 15113 22235 15147
rect 23213 15113 23247 15147
rect 25605 15113 25639 15147
rect 26341 15113 26375 15147
rect 31953 15113 31987 15147
rect 37749 15113 37783 15147
rect 38485 15113 38519 15147
rect 39497 15113 39531 15147
rect 39681 15113 39715 15147
rect 46489 15113 46523 15147
rect 49893 15113 49927 15147
rect 49985 15113 50019 15147
rect 51641 15113 51675 15147
rect 52285 15113 52319 15147
rect 13277 15045 13311 15079
rect 18153 15045 18187 15079
rect 19993 15045 20027 15079
rect 25881 15045 25915 15079
rect 25973 15045 26007 15079
rect 30481 15045 30515 15079
rect 33425 15045 33459 15079
rect 33609 15045 33643 15079
rect 46857 15045 46891 15079
rect 52009 15045 52043 15079
rect 52377 15045 52411 15079
rect 52745 15045 52779 15079
rect 53297 15045 53331 15079
rect 56425 15045 56459 15079
rect 12633 14977 12667 15011
rect 12725 14977 12759 15011
rect 12909 14977 12943 15011
rect 13001 14977 13035 15011
rect 15117 14977 15151 15011
rect 15393 14977 15427 15011
rect 19855 14977 19889 15011
rect 20085 14977 20119 15011
rect 20268 14977 20302 15011
rect 20361 14977 20395 15011
rect 20545 14977 20579 15011
rect 20913 14977 20947 15011
rect 22380 14977 22414 15011
rect 22477 14977 22511 15011
rect 22569 14977 22603 15011
rect 22752 14977 22786 15011
rect 22845 14977 22879 15011
rect 23029 14977 23063 15011
rect 23581 14977 23615 15011
rect 25743 14977 25777 15011
rect 26156 14977 26190 15011
rect 26249 14977 26283 15011
rect 33241 14977 33275 15011
rect 36645 14977 36679 15011
rect 37933 14977 37967 15011
rect 38025 14977 38059 15011
rect 38301 14977 38335 15011
rect 38669 14977 38703 15011
rect 39221 14977 39255 15011
rect 42717 14977 42751 15011
rect 42809 14977 42843 15011
rect 43085 14977 43119 15011
rect 44925 14977 44959 15011
rect 46668 14977 46702 15011
rect 46765 14977 46799 15011
rect 47040 14977 47074 15011
rect 47133 14977 47167 15011
rect 48145 14977 48179 15011
rect 51825 14977 51859 15011
rect 56701 14977 56735 15011
rect 15301 14909 15335 14943
rect 17877 14909 17911 14943
rect 30205 14909 30239 14943
rect 44649 14909 44683 14943
rect 53021 14909 53055 14943
rect 54769 14909 54803 14943
rect 54953 14909 54987 14943
rect 34621 14841 34655 14875
rect 43177 14841 43211 14875
rect 12909 14773 12943 14807
rect 14749 14773 14783 14807
rect 15117 14773 15151 14807
rect 15577 14773 15611 14807
rect 36553 14773 36587 14807
rect 38209 14773 38243 14807
rect 42533 14773 42567 14807
rect 42993 14773 43027 14807
rect 47225 14773 47259 14807
rect 48408 14773 48442 14807
rect 13277 14569 13311 14603
rect 19257 14569 19291 14603
rect 23305 14569 23339 14603
rect 24501 14569 24535 14603
rect 24777 14569 24811 14603
rect 26709 14569 26743 14603
rect 34345 14569 34379 14603
rect 34759 14569 34793 14603
rect 37105 14569 37139 14603
rect 43729 14569 43763 14603
rect 47317 14569 47351 14603
rect 48421 14569 48455 14603
rect 36829 14501 36863 14535
rect 12725 14433 12759 14467
rect 13001 14433 13035 14467
rect 13829 14433 13863 14467
rect 14749 14433 14783 14467
rect 15117 14433 15151 14467
rect 15393 14433 15427 14467
rect 16957 14433 16991 14467
rect 17233 14433 17267 14467
rect 20729 14433 20763 14467
rect 21741 14433 21775 14467
rect 26249 14433 26283 14467
rect 26525 14433 26559 14467
rect 27353 14433 27387 14467
rect 29377 14433 29411 14467
rect 32597 14433 32631 14467
rect 36553 14433 36587 14467
rect 40601 14433 40635 14467
rect 42533 14433 42567 14467
rect 43637 14433 43671 14467
rect 51457 14433 51491 14467
rect 1409 14365 1443 14399
rect 1685 14365 1719 14399
rect 12173 14365 12207 14399
rect 12357 14365 12391 14399
rect 12633 14365 12667 14399
rect 15025 14365 15059 14399
rect 21005 14365 21039 14399
rect 21465 14365 21499 14399
rect 23443 14365 23477 14399
rect 23581 14365 23615 14399
rect 23856 14365 23890 14399
rect 23949 14365 23983 14399
rect 24685 14365 24719 14399
rect 26893 14365 26927 14399
rect 27169 14365 27203 14399
rect 29745 14365 29779 14399
rect 29837 14365 29871 14399
rect 29929 14365 29963 14399
rect 30021 14365 30055 14399
rect 30757 14365 30791 14399
rect 30941 14365 30975 14399
rect 31033 14365 31067 14399
rect 36185 14365 36219 14399
rect 36645 14365 36679 14399
rect 37013 14365 37047 14399
rect 37197 14365 37231 14399
rect 40785 14365 40819 14399
rect 40969 14365 41003 14399
rect 41061 14365 41095 14399
rect 41153 14365 41187 14399
rect 41521 14365 41555 14399
rect 42257 14365 42291 14399
rect 42349 14365 42383 14399
rect 42625 14365 42659 14399
rect 43361 14365 43395 14399
rect 43913 14365 43947 14399
rect 44281 14365 44315 14399
rect 46581 14365 46615 14399
rect 46765 14365 46799 14399
rect 46857 14365 46891 14399
rect 48605 14365 48639 14399
rect 48789 14365 48823 14399
rect 48973 14365 49007 14399
rect 49249 14365 49283 14399
rect 49341 14365 49375 14399
rect 49433 14365 49467 14399
rect 49617 14365 49651 14399
rect 49985 14365 50019 14399
rect 50261 14365 50295 14399
rect 50537 14365 50571 14399
rect 50629 14365 50663 14399
rect 14105 14297 14139 14331
rect 18521 14297 18555 14331
rect 18889 14297 18923 14331
rect 23673 14297 23707 14331
rect 26985 14297 27019 14331
rect 29101 14297 29135 14331
rect 30297 14297 30331 14331
rect 32873 14297 32907 14331
rect 44005 14297 44039 14331
rect 44097 14297 44131 14331
rect 47041 14297 47075 14331
rect 47225 14297 47259 14331
rect 48697 14297 48731 14331
rect 50445 14297 50479 14331
rect 51733 14297 51767 14331
rect 1593 14229 1627 14263
rect 12265 14229 12299 14263
rect 15485 14229 15519 14263
rect 18705 14229 18739 14263
rect 18981 14229 19015 14263
rect 23213 14229 23247 14263
rect 24225 14229 24259 14263
rect 27629 14229 27663 14263
rect 29561 14229 29595 14263
rect 30389 14229 30423 14263
rect 40049 14229 40083 14263
rect 41337 14229 41371 14263
rect 42073 14229 42107 14263
rect 46397 14229 46431 14263
rect 47593 14229 47627 14263
rect 47777 14229 47811 14263
rect 49065 14229 49099 14263
rect 49801 14229 49835 14263
rect 50813 14229 50847 14263
rect 53205 14229 53239 14263
rect 15301 14025 15335 14059
rect 18337 14025 18371 14059
rect 18981 14025 19015 14059
rect 33057 14025 33091 14059
rect 33425 14025 33459 14059
rect 34437 14025 34471 14059
rect 35725 14025 35759 14059
rect 44189 14025 44223 14059
rect 44281 14025 44315 14059
rect 46121 14025 46155 14059
rect 46305 14025 46339 14059
rect 47133 14025 47167 14059
rect 47593 14025 47627 14059
rect 53113 14025 53147 14059
rect 13185 13957 13219 13991
rect 19349 13957 19383 13991
rect 22109 13957 22143 13991
rect 25329 13957 25363 13991
rect 32781 13957 32815 13991
rect 34253 13957 34287 13991
rect 36001 13957 36035 13991
rect 36093 13957 36127 13991
rect 41981 13957 42015 13991
rect 42717 13957 42751 13991
rect 46673 13957 46707 13991
rect 50721 13957 50755 13991
rect 52193 13957 52227 13991
rect 52837 13957 52871 13991
rect 53297 13957 53331 13991
rect 15853 13889 15887 13923
rect 18153 13889 18187 13923
rect 18429 13889 18463 13923
rect 18613 13889 18647 13923
rect 18797 13889 18831 13923
rect 19165 13889 19199 13923
rect 19625 13889 19659 13923
rect 20269 13889 20303 13923
rect 21833 13889 21867 13923
rect 23857 13889 23891 13923
rect 24225 13889 24259 13923
rect 24317 13889 24351 13923
rect 24410 13889 24444 13923
rect 24593 13889 24627 13923
rect 24685 13889 24719 13923
rect 24823 13889 24857 13923
rect 25053 13889 25087 13923
rect 28641 13889 28675 13923
rect 32137 13889 32171 13923
rect 32597 13889 32631 13923
rect 32965 13889 32999 13923
rect 33885 13889 33919 13923
rect 35909 13889 35943 13923
rect 36277 13889 36311 13923
rect 36645 13889 36679 13923
rect 36737 13889 36771 13923
rect 36921 13889 36955 13923
rect 37013 13889 37047 13923
rect 38669 13889 38703 13923
rect 42257 13889 42291 13923
rect 42441 13889 42475 13923
rect 44465 13889 44499 13923
rect 44557 13889 44591 13923
rect 44833 13889 44867 13923
rect 45937 13889 45971 13923
rect 46484 13889 46518 13923
rect 46581 13889 46615 13923
rect 46856 13889 46890 13923
rect 46949 13889 46983 13923
rect 47317 13889 47351 13923
rect 48237 13889 48271 13923
rect 49065 13889 49099 13923
rect 49157 13889 49191 13923
rect 49433 13889 49467 13923
rect 49801 13889 49835 13923
rect 51273 13889 51307 13923
rect 51641 13889 51675 13923
rect 51733 13889 51767 13923
rect 52009 13889 52043 13923
rect 58265 13889 58299 13923
rect 12909 13821 12943 13855
rect 14657 13821 14691 13855
rect 19901 13821 19935 13855
rect 20085 13821 20119 13855
rect 26801 13821 26835 13855
rect 28917 13821 28951 13855
rect 31033 13821 31067 13855
rect 32229 13821 32263 13855
rect 33517 13821 33551 13855
rect 33701 13821 33735 13855
rect 38945 13821 38979 13855
rect 40417 13821 40451 13855
rect 40509 13821 40543 13855
rect 44741 13821 44775 13855
rect 48421 13821 48455 13855
rect 23581 13753 23615 13787
rect 30389 13753 30423 13787
rect 34069 13753 34103 13787
rect 34621 13753 34655 13787
rect 19533 13685 19567 13719
rect 24961 13685 24995 13719
rect 30481 13685 30515 13719
rect 36461 13685 36495 13719
rect 48697 13685 48731 13719
rect 48881 13685 48915 13719
rect 49341 13685 49375 13719
rect 51457 13685 51491 13719
rect 51917 13685 51951 13719
rect 52285 13685 52319 13719
rect 53481 13685 53515 13719
rect 58449 13685 58483 13719
rect 13737 13481 13771 13515
rect 15301 13481 15335 13515
rect 24041 13481 24075 13515
rect 24685 13481 24719 13515
rect 29561 13481 29595 13515
rect 33057 13481 33091 13515
rect 36001 13481 36035 13515
rect 36277 13481 36311 13515
rect 36461 13481 36495 13515
rect 37657 13481 37691 13515
rect 37749 13481 37783 13515
rect 39037 13481 39071 13515
rect 41061 13481 41095 13515
rect 42165 13481 42199 13515
rect 45845 13481 45879 13515
rect 48513 13481 48547 13515
rect 48789 13481 48823 13515
rect 51917 13481 51951 13515
rect 52009 13481 52043 13515
rect 54861 13481 54895 13515
rect 54953 13481 54987 13515
rect 37933 13413 37967 13447
rect 54585 13413 54619 13447
rect 55321 13413 55355 13447
rect 12265 13345 12299 13379
rect 16405 13345 16439 13379
rect 16681 13345 16715 13379
rect 17325 13345 17359 13379
rect 20085 13345 20119 13379
rect 23673 13345 23707 13379
rect 26617 13345 26651 13379
rect 30021 13345 30055 13379
rect 35909 13345 35943 13379
rect 37013 13345 37047 13379
rect 37105 13345 37139 13379
rect 37565 13345 37599 13379
rect 39681 13345 39715 13379
rect 40785 13345 40819 13379
rect 46029 13345 46063 13379
rect 46305 13345 46339 13379
rect 47777 13345 47811 13379
rect 49801 13345 49835 13379
rect 50169 13345 50203 13379
rect 50445 13345 50479 13379
rect 55505 13345 55539 13379
rect 55781 13345 55815 13379
rect 11989 13277 12023 13311
rect 14933 13277 14967 13311
rect 15025 13277 15059 13311
rect 15393 13277 15427 13311
rect 16773 13277 16807 13311
rect 17049 13277 17083 13311
rect 17233 13277 17267 13311
rect 19809 13277 19843 13311
rect 20361 13277 20395 13311
rect 24133 13277 24167 13311
rect 24869 13277 24903 13311
rect 26893 13277 26927 13311
rect 29745 13277 29779 13311
rect 29837 13277 29871 13311
rect 30113 13277 30147 13311
rect 30849 13277 30883 13311
rect 31125 13277 31159 13311
rect 32137 13277 32171 13311
rect 32321 13277 32355 13311
rect 32413 13277 32447 13311
rect 36093 13277 36127 13311
rect 36185 13277 36219 13311
rect 36461 13277 36495 13311
rect 36553 13277 36587 13311
rect 37289 13277 37323 13311
rect 39162 13277 39196 13311
rect 39589 13277 39623 13311
rect 40049 13277 40083 13311
rect 45569 13277 45603 13311
rect 45661 13277 45695 13311
rect 45937 13277 45971 13311
rect 48053 13277 48087 13311
rect 48145 13277 48179 13311
rect 48237 13277 48271 13311
rect 48421 13277 48455 13311
rect 48973 13277 49007 13311
rect 54677 13277 54711 13311
rect 54861 13277 54895 13311
rect 14749 13209 14783 13243
rect 16221 13209 16255 13243
rect 17601 13209 17635 13243
rect 24501 13209 24535 13243
rect 30665 13209 30699 13243
rect 36921 13209 36955 13243
rect 37473 13209 37507 13243
rect 37933 13209 37967 13243
rect 42073 13209 42107 13243
rect 49065 13209 49099 13243
rect 15117 13141 15151 13175
rect 17141 13141 17175 13175
rect 19073 13141 19107 13175
rect 19257 13141 19291 13175
rect 25513 13141 25547 13175
rect 31033 13141 31067 13175
rect 31953 13141 31987 13175
rect 39221 13141 39255 13175
rect 45385 13141 45419 13175
rect 47869 13141 47903 13175
rect 57253 13141 57287 13175
rect 16497 12937 16531 12971
rect 16865 12937 16899 12971
rect 17601 12937 17635 12971
rect 23765 12937 23799 12971
rect 25605 12937 25639 12971
rect 26525 12937 26559 12971
rect 27629 12937 27663 12971
rect 32137 12937 32171 12971
rect 32505 12937 32539 12971
rect 33333 12937 33367 12971
rect 33517 12937 33551 12971
rect 36645 12937 36679 12971
rect 37289 12937 37323 12971
rect 38577 12937 38611 12971
rect 39313 12937 39347 12971
rect 50537 12937 50571 12971
rect 57621 12937 57655 12971
rect 18429 12869 18463 12903
rect 18613 12869 18647 12903
rect 26709 12869 26743 12903
rect 39129 12869 39163 12903
rect 45477 12869 45511 12903
rect 49065 12869 49099 12903
rect 16037 12801 16071 12835
rect 17509 12801 17543 12835
rect 18337 12801 18371 12835
rect 19625 12801 19659 12835
rect 19809 12801 19843 12835
rect 25513 12801 25547 12835
rect 25789 12801 25823 12835
rect 25973 12801 26007 12835
rect 26341 12801 26375 12835
rect 26617 12801 26651 12835
rect 27721 12801 27755 12835
rect 28549 12801 28583 12835
rect 28733 12801 28767 12835
rect 29009 12801 29043 12835
rect 29469 12801 29503 12835
rect 29653 12801 29687 12835
rect 32321 12801 32355 12835
rect 32597 12801 32631 12835
rect 33336 12801 33370 12835
rect 36553 12801 36587 12835
rect 36829 12801 36863 12835
rect 37013 12801 37047 12835
rect 37473 12801 37507 12835
rect 37657 12801 37691 12835
rect 38485 12801 38519 12835
rect 38761 12801 38795 12835
rect 38853 12801 38887 12835
rect 39037 12801 39071 12835
rect 39221 12801 39255 12835
rect 39405 12801 39439 12835
rect 39497 12801 39531 12835
rect 42809 12801 42843 12835
rect 43637 12801 43671 12835
rect 45201 12801 45235 12835
rect 48789 12801 48823 12835
rect 57437 12801 57471 12835
rect 18245 12733 18279 12767
rect 21097 12733 21131 12767
rect 25237 12733 25271 12767
rect 26065 12733 26099 12767
rect 27905 12733 27939 12767
rect 28825 12733 28859 12767
rect 32873 12733 32907 12767
rect 38669 12733 38703 12767
rect 42901 12733 42935 12767
rect 42993 12733 43027 12767
rect 44281 12733 44315 12767
rect 18613 12665 18647 12699
rect 26157 12665 26191 12699
rect 28917 12665 28951 12699
rect 19625 12597 19659 12631
rect 20453 12597 20487 12631
rect 27261 12597 27295 12631
rect 29653 12597 29687 12631
rect 32965 12597 32999 12631
rect 42441 12597 42475 12631
rect 46949 12597 46983 12631
rect 17233 12393 17267 12427
rect 18337 12393 18371 12427
rect 19533 12393 19567 12427
rect 26617 12393 26651 12427
rect 27997 12393 28031 12427
rect 29561 12393 29595 12427
rect 30297 12393 30331 12427
rect 30481 12393 30515 12427
rect 31677 12393 31711 12427
rect 33517 12393 33551 12427
rect 43453 12393 43487 12427
rect 46213 12393 46247 12427
rect 46673 12393 46707 12427
rect 13921 12325 13955 12359
rect 17785 12325 17819 12359
rect 26433 12325 26467 12359
rect 26985 12325 27019 12359
rect 28641 12325 28675 12359
rect 12173 12257 12207 12291
rect 14749 12257 14783 12291
rect 15393 12257 15427 12291
rect 15669 12257 15703 12291
rect 17141 12257 17175 12291
rect 18153 12257 18187 12291
rect 19901 12257 19935 12291
rect 20177 12257 20211 12291
rect 22477 12257 22511 12291
rect 22753 12257 22787 12291
rect 24593 12257 24627 12291
rect 24869 12257 24903 12291
rect 29745 12257 29779 12291
rect 32965 12257 32999 12291
rect 34253 12257 34287 12291
rect 41705 12257 41739 12291
rect 14841 12189 14875 12223
rect 15025 12189 15059 12223
rect 17601 12189 17635 12223
rect 18061 12189 18095 12223
rect 18337 12189 18371 12223
rect 18613 12189 18647 12223
rect 18797 12189 18831 12223
rect 19257 12189 19291 12223
rect 19349 12189 19383 12223
rect 19533 12189 19567 12223
rect 19809 12189 19843 12223
rect 20269 12189 20303 12223
rect 20821 12189 20855 12223
rect 27169 12189 27203 12223
rect 27813 12189 27847 12223
rect 27997 12189 28031 12223
rect 28825 12189 28859 12223
rect 28917 12189 28951 12223
rect 29009 12189 29043 12223
rect 29101 12189 29135 12223
rect 29285 12189 29319 12223
rect 29837 12189 29871 12223
rect 30481 12189 30515 12223
rect 30573 12189 30607 12223
rect 31493 12189 31527 12223
rect 31769 12189 31803 12223
rect 33057 12189 33091 12223
rect 33149 12189 33183 12223
rect 33241 12189 33275 12223
rect 33425 12189 33459 12223
rect 33701 12189 33735 12223
rect 33793 12189 33827 12223
rect 33885 12189 33919 12223
rect 33977 12189 34011 12223
rect 34897 12189 34931 12223
rect 34989 12189 35023 12223
rect 35173 12189 35207 12223
rect 35265 12189 35299 12223
rect 35720 12189 35754 12223
rect 35817 12189 35851 12223
rect 36092 12189 36126 12223
rect 36185 12189 36219 12223
rect 38669 12189 38703 12223
rect 39037 12189 39071 12223
rect 39221 12189 39255 12223
rect 39865 12189 39899 12223
rect 39958 12189 39992 12223
rect 40233 12189 40267 12223
rect 40330 12189 40364 12223
rect 40601 12189 40635 12223
rect 40877 12189 40911 12223
rect 40969 12189 41003 12223
rect 46765 12189 46799 12223
rect 12449 12121 12483 12155
rect 14933 12121 14967 12155
rect 17417 12121 17451 12155
rect 26801 12121 26835 12155
rect 30757 12121 30791 12155
rect 35909 12121 35943 12155
rect 40141 12121 40175 12155
rect 40785 12121 40819 12155
rect 41981 12121 42015 12155
rect 14105 12053 14139 12087
rect 17509 12053 17543 12087
rect 17877 12053 17911 12087
rect 18429 12053 18463 12087
rect 21005 12053 21039 12087
rect 26341 12053 26375 12087
rect 26601 12053 26635 12087
rect 27261 12053 27295 12087
rect 30205 12053 30239 12087
rect 31217 12053 31251 12087
rect 32689 12053 32723 12087
rect 35449 12053 35483 12087
rect 35541 12053 35575 12087
rect 38853 12053 38887 12087
rect 39129 12053 39163 12087
rect 40509 12053 40543 12087
rect 41153 12053 41187 12087
rect 29561 11849 29595 11883
rect 32413 11849 32447 11883
rect 33241 11849 33275 11883
rect 33333 11849 33367 11883
rect 34989 11849 35023 11883
rect 35173 11849 35207 11883
rect 36645 11849 36679 11883
rect 37657 11849 37691 11883
rect 38485 11849 38519 11883
rect 39405 11849 39439 11883
rect 39773 11849 39807 11883
rect 44281 11849 44315 11883
rect 19717 11781 19751 11815
rect 29837 11781 29871 11815
rect 29929 11781 29963 11815
rect 31033 11781 31067 11815
rect 31151 11781 31185 11815
rect 32965 11781 32999 11815
rect 33701 11781 33735 11815
rect 36001 11781 36035 11815
rect 36369 11781 36403 11815
rect 40141 11781 40175 11815
rect 42809 11781 42843 11815
rect 12173 11713 12207 11747
rect 14749 11713 14783 11747
rect 14933 11713 14967 11747
rect 19441 11713 19475 11747
rect 26985 11713 27019 11747
rect 27353 11713 27387 11747
rect 28825 11713 28859 11747
rect 29377 11713 29411 11747
rect 29740 11713 29774 11747
rect 30112 11713 30146 11747
rect 30205 11713 30239 11747
rect 30849 11713 30883 11747
rect 30941 11713 30975 11747
rect 32229 11713 32263 11747
rect 32505 11713 32539 11747
rect 32597 11713 32631 11747
rect 32745 11713 32779 11747
rect 32873 11713 32907 11747
rect 33062 11713 33096 11747
rect 33333 11713 33367 11747
rect 33517 11713 33551 11747
rect 33609 11713 33643 11747
rect 33793 11713 33827 11747
rect 35114 11713 35148 11747
rect 35817 11713 35851 11747
rect 36277 11713 36311 11747
rect 36461 11713 36495 11747
rect 36737 11713 36771 11747
rect 37841 11713 37875 11747
rect 38117 11713 38151 11747
rect 38298 11713 38332 11747
rect 38393 11713 38427 11747
rect 38577 11711 38611 11745
rect 38853 11713 38887 11747
rect 38946 11713 38980 11747
rect 39313 11713 39347 11747
rect 39589 11713 39623 11747
rect 39865 11713 39899 11747
rect 39957 11713 39991 11747
rect 42533 11713 42567 11747
rect 12449 11645 12483 11679
rect 13921 11645 13955 11679
rect 14565 11645 14599 11679
rect 21189 11645 21223 11679
rect 22845 11645 22879 11679
rect 29101 11645 29135 11679
rect 29193 11645 29227 11679
rect 31309 11645 31343 11679
rect 35633 11645 35667 11679
rect 36185 11645 36219 11679
rect 38025 11645 38059 11679
rect 38669 11645 38703 11679
rect 39037 11645 39071 11679
rect 39129 11645 39163 11679
rect 27169 11577 27203 11611
rect 32229 11577 32263 11611
rect 35541 11577 35575 11611
rect 37933 11577 37967 11611
rect 40141 11577 40175 11611
rect 14013 11509 14047 11543
rect 15117 11509 15151 11543
rect 22293 11509 22327 11543
rect 27445 11509 27479 11543
rect 29009 11509 29043 11543
rect 29193 11509 29227 11543
rect 30665 11509 30699 11543
rect 12265 11305 12299 11339
rect 15025 11305 15059 11339
rect 16405 11305 16439 11339
rect 16773 11305 16807 11339
rect 22477 11305 22511 11339
rect 27997 11305 28031 11339
rect 28917 11305 28951 11339
rect 30297 11305 30331 11339
rect 38393 11305 38427 11339
rect 38761 11305 38795 11339
rect 39129 11305 39163 11339
rect 39313 11305 39347 11339
rect 14105 11237 14139 11271
rect 15209 11237 15243 11271
rect 15301 11237 15335 11271
rect 16589 11237 16623 11271
rect 18797 11237 18831 11271
rect 32505 11237 32539 11271
rect 35449 11237 35483 11271
rect 40509 11237 40543 11271
rect 12725 11169 12759 11203
rect 14841 11169 14875 11203
rect 16313 11169 16347 11203
rect 21925 11169 21959 11203
rect 22385 11169 22419 11203
rect 23949 11169 23983 11203
rect 28457 11169 28491 11203
rect 32321 11169 32355 11203
rect 39497 11169 39531 11203
rect 40325 11169 40359 11203
rect 12633 11101 12667 11135
rect 14105 11101 14139 11135
rect 14289 11101 14323 11135
rect 14381 11101 14415 11135
rect 15025 11101 15059 11135
rect 15485 11101 15519 11135
rect 16129 11101 16163 11135
rect 16405 11101 16439 11135
rect 16957 11101 16991 11135
rect 17325 11101 17359 11135
rect 18521 11101 18555 11135
rect 19901 11101 19935 11135
rect 20269 11101 20303 11135
rect 20453 11101 20487 11135
rect 22017 11101 22051 11135
rect 24225 11101 24259 11135
rect 27537 11101 27571 11135
rect 28181 11101 28215 11135
rect 28273 11101 28307 11135
rect 28549 11101 28583 11135
rect 29101 11101 29135 11135
rect 30481 11101 30515 11135
rect 30665 11101 30699 11135
rect 30757 11101 30791 11135
rect 32137 11101 32171 11135
rect 32505 11101 32539 11135
rect 34805 11101 34839 11135
rect 34897 11101 34931 11135
rect 35173 11101 35207 11135
rect 35265 11101 35299 11135
rect 38301 11101 38335 11135
rect 38485 11101 38519 11135
rect 38577 11101 38611 11135
rect 39313 11101 39347 11135
rect 39865 11101 39899 11135
rect 40233 11101 40267 11135
rect 14749 11033 14783 11067
rect 15853 11033 15887 11067
rect 17049 11033 17083 11067
rect 18797 11033 18831 11067
rect 19349 11033 19383 11067
rect 27721 11033 27755 11067
rect 27905 11033 27939 11067
rect 35081 11033 35115 11067
rect 39589 11033 39623 11067
rect 15577 10965 15611 10999
rect 15669 10965 15703 10999
rect 17141 10965 17175 10999
rect 18613 10965 18647 10999
rect 20085 10965 20119 10999
rect 13553 10761 13587 10795
rect 16681 10761 16715 10795
rect 20177 10761 20211 10795
rect 26709 10761 26743 10795
rect 27169 10761 27203 10795
rect 27905 10761 27939 10795
rect 28917 10761 28951 10795
rect 29101 10761 29135 10795
rect 29653 10761 29687 10795
rect 31401 10761 31435 10795
rect 32689 10761 32723 10795
rect 32965 10761 32999 10795
rect 35357 10761 35391 10795
rect 37105 10761 37139 10795
rect 37381 10761 37415 10795
rect 37999 10761 38033 10795
rect 39037 10761 39071 10795
rect 13705 10693 13739 10727
rect 13921 10693 13955 10727
rect 16957 10693 16991 10727
rect 18153 10693 18187 10727
rect 18613 10693 18647 10727
rect 21465 10693 21499 10727
rect 28641 10693 28675 10727
rect 30757 10693 30791 10727
rect 30849 10693 30883 10727
rect 35081 10693 35115 10727
rect 37565 10693 37599 10727
rect 37749 10693 37783 10727
rect 38209 10693 38243 10727
rect 39405 10693 39439 10727
rect 13093 10625 13127 10659
rect 14013 10625 14047 10659
rect 14657 10625 14691 10659
rect 16865 10625 16899 10659
rect 17049 10625 17083 10659
rect 18061 10625 18095 10659
rect 18245 10625 18279 10659
rect 20361 10625 20395 10659
rect 20729 10625 20763 10659
rect 21373 10625 21407 10659
rect 21649 10625 21683 10659
rect 27077 10625 27111 10659
rect 27813 10625 27847 10659
rect 27997 10625 28031 10659
rect 28273 10625 28307 10659
rect 28366 10625 28400 10659
rect 28549 10625 28583 10659
rect 28779 10625 28813 10659
rect 29009 10625 29043 10659
rect 29193 10625 29227 10659
rect 29285 10625 29319 10659
rect 29469 10625 29503 10659
rect 31125 10625 31159 10659
rect 32597 10625 32631 10659
rect 32781 10625 32815 10659
rect 32873 10625 32907 10659
rect 33057 10625 33091 10659
rect 34437 10625 34471 10659
rect 35541 10625 35575 10659
rect 35633 10625 35667 10659
rect 35909 10625 35943 10659
rect 36185 10625 36219 10659
rect 36277 10625 36311 10659
rect 36461 10625 36495 10659
rect 36553 10625 36587 10659
rect 38945 10625 38979 10659
rect 39129 10625 39163 10659
rect 39313 10625 39347 10659
rect 39497 10625 39531 10659
rect 13185 10557 13219 10591
rect 18337 10557 18371 10591
rect 20821 10557 20855 10591
rect 23489 10557 23523 10591
rect 23765 10557 23799 10591
rect 24961 10557 24995 10591
rect 25237 10557 25271 10591
rect 31217 10557 31251 10591
rect 34529 10557 34563 10591
rect 17233 10489 17267 10523
rect 22017 10489 22051 10523
rect 34713 10489 34747 10523
rect 13461 10421 13495 10455
rect 13737 10421 13771 10455
rect 20085 10421 20119 10455
rect 20361 10421 20395 10455
rect 21649 10421 21683 10455
rect 27629 10421 27663 10455
rect 29469 10421 29503 10455
rect 35081 10421 35115 10455
rect 35265 10421 35299 10455
rect 35817 10421 35851 10455
rect 36001 10421 36035 10455
rect 37565 10421 37599 10455
rect 37841 10421 37875 10455
rect 38025 10421 38059 10455
rect 14473 10217 14507 10251
rect 18337 10217 18371 10251
rect 22385 10217 22419 10251
rect 22569 10217 22603 10251
rect 22845 10217 22879 10251
rect 25881 10217 25915 10251
rect 27721 10217 27755 10251
rect 29285 10217 29319 10251
rect 29929 10217 29963 10251
rect 31033 10217 31067 10251
rect 31125 10217 31159 10251
rect 32045 10217 32079 10251
rect 38301 10217 38335 10251
rect 13921 10149 13955 10183
rect 14381 10149 14415 10183
rect 19901 10149 19935 10183
rect 22753 10149 22787 10183
rect 36185 10149 36219 10183
rect 36737 10149 36771 10183
rect 12449 10081 12483 10115
rect 16221 10081 16255 10115
rect 16589 10081 16623 10115
rect 22937 10081 22971 10115
rect 26249 10081 26283 10115
rect 27261 10081 27295 10115
rect 30389 10081 30423 10115
rect 30573 10081 30607 10115
rect 32413 10081 32447 10115
rect 32689 10081 32723 10115
rect 32965 10081 32999 10115
rect 33425 10081 33459 10115
rect 35449 10081 35483 10115
rect 35541 10081 35575 10115
rect 35909 10081 35943 10115
rect 39221 10081 39255 10115
rect 41981 10081 42015 10115
rect 12173 10013 12207 10047
rect 14105 10013 14139 10047
rect 14473 10013 14507 10047
rect 14657 10013 14691 10047
rect 16129 10013 16163 10047
rect 18797 10013 18831 10047
rect 20177 10013 20211 10047
rect 20269 10013 20303 10047
rect 22661 10013 22695 10047
rect 23029 10013 23063 10047
rect 23213 10013 23247 10047
rect 26157 10013 26191 10047
rect 27169 10013 27203 10047
rect 27353 10013 27387 10047
rect 27813 10013 27847 10047
rect 30297 10013 30331 10047
rect 30849 10013 30883 10047
rect 31033 10013 31067 10047
rect 31125 10013 31159 10047
rect 31309 10013 31343 10047
rect 32045 10013 32079 10047
rect 32229 10013 32263 10047
rect 32505 10013 32539 10047
rect 32597 10013 32631 10047
rect 33057 10013 33091 10047
rect 33241 10013 33275 10047
rect 35357 10013 35391 10047
rect 36372 10013 36406 10047
rect 36553 10013 36587 10047
rect 36921 10013 36955 10047
rect 37105 10013 37139 10047
rect 37197 10013 37231 10047
rect 37933 10013 37967 10047
rect 38117 10013 38151 10047
rect 39313 10013 39347 10047
rect 40233 10013 40267 10047
rect 14381 9945 14415 9979
rect 16865 9945 16899 9979
rect 18429 9945 18463 9979
rect 20453 9945 20487 9979
rect 22201 9945 22235 9979
rect 28641 9945 28675 9979
rect 28917 9945 28951 9979
rect 29101 9945 29135 9979
rect 36645 9945 36679 9979
rect 40509 9945 40543 9979
rect 14197 9877 14231 9911
rect 16497 9877 16531 9911
rect 20085 9877 20119 9911
rect 22401 9877 22435 9911
rect 23121 9877 23155 9911
rect 32873 9877 32907 9911
rect 39681 9877 39715 9911
rect 14841 9673 14875 9707
rect 16865 9673 16899 9707
rect 29285 9673 29319 9707
rect 30297 9673 30331 9707
rect 40693 9673 40727 9707
rect 13369 9605 13403 9639
rect 33977 9605 34011 9639
rect 34161 9605 34195 9639
rect 36553 9605 36587 9639
rect 16773 9537 16807 9571
rect 16957 9537 16991 9571
rect 21833 9537 21867 9571
rect 21925 9537 21959 9571
rect 22109 9537 22143 9571
rect 22201 9537 22235 9571
rect 28733 9537 28767 9571
rect 29101 9537 29135 9571
rect 29377 9537 29411 9571
rect 30205 9537 30239 9571
rect 30389 9537 30423 9571
rect 32229 9537 32263 9571
rect 32505 9537 32539 9571
rect 32597 9537 32631 9571
rect 32965 9537 32999 9571
rect 33057 9537 33091 9571
rect 33241 9537 33275 9571
rect 33333 9537 33367 9571
rect 33793 9537 33827 9571
rect 36461 9537 36495 9571
rect 36829 9537 36863 9571
rect 37105 9537 37139 9571
rect 37565 9537 37599 9571
rect 41245 9537 41279 9571
rect 13093 9469 13127 9503
rect 22753 9469 22787 9503
rect 23489 9469 23523 9503
rect 33517 9469 33551 9503
rect 36553 9469 36587 9503
rect 22109 9401 22143 9435
rect 33701 9401 33735 9435
rect 22937 9333 22971 9367
rect 32321 9333 32355 9367
rect 32781 9333 32815 9367
rect 33425 9333 33459 9367
rect 33517 9333 33551 9367
rect 36737 9333 36771 9367
rect 37013 9333 37047 9367
rect 37657 9333 37691 9367
rect 21005 9129 21039 9163
rect 21925 9129 21959 9163
rect 22201 9129 22235 9163
rect 27721 9129 27755 9163
rect 28457 9129 28491 9163
rect 28825 9129 28859 9163
rect 32229 9129 32263 9163
rect 33425 9129 33459 9163
rect 22109 9061 22143 9095
rect 28365 9061 28399 9095
rect 23673 8993 23707 9027
rect 28549 8993 28583 9027
rect 36829 8993 36863 9027
rect 39681 8993 39715 9027
rect 17417 8925 17451 8959
rect 21281 8925 21315 8959
rect 23949 8925 23983 8959
rect 27261 8925 27295 8959
rect 27629 8925 27663 8959
rect 27905 8925 27939 8959
rect 27997 8925 28031 8959
rect 32045 8925 32079 8959
rect 32321 8925 32355 8959
rect 32689 8925 32723 8959
rect 37105 8925 37139 8959
rect 37197 8925 37231 8959
rect 37381 8925 37415 8959
rect 20453 8857 20487 8891
rect 21557 8857 21591 8891
rect 21741 8857 21775 8891
rect 21941 8857 21975 8891
rect 39405 8857 39439 8891
rect 18061 8789 18095 8823
rect 20729 8789 20763 8823
rect 21189 8789 21223 8823
rect 21373 8789 21407 8823
rect 27445 8789 27479 8823
rect 32505 8789 32539 8823
rect 35357 8789 35391 8823
rect 37289 8789 37323 8823
rect 37933 8789 37967 8823
rect 21189 8585 21223 8619
rect 23029 8585 23063 8619
rect 29009 8585 29043 8619
rect 31493 8585 31527 8619
rect 32965 8585 32999 8619
rect 37013 8585 37047 8619
rect 37657 8585 37691 8619
rect 38393 8585 38427 8619
rect 36093 8517 36127 8551
rect 36185 8517 36219 8551
rect 15577 8449 15611 8483
rect 15761 8449 15795 8483
rect 15853 8449 15887 8483
rect 16037 8449 16071 8483
rect 18429 8449 18463 8483
rect 19165 8449 19199 8483
rect 21005 8449 21039 8483
rect 21373 8449 21407 8483
rect 21649 8449 21683 8483
rect 22477 8449 22511 8483
rect 31309 8449 31343 8483
rect 31677 8449 31711 8483
rect 31953 8449 31987 8483
rect 35541 8449 35575 8483
rect 35817 8449 35851 8483
rect 36001 8449 36035 8483
rect 36277 8449 36311 8483
rect 36645 8449 36679 8483
rect 36737 8449 36771 8483
rect 37381 8449 37415 8483
rect 37841 8449 37875 8483
rect 38301 8449 38335 8483
rect 40601 8449 40635 8483
rect 16681 8381 16715 8415
rect 18153 8381 18187 8415
rect 19441 8381 19475 8415
rect 20913 8381 20947 8415
rect 22385 8381 22419 8415
rect 22845 8381 22879 8415
rect 24501 8381 24535 8415
rect 24777 8381 24811 8415
rect 25053 8381 25087 8415
rect 25329 8381 25363 8415
rect 26801 8381 26835 8415
rect 27537 8381 27571 8415
rect 28181 8381 28215 8415
rect 28733 8381 28767 8415
rect 32689 8381 32723 8415
rect 38853 8381 38887 8415
rect 40325 8381 40359 8415
rect 32137 8313 32171 8347
rect 36461 8313 36495 8347
rect 38209 8313 38243 8347
rect 16037 8245 16071 8279
rect 21373 8245 21407 8279
rect 26985 8245 27019 8279
rect 28549 8245 28583 8279
rect 28641 8245 28675 8279
rect 31769 8245 31803 8279
rect 32505 8245 32539 8279
rect 32597 8245 32631 8279
rect 36553 8245 36587 8279
rect 37933 8245 37967 8279
rect 16129 8041 16163 8075
rect 19809 8041 19843 8075
rect 21741 8041 21775 8075
rect 21925 8041 21959 8075
rect 26065 8041 26099 8075
rect 28549 8041 28583 8075
rect 28917 8041 28951 8075
rect 32137 8041 32171 8075
rect 37841 8041 37875 8075
rect 38853 8041 38887 8075
rect 40969 8041 41003 8075
rect 16313 7973 16347 8007
rect 27537 7973 27571 8007
rect 28457 7973 28491 8007
rect 32321 7973 32355 8007
rect 32413 7973 32447 8007
rect 36737 7973 36771 8007
rect 12173 7905 12207 7939
rect 14105 7905 14139 7939
rect 15853 7905 15887 7939
rect 20269 7905 20303 7939
rect 21281 7905 21315 7939
rect 26709 7905 26743 7939
rect 27169 7905 27203 7939
rect 27445 7905 27479 7939
rect 28641 7905 28675 7939
rect 32229 7905 32263 7939
rect 32965 7905 32999 7939
rect 33425 7905 33459 7939
rect 36645 7905 36679 7939
rect 37013 7905 37047 7939
rect 16681 7837 16715 7871
rect 16865 7837 16899 7871
rect 17233 7837 17267 7871
rect 17877 7837 17911 7871
rect 17969 7837 18003 7871
rect 18153 7837 18187 7871
rect 20177 7837 20211 7871
rect 20637 7837 20671 7871
rect 26433 7837 26467 7871
rect 27077 7837 27111 7871
rect 28089 7837 28123 7871
rect 29561 7837 29595 7871
rect 32781 7837 32815 7871
rect 33057 7837 33091 7871
rect 36369 7837 36403 7871
rect 36553 7837 36587 7871
rect 36829 7837 36863 7871
rect 37657 7837 37691 7871
rect 38025 7837 38059 7871
rect 38761 7837 38795 7871
rect 39497 7837 39531 7871
rect 40049 7837 40083 7871
rect 40785 7837 40819 7871
rect 12449 7769 12483 7803
rect 14381 7769 14415 7803
rect 15945 7769 15979 7803
rect 21557 7769 21591 7803
rect 29837 7769 29871 7803
rect 13921 7701 13955 7735
rect 16145 7701 16179 7735
rect 16681 7701 16715 7735
rect 18061 7701 18095 7735
rect 21757 7701 21791 7735
rect 26525 7701 26559 7735
rect 31309 7701 31343 7735
rect 37105 7701 37139 7735
rect 38669 7701 38703 7735
rect 16129 7497 16163 7531
rect 16865 7497 16899 7531
rect 17509 7497 17543 7531
rect 20177 7497 20211 7531
rect 23305 7497 23339 7531
rect 28273 7497 28307 7531
rect 31861 7497 31895 7531
rect 33885 7497 33919 7531
rect 35817 7497 35851 7531
rect 36277 7497 36311 7531
rect 37105 7497 37139 7531
rect 15301 7429 15335 7463
rect 16037 7429 16071 7463
rect 22017 7429 22051 7463
rect 28457 7429 28491 7463
rect 35173 7429 35207 7463
rect 35378 7429 35412 7463
rect 36829 7429 36863 7463
rect 12817 7361 12851 7395
rect 13461 7361 13495 7395
rect 14013 7361 14047 7395
rect 16129 7361 16163 7395
rect 16221 7361 16255 7395
rect 16681 7361 16715 7395
rect 17049 7361 17083 7395
rect 17325 7361 17359 7395
rect 17417 7361 17451 7395
rect 17601 7361 17635 7395
rect 20361 7361 20395 7395
rect 20453 7361 20487 7395
rect 20545 7361 20579 7395
rect 21189 7361 21223 7395
rect 21373 7361 21407 7395
rect 23029 7361 23063 7395
rect 23213 7361 23247 7395
rect 26341 7361 26375 7395
rect 26985 7361 27019 7395
rect 27629 7361 27663 7395
rect 28089 7361 28123 7395
rect 28641 7361 28675 7395
rect 29929 7361 29963 7395
rect 30665 7361 30699 7395
rect 31309 7361 31343 7395
rect 32137 7361 32171 7395
rect 34529 7361 34563 7395
rect 36001 7361 36035 7395
rect 36553 7361 36587 7395
rect 36737 7361 36771 7395
rect 36921 7361 36955 7395
rect 38761 7361 38795 7395
rect 39129 7361 39163 7395
rect 12449 7293 12483 7327
rect 12909 7293 12943 7327
rect 16405 7293 16439 7327
rect 22753 7293 22787 7327
rect 26433 7293 26467 7327
rect 26525 7293 26559 7327
rect 30021 7293 30055 7327
rect 30205 7293 30239 7327
rect 32413 7293 32447 7327
rect 35633 7293 35667 7327
rect 35725 7293 35759 7327
rect 36093 7293 36127 7327
rect 37335 7293 37369 7327
rect 20729 7225 20763 7259
rect 25881 7225 25915 7259
rect 29561 7225 29595 7259
rect 17049 7157 17083 7191
rect 21373 7157 21407 7191
rect 23029 7157 23063 7191
rect 25973 7157 26007 7191
rect 27997 7157 28031 7191
rect 30481 7157 30515 7191
rect 33977 7157 34011 7191
rect 35357 7157 35391 7191
rect 35541 7157 35575 7191
rect 23961 6953 23995 6987
rect 25500 6953 25534 6987
rect 32321 6953 32355 6987
rect 36553 6953 36587 6987
rect 36829 6953 36863 6987
rect 15945 6885 15979 6919
rect 27353 6885 27387 6919
rect 33241 6885 33275 6919
rect 16589 6817 16623 6851
rect 20361 6817 20395 6851
rect 20913 6817 20947 6851
rect 21281 6817 21315 6851
rect 22477 6817 22511 6851
rect 24225 6817 24259 6851
rect 25237 6817 25271 6851
rect 30665 6817 30699 6851
rect 32873 6817 32907 6851
rect 34345 6817 34379 6851
rect 14749 6749 14783 6783
rect 16129 6749 16163 6783
rect 16221 6749 16255 6783
rect 18337 6749 18371 6783
rect 20545 6749 20579 6783
rect 21189 6749 21223 6783
rect 22017 6749 22051 6783
rect 27077 6749 27111 6783
rect 27353 6749 27387 6783
rect 27445 6749 27479 6783
rect 27629 6749 27663 6783
rect 30757 6749 30791 6783
rect 32689 6749 32723 6783
rect 34253 6749 34287 6783
rect 34437 6749 34471 6783
rect 35633 6749 35667 6783
rect 35725 6749 35759 6783
rect 36277 6749 36311 6783
rect 36737 6749 36771 6783
rect 36921 6749 36955 6783
rect 16497 6681 16531 6715
rect 18521 6681 18555 6715
rect 35449 6681 35483 6715
rect 36369 6681 36403 6715
rect 36553 6681 36587 6715
rect 14105 6613 14139 6647
rect 16313 6613 16347 6647
rect 18153 6613 18187 6647
rect 20637 6613 20671 6647
rect 20729 6613 20763 6647
rect 21557 6613 21591 6647
rect 26985 6613 27019 6647
rect 27169 6613 27203 6647
rect 27445 6613 27479 6647
rect 30389 6613 30423 6647
rect 32781 6613 32815 6647
rect 35725 6613 35759 6647
rect 13829 6409 13863 6443
rect 15209 6409 15243 6443
rect 15577 6409 15611 6443
rect 19717 6409 19751 6443
rect 20545 6409 20579 6443
rect 29101 6409 29135 6443
rect 30389 6409 30423 6443
rect 30573 6409 30607 6443
rect 30849 6409 30883 6443
rect 35909 6409 35943 6443
rect 14933 6341 14967 6375
rect 16037 6341 16071 6375
rect 30481 6341 30515 6375
rect 30757 6341 30791 6375
rect 13921 6273 13955 6307
rect 14105 6273 14139 6307
rect 14565 6273 14599 6307
rect 14657 6273 14691 6307
rect 14841 6273 14875 6307
rect 15117 6273 15151 6307
rect 15301 6273 15335 6307
rect 15761 6273 15795 6307
rect 17417 6273 17451 6307
rect 17601 6273 17635 6307
rect 19717 6273 19751 6307
rect 19901 6273 19935 6307
rect 20729 6273 20763 6307
rect 20913 6273 20947 6307
rect 27261 6273 27295 6307
rect 27721 6273 27755 6307
rect 28733 6273 28767 6307
rect 29745 6273 29779 6307
rect 31217 6273 31251 6307
rect 33609 6273 33643 6307
rect 36184 6273 36218 6307
rect 36277 6273 36311 6307
rect 12081 6205 12115 6239
rect 12357 6205 12391 6239
rect 15853 6205 15887 6239
rect 17693 6205 17727 6239
rect 19165 6205 19199 6239
rect 19441 6205 19475 6239
rect 21189 6205 21223 6239
rect 21281 6205 21315 6239
rect 21373 6205 21407 6239
rect 21465 6205 21499 6239
rect 21833 6205 21867 6239
rect 23305 6205 23339 6239
rect 23581 6205 23615 6239
rect 27353 6205 27387 6239
rect 28641 6205 28675 6239
rect 31309 6205 31343 6239
rect 33701 6205 33735 6239
rect 33977 6205 34011 6239
rect 36461 6205 36495 6239
rect 15485 6137 15519 6171
rect 27629 6137 27663 6171
rect 30205 6137 30239 6171
rect 13921 6069 13955 6103
rect 14841 6069 14875 6103
rect 15761 6069 15795 6103
rect 17509 6069 17543 6103
rect 21005 6069 21039 6103
rect 28365 6069 28399 6103
rect 29193 6069 29227 6103
rect 37013 6069 37047 6103
rect 13001 5865 13035 5899
rect 14565 5865 14599 5899
rect 14841 5865 14875 5899
rect 18153 5865 18187 5899
rect 18337 5865 18371 5899
rect 21005 5865 21039 5899
rect 21465 5865 21499 5899
rect 27445 5865 27479 5899
rect 29285 5865 29319 5899
rect 29561 5865 29595 5899
rect 31861 5865 31895 5899
rect 34529 5865 34563 5899
rect 36645 5865 36679 5899
rect 37473 5865 37507 5899
rect 14381 5797 14415 5831
rect 27537 5797 27571 5831
rect 37565 5797 37599 5831
rect 15485 5729 15519 5763
rect 15853 5729 15887 5763
rect 16313 5729 16347 5763
rect 18521 5729 18555 5763
rect 19257 5729 19291 5763
rect 21097 5729 21131 5763
rect 25973 5729 26007 5763
rect 28181 5729 28215 5763
rect 29009 5729 29043 5763
rect 30113 5729 30147 5763
rect 35265 5729 35299 5763
rect 36093 5729 36127 5763
rect 12817 5661 12851 5695
rect 13001 5661 13035 5695
rect 14105 5661 14139 5695
rect 14289 5661 14323 5695
rect 16037 5661 16071 5695
rect 17785 5661 17819 5695
rect 18613 5661 18647 5695
rect 21281 5661 21315 5695
rect 25697 5661 25731 5695
rect 27905 5661 27939 5695
rect 28733 5661 28767 5695
rect 32505 5661 32539 5695
rect 32781 5661 32815 5695
rect 37289 5661 37323 5695
rect 37933 5661 37967 5695
rect 14549 5593 14583 5627
rect 14749 5593 14783 5627
rect 16497 5593 16531 5627
rect 16681 5593 16715 5627
rect 18153 5593 18187 5627
rect 19533 5593 19567 5627
rect 30389 5593 30423 5627
rect 33057 5593 33091 5627
rect 14197 5525 14231 5559
rect 16221 5525 16255 5559
rect 18981 5525 19015 5559
rect 27997 5525 28031 5559
rect 28365 5525 28399 5559
rect 28825 5525 28859 5559
rect 31953 5525 31987 5559
rect 34713 5525 34747 5559
rect 36185 5525 36219 5559
rect 36277 5525 36311 5559
rect 36737 5525 36771 5559
rect 14565 5321 14599 5355
rect 14749 5321 14783 5355
rect 16681 5321 16715 5355
rect 19901 5321 19935 5355
rect 25421 5321 25455 5355
rect 29469 5321 29503 5355
rect 30941 5321 30975 5355
rect 31309 5321 31343 5355
rect 33333 5321 33367 5355
rect 33701 5321 33735 5355
rect 35541 5321 35575 5355
rect 16221 5253 16255 5287
rect 27997 5253 28031 5287
rect 31769 5253 31803 5287
rect 36676 5253 36710 5287
rect 12817 5185 12851 5219
rect 16497 5185 16531 5219
rect 16681 5185 16715 5219
rect 16865 5185 16899 5219
rect 20545 5185 20579 5219
rect 23673 5185 23707 5219
rect 36921 5185 36955 5219
rect 13093 5117 13127 5151
rect 23949 5117 23983 5151
rect 27721 5117 27755 5151
rect 31401 5117 31435 5151
rect 31585 5117 31619 5151
rect 33793 5117 33827 5151
rect 33977 5117 34011 5151
rect 34161 5117 34195 5151
rect 34805 4981 34839 5015
rect 23765 4777 23799 4811
rect 26157 4777 26191 4811
rect 27721 4777 27755 4811
rect 33241 4777 33275 4811
rect 34529 4777 34563 4811
rect 36461 4777 36495 4811
rect 15577 4641 15611 4675
rect 21189 4641 21223 4675
rect 22569 4641 22603 4675
rect 24409 4641 24443 4675
rect 31493 4641 31527 4675
rect 34713 4641 34747 4675
rect 34989 4641 35023 4675
rect 15301 4573 15335 4607
rect 15485 4573 15519 4607
rect 23581 4573 23615 4607
rect 23765 4573 23799 4607
rect 28825 4573 28859 4607
rect 30849 4573 30883 4607
rect 15393 4505 15427 4539
rect 15853 4505 15887 4539
rect 20913 4505 20947 4539
rect 24685 4505 24719 4539
rect 28089 4505 28123 4539
rect 30941 4505 30975 4539
rect 31769 4505 31803 4539
rect 17325 4437 17359 4471
rect 20545 4437 20579 4471
rect 21005 4437 21039 4471
rect 23213 4437 23247 4471
rect 22661 4233 22695 4267
rect 19993 4165 20027 4199
rect 22845 4165 22879 4199
rect 27261 4165 27295 4199
rect 16681 4097 16715 4131
rect 17325 4097 17359 4131
rect 22569 4097 22603 4131
rect 22937 4097 22971 4131
rect 23121 4097 23155 4131
rect 26341 4097 26375 4131
rect 26525 4097 26559 4131
rect 19717 4029 19751 4063
rect 22385 4029 22419 4063
rect 23305 4029 23339 4063
rect 23489 4029 23523 4063
rect 23765 4029 23799 4063
rect 25237 4029 25271 4063
rect 25605 4029 25639 4063
rect 26433 4029 26467 4063
rect 26985 4029 27019 4063
rect 28733 4029 28767 4063
rect 21465 3893 21499 3927
rect 21833 3893 21867 3927
rect 22845 3893 22879 3927
rect 26249 3893 26283 3927
rect 23397 3689 23431 3723
rect 25329 3689 25363 3723
rect 27997 3689 28031 3723
rect 32413 3689 32447 3723
rect 23489 3621 23523 3655
rect 19717 3553 19751 3587
rect 26249 3553 26283 3587
rect 30665 3553 30699 3587
rect 22385 3485 22419 3519
rect 23029 3485 23063 3519
rect 23213 3485 23247 3519
rect 23397 3485 23431 3519
rect 23489 3485 23523 3519
rect 23673 3485 23707 3519
rect 24685 3485 24719 3519
rect 25789 3485 25823 3519
rect 25973 3485 26007 3519
rect 28641 3485 28675 3519
rect 30297 3485 30331 3519
rect 19993 3417 20027 3451
rect 22109 3417 22143 3451
rect 22293 3417 22327 3451
rect 25881 3417 25915 3451
rect 26525 3417 26559 3451
rect 30941 3417 30975 3451
rect 21465 3349 21499 3383
rect 21925 3349 21959 3383
rect 28457 3349 28491 3383
rect 30481 3349 30515 3383
rect 20821 3145 20855 3179
rect 22017 3145 22051 3179
rect 22937 3145 22971 3179
rect 23397 3145 23431 3179
rect 23765 3145 23799 3179
rect 25697 3145 25731 3179
rect 31769 3145 31803 3179
rect 33885 3145 33919 3179
rect 22109 3077 22143 3111
rect 22661 3077 22695 3111
rect 24225 3077 24259 3111
rect 28365 3077 28399 3111
rect 32413 3077 32447 3111
rect 21005 3009 21039 3043
rect 22201 3009 22235 3043
rect 23949 3009 23983 3043
rect 28089 3009 28123 3043
rect 30021 3009 30055 3043
rect 34345 3009 34379 3043
rect 34437 3009 34471 3043
rect 35081 3009 35115 3043
rect 35265 3009 35299 3043
rect 36185 3009 36219 3043
rect 36277 3009 36311 3043
rect 36829 3009 36863 3043
rect 36921 3009 36955 3043
rect 37289 3009 37323 3043
rect 38117 3009 38151 3043
rect 38209 3009 38243 3043
rect 38761 3009 38795 3043
rect 38853 3009 38887 3043
rect 39405 3009 39439 3043
rect 39497 3009 39531 3043
rect 40049 3009 40083 3043
rect 40141 3009 40175 3043
rect 40693 3009 40727 3043
rect 40785 3009 40819 3043
rect 41337 3009 41371 3043
rect 41429 3009 41463 3043
rect 41981 3009 42015 3043
rect 42073 3009 42107 3043
rect 42441 3009 42475 3043
rect 43269 3009 43303 3043
rect 43361 3009 43395 3043
rect 43637 3009 43671 3043
rect 44373 3009 44407 3043
rect 44741 3009 44775 3043
rect 45109 3009 45143 3043
rect 21189 2941 21223 2975
rect 21281 2941 21315 2975
rect 21833 2941 21867 2975
rect 22293 2941 22327 2975
rect 22569 2941 22603 2975
rect 22778 2941 22812 2975
rect 23121 2941 23155 2975
rect 23305 2941 23339 2975
rect 30297 2941 30331 2975
rect 32137 2941 32171 2975
rect 35633 2941 35667 2975
rect 44833 2941 44867 2975
rect 21925 2873 21959 2907
rect 29837 2805 29871 2839
rect 34621 2805 34655 2839
rect 34897 2805 34931 2839
rect 35449 2805 35483 2839
rect 36001 2805 36035 2839
rect 36645 2805 36679 2839
rect 37473 2805 37507 2839
rect 37933 2805 37967 2839
rect 38577 2805 38611 2839
rect 39221 2805 39255 2839
rect 39865 2805 39899 2839
rect 40509 2805 40543 2839
rect 41153 2805 41187 2839
rect 41797 2805 41831 2839
rect 42625 2805 42659 2839
rect 43085 2805 43119 2839
rect 43821 2805 43855 2839
rect 44189 2805 44223 2839
rect 44557 2805 44591 2839
rect 19441 2601 19475 2635
rect 28917 2601 28951 2635
rect 29377 2601 29411 2635
rect 31033 2601 31067 2635
rect 22845 2533 22879 2567
rect 29745 2533 29779 2567
rect 30757 2533 30791 2567
rect 22661 2465 22695 2499
rect 28365 2465 28399 2499
rect 31493 2465 31527 2499
rect 35357 2465 35391 2499
rect 37289 2465 37323 2499
rect 42441 2465 42475 2499
rect 43637 2465 43671 2499
rect 19625 2397 19659 2431
rect 21005 2397 21039 2431
rect 21649 2397 21683 2431
rect 22201 2397 22235 2431
rect 22293 2397 22327 2431
rect 23029 2397 23063 2431
rect 23581 2397 23615 2431
rect 28457 2397 28491 2431
rect 28733 2397 28767 2431
rect 29193 2397 29227 2431
rect 29561 2397 29595 2431
rect 29837 2397 29871 2431
rect 30113 2397 30147 2431
rect 30297 2397 30331 2431
rect 30481 2397 30515 2431
rect 30665 2397 30699 2431
rect 30941 2397 30975 2431
rect 31217 2397 31251 2431
rect 22385 2329 22419 2363
rect 22477 2329 22511 2363
rect 29101 2329 29135 2363
rect 31309 2329 31343 2363
rect 19349 2261 19383 2295
rect 20821 2261 20855 2295
rect 21465 2261 21499 2295
rect 23397 2261 23431 2295
rect 28641 2261 28675 2295
<< metal1 >>
rect 1104 37562 58880 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 58880 37562
rect 1104 37488 58880 37510
rect 22554 37408 22560 37460
rect 22612 37448 22618 37460
rect 22741 37451 22799 37457
rect 22741 37448 22753 37451
rect 22612 37420 22753 37448
rect 22612 37408 22618 37420
rect 22741 37417 22753 37420
rect 22787 37417 22799 37451
rect 22741 37411 22799 37417
rect 23198 37408 23204 37460
rect 23256 37448 23262 37460
rect 23385 37451 23443 37457
rect 23385 37448 23397 37451
rect 23256 37420 23397 37448
rect 23256 37408 23262 37420
rect 23385 37417 23397 37420
rect 23431 37417 23443 37451
rect 23385 37411 23443 37417
rect 26418 37408 26424 37460
rect 26476 37448 26482 37460
rect 27065 37451 27123 37457
rect 27065 37448 27077 37451
rect 26476 37420 27077 37448
rect 26476 37408 26482 37420
rect 27065 37417 27077 37420
rect 27111 37417 27123 37451
rect 27065 37411 27123 37417
rect 28350 37408 28356 37460
rect 28408 37448 28414 37460
rect 28537 37451 28595 37457
rect 28537 37448 28549 37451
rect 28408 37420 28549 37448
rect 28408 37408 28414 37420
rect 28537 37417 28549 37420
rect 28583 37417 28595 37451
rect 28537 37411 28595 37417
rect 27341 37247 27399 37253
rect 27341 37213 27353 37247
rect 27387 37244 27399 37247
rect 31662 37244 31668 37256
rect 27387 37216 31668 37244
rect 27387 37213 27399 37216
rect 27341 37207 27399 37213
rect 31662 37204 31668 37216
rect 31720 37204 31726 37256
rect 23014 37136 23020 37188
rect 23072 37136 23078 37188
rect 23661 37179 23719 37185
rect 23661 37145 23673 37179
rect 23707 37176 23719 37179
rect 24210 37176 24216 37188
rect 23707 37148 24216 37176
rect 23707 37145 23719 37148
rect 23661 37139 23719 37145
rect 24210 37136 24216 37148
rect 24268 37136 24274 37188
rect 28813 37179 28871 37185
rect 28813 37145 28825 37179
rect 28859 37176 28871 37179
rect 29730 37176 29736 37188
rect 28859 37148 29736 37176
rect 28859 37145 28871 37148
rect 28813 37139 28871 37145
rect 29730 37136 29736 37148
rect 29788 37136 29794 37188
rect 1104 37018 58880 37040
rect 1104 36966 4874 37018
rect 4926 36966 4938 37018
rect 4990 36966 5002 37018
rect 5054 36966 5066 37018
rect 5118 36966 5130 37018
rect 5182 36966 35594 37018
rect 35646 36966 35658 37018
rect 35710 36966 35722 37018
rect 35774 36966 35786 37018
rect 35838 36966 35850 37018
rect 35902 36966 58880 37018
rect 1104 36944 58880 36966
rect 24486 36864 24492 36916
rect 24544 36904 24550 36916
rect 24949 36907 25007 36913
rect 24949 36904 24961 36907
rect 24544 36876 24961 36904
rect 24544 36864 24550 36876
rect 24949 36873 24961 36876
rect 24995 36873 25007 36907
rect 24949 36867 25007 36873
rect 25130 36864 25136 36916
rect 25188 36904 25194 36916
rect 25225 36907 25283 36913
rect 25225 36904 25237 36907
rect 25188 36876 25237 36904
rect 25188 36864 25194 36876
rect 25225 36873 25237 36876
rect 25271 36873 25283 36907
rect 25225 36867 25283 36873
rect 25685 36907 25743 36913
rect 25685 36873 25697 36907
rect 25731 36904 25743 36907
rect 25774 36904 25780 36916
rect 25731 36876 25780 36904
rect 25731 36873 25743 36876
rect 25685 36867 25743 36873
rect 25774 36864 25780 36876
rect 25832 36864 25838 36916
rect 27062 36864 27068 36916
rect 27120 36904 27126 36916
rect 27157 36907 27215 36913
rect 27157 36904 27169 36907
rect 27120 36876 27169 36904
rect 27120 36864 27126 36876
rect 27157 36873 27169 36876
rect 27203 36873 27215 36907
rect 27157 36867 27215 36873
rect 27617 36907 27675 36913
rect 27617 36873 27629 36907
rect 27663 36904 27675 36907
rect 27706 36904 27712 36916
rect 27663 36876 27712 36904
rect 27663 36873 27675 36876
rect 27617 36867 27675 36873
rect 27706 36864 27712 36876
rect 27764 36864 27770 36916
rect 28813 36907 28871 36913
rect 28813 36873 28825 36907
rect 28859 36904 28871 36907
rect 28994 36904 29000 36916
rect 28859 36876 29000 36904
rect 28859 36873 28871 36876
rect 28813 36867 28871 36873
rect 28994 36864 29000 36876
rect 29052 36864 29058 36916
rect 29457 36907 29515 36913
rect 29457 36873 29469 36907
rect 29503 36904 29515 36907
rect 29638 36904 29644 36916
rect 29503 36876 29644 36904
rect 29503 36873 29515 36876
rect 29457 36867 29515 36873
rect 29638 36864 29644 36876
rect 29696 36864 29702 36916
rect 30101 36907 30159 36913
rect 30101 36873 30113 36907
rect 30147 36904 30159 36907
rect 30282 36904 30288 36916
rect 30147 36876 30288 36904
rect 30147 36873 30159 36876
rect 30101 36867 30159 36873
rect 30282 36864 30288 36876
rect 30340 36864 30346 36916
rect 30837 36907 30895 36913
rect 30837 36873 30849 36907
rect 30883 36904 30895 36907
rect 30926 36904 30932 36916
rect 30883 36876 30932 36904
rect 30883 36873 30895 36876
rect 30837 36867 30895 36873
rect 30926 36864 30932 36876
rect 30984 36864 30990 36916
rect 31481 36907 31539 36913
rect 31481 36873 31493 36907
rect 31527 36904 31539 36907
rect 31570 36904 31576 36916
rect 31527 36876 31576 36904
rect 31527 36873 31539 36876
rect 31481 36867 31539 36873
rect 31570 36864 31576 36876
rect 31628 36864 31634 36916
rect 32214 36864 32220 36916
rect 32272 36904 32278 36916
rect 32309 36907 32367 36913
rect 32309 36904 32321 36907
rect 32272 36876 32321 36904
rect 32272 36864 32278 36876
rect 32309 36873 32321 36876
rect 32355 36873 32367 36907
rect 32309 36867 32367 36873
rect 32769 36907 32827 36913
rect 32769 36873 32781 36907
rect 32815 36904 32827 36907
rect 32858 36904 32864 36916
rect 32815 36876 32864 36904
rect 32815 36873 32827 36876
rect 32769 36867 32827 36873
rect 32858 36864 32864 36876
rect 32916 36864 32922 36916
rect 33413 36907 33471 36913
rect 33413 36873 33425 36907
rect 33459 36904 33471 36907
rect 33502 36904 33508 36916
rect 33459 36876 33508 36904
rect 33459 36873 33471 36876
rect 33413 36867 33471 36873
rect 33502 36864 33508 36876
rect 33560 36864 33566 36916
rect 34057 36907 34115 36913
rect 34057 36873 34069 36907
rect 34103 36904 34115 36907
rect 34146 36904 34152 36916
rect 34103 36876 34152 36904
rect 34103 36873 34115 36876
rect 34057 36867 34115 36873
rect 34146 36864 34152 36876
rect 34204 36864 34210 36916
rect 34701 36907 34759 36913
rect 34701 36873 34713 36907
rect 34747 36904 34759 36907
rect 34790 36904 34796 36916
rect 34747 36876 34796 36904
rect 34747 36873 34759 36876
rect 34701 36867 34759 36873
rect 34790 36864 34796 36876
rect 34848 36864 34854 36916
rect 35434 36864 35440 36916
rect 35492 36864 35498 36916
rect 35897 36907 35955 36913
rect 35897 36873 35909 36907
rect 35943 36904 35955 36907
rect 36078 36904 36084 36916
rect 35943 36876 36084 36904
rect 35943 36873 35955 36876
rect 35897 36867 35955 36873
rect 36078 36864 36084 36876
rect 36136 36864 36142 36916
rect 36541 36907 36599 36913
rect 36541 36873 36553 36907
rect 36587 36904 36599 36907
rect 36722 36904 36728 36916
rect 36587 36876 36728 36904
rect 36587 36873 36599 36876
rect 36541 36867 36599 36873
rect 36722 36864 36728 36876
rect 36780 36864 36786 36916
rect 37366 36864 37372 36916
rect 37424 36904 37430 36916
rect 37461 36907 37519 36913
rect 37461 36904 37473 36907
rect 37424 36876 37473 36904
rect 37424 36864 37430 36876
rect 37461 36873 37473 36876
rect 37507 36873 37519 36907
rect 37461 36867 37519 36873
rect 37921 36907 37979 36913
rect 37921 36873 37933 36907
rect 37967 36904 37979 36907
rect 38010 36904 38016 36916
rect 37967 36876 38016 36904
rect 37967 36873 37979 36876
rect 37921 36867 37979 36873
rect 38010 36864 38016 36876
rect 38068 36864 38074 36916
rect 38565 36907 38623 36913
rect 38565 36873 38577 36907
rect 38611 36904 38623 36907
rect 38654 36904 38660 36916
rect 38611 36876 38660 36904
rect 38611 36873 38623 36876
rect 38565 36867 38623 36873
rect 38654 36864 38660 36876
rect 38712 36864 38718 36916
rect 39209 36907 39267 36913
rect 39209 36873 39221 36907
rect 39255 36904 39267 36907
rect 39298 36904 39304 36916
rect 39255 36876 39304 36904
rect 39255 36873 39267 36876
rect 39209 36867 39267 36873
rect 39298 36864 39304 36876
rect 39356 36864 39362 36916
rect 39853 36907 39911 36913
rect 39853 36873 39865 36907
rect 39899 36904 39911 36907
rect 39942 36904 39948 36916
rect 39899 36876 39948 36904
rect 39899 36873 39911 36876
rect 39853 36867 39911 36873
rect 39942 36864 39948 36876
rect 40000 36864 40006 36916
rect 40497 36907 40555 36913
rect 40497 36873 40509 36907
rect 40543 36904 40555 36907
rect 40586 36904 40592 36916
rect 40543 36876 40592 36904
rect 40543 36873 40555 36876
rect 40497 36867 40555 36873
rect 40586 36864 40592 36876
rect 40644 36864 40650 36916
rect 41141 36907 41199 36913
rect 41141 36873 41153 36907
rect 41187 36904 41199 36907
rect 41230 36904 41236 36916
rect 41187 36876 41236 36904
rect 41187 36873 41199 36876
rect 41141 36867 41199 36873
rect 41230 36864 41236 36876
rect 41288 36864 41294 36916
rect 41785 36907 41843 36913
rect 41785 36873 41797 36907
rect 41831 36904 41843 36907
rect 41874 36904 41880 36916
rect 41831 36876 41880 36904
rect 41831 36873 41843 36876
rect 41785 36867 41843 36873
rect 41874 36864 41880 36876
rect 41932 36864 41938 36916
rect 42518 36864 42524 36916
rect 42576 36904 42582 36916
rect 42613 36907 42671 36913
rect 42613 36904 42625 36907
rect 42576 36876 42625 36904
rect 42576 36864 42582 36876
rect 42613 36873 42625 36876
rect 42659 36873 42671 36907
rect 42613 36867 42671 36873
rect 43073 36907 43131 36913
rect 43073 36873 43085 36907
rect 43119 36904 43131 36907
rect 43162 36904 43168 36916
rect 43119 36876 43168 36904
rect 43119 36873 43131 36876
rect 43073 36867 43131 36873
rect 43162 36864 43168 36876
rect 43220 36864 43226 36916
rect 43717 36907 43775 36913
rect 43717 36873 43729 36907
rect 43763 36904 43775 36907
rect 43806 36904 43812 36916
rect 43763 36876 43812 36904
rect 43763 36873 43775 36876
rect 43717 36867 43775 36873
rect 43806 36864 43812 36876
rect 43864 36864 43870 36916
rect 44361 36907 44419 36913
rect 44361 36873 44373 36907
rect 44407 36904 44419 36907
rect 44450 36904 44456 36916
rect 44407 36876 44456 36904
rect 44407 36873 44419 36876
rect 44361 36867 44419 36873
rect 44450 36864 44456 36876
rect 44508 36864 44514 36916
rect 45005 36907 45063 36913
rect 45005 36873 45017 36907
rect 45051 36904 45063 36907
rect 45094 36904 45100 36916
rect 45051 36876 45100 36904
rect 45051 36873 45063 36876
rect 45005 36867 45063 36873
rect 45094 36864 45100 36876
rect 45152 36864 45158 36916
rect 45649 36907 45707 36913
rect 45649 36873 45661 36907
rect 45695 36904 45707 36907
rect 45738 36904 45744 36916
rect 45695 36876 45744 36904
rect 45695 36873 45707 36876
rect 45649 36867 45707 36873
rect 45738 36864 45744 36876
rect 45796 36864 45802 36916
rect 46382 36864 46388 36916
rect 46440 36864 46446 36916
rect 46753 36907 46811 36913
rect 46753 36873 46765 36907
rect 46799 36904 46811 36907
rect 47026 36904 47032 36916
rect 46799 36876 47032 36904
rect 46799 36873 46811 36876
rect 46753 36867 46811 36873
rect 47026 36864 47032 36876
rect 47084 36864 47090 36916
rect 47121 36907 47179 36913
rect 47121 36873 47133 36907
rect 47167 36904 47179 36907
rect 47670 36904 47676 36916
rect 47167 36876 47676 36904
rect 47167 36873 47179 36876
rect 47121 36867 47179 36873
rect 47670 36864 47676 36876
rect 47728 36864 47734 36916
rect 24673 36771 24731 36777
rect 24673 36737 24685 36771
rect 24719 36768 24731 36771
rect 24765 36771 24823 36777
rect 24765 36768 24777 36771
rect 24719 36740 24777 36768
rect 24719 36737 24731 36740
rect 24673 36731 24731 36737
rect 24765 36737 24777 36740
rect 24811 36737 24823 36771
rect 24765 36731 24823 36737
rect 25314 36728 25320 36780
rect 25372 36768 25378 36780
rect 25409 36771 25467 36777
rect 25409 36768 25421 36771
rect 25372 36740 25421 36768
rect 25372 36728 25378 36740
rect 25409 36737 25421 36740
rect 25455 36737 25467 36771
rect 25409 36731 25467 36737
rect 25869 36771 25927 36777
rect 25869 36737 25881 36771
rect 25915 36768 25927 36771
rect 25961 36771 26019 36777
rect 25961 36768 25973 36771
rect 25915 36740 25973 36768
rect 25915 36737 25927 36740
rect 25869 36731 25927 36737
rect 25961 36737 25973 36740
rect 26007 36737 26019 36771
rect 25961 36731 26019 36737
rect 26789 36771 26847 36777
rect 26789 36737 26801 36771
rect 26835 36768 26847 36771
rect 26973 36771 27031 36777
rect 26973 36768 26985 36771
rect 26835 36740 26985 36768
rect 26835 36737 26847 36740
rect 26789 36731 26847 36737
rect 26973 36737 26985 36740
rect 27019 36737 27031 36771
rect 26973 36731 27031 36737
rect 27801 36771 27859 36777
rect 27801 36737 27813 36771
rect 27847 36768 27859 36771
rect 27893 36771 27951 36777
rect 27893 36768 27905 36771
rect 27847 36740 27905 36768
rect 27847 36737 27859 36740
rect 27801 36731 27859 36737
rect 27893 36737 27905 36740
rect 27939 36737 27951 36771
rect 27893 36731 27951 36737
rect 28997 36771 29055 36777
rect 28997 36737 29009 36771
rect 29043 36768 29055 36771
rect 29089 36771 29147 36777
rect 29089 36768 29101 36771
rect 29043 36740 29101 36768
rect 29043 36737 29055 36740
rect 28997 36731 29055 36737
rect 29089 36737 29101 36740
rect 29135 36737 29147 36771
rect 29089 36731 29147 36737
rect 29641 36771 29699 36777
rect 29641 36737 29653 36771
rect 29687 36768 29699 36771
rect 29733 36771 29791 36777
rect 29733 36768 29745 36771
rect 29687 36740 29745 36768
rect 29687 36737 29699 36740
rect 29641 36731 29699 36737
rect 29733 36737 29745 36740
rect 29779 36737 29791 36771
rect 29733 36731 29791 36737
rect 30285 36771 30343 36777
rect 30285 36737 30297 36771
rect 30331 36768 30343 36771
rect 30377 36771 30435 36777
rect 30377 36768 30389 36771
rect 30331 36740 30389 36768
rect 30331 36737 30343 36740
rect 30285 36731 30343 36737
rect 30377 36737 30389 36740
rect 30423 36737 30435 36771
rect 30377 36731 30435 36737
rect 31021 36771 31079 36777
rect 31021 36737 31033 36771
rect 31067 36768 31079 36771
rect 31113 36771 31171 36777
rect 31113 36768 31125 36771
rect 31067 36740 31125 36768
rect 31067 36737 31079 36740
rect 31021 36731 31079 36737
rect 31113 36737 31125 36740
rect 31159 36737 31171 36771
rect 31113 36731 31171 36737
rect 31665 36771 31723 36777
rect 31665 36737 31677 36771
rect 31711 36768 31723 36771
rect 31757 36771 31815 36777
rect 31757 36768 31769 36771
rect 31711 36740 31769 36768
rect 31711 36737 31723 36740
rect 31665 36731 31723 36737
rect 31757 36737 31769 36740
rect 31803 36737 31815 36771
rect 31757 36731 31815 36737
rect 32125 36771 32183 36777
rect 32125 36737 32137 36771
rect 32171 36768 32183 36771
rect 32214 36768 32220 36780
rect 32171 36740 32220 36768
rect 32171 36737 32183 36740
rect 32125 36731 32183 36737
rect 32214 36728 32220 36740
rect 32272 36728 32278 36780
rect 32953 36771 33011 36777
rect 32953 36737 32965 36771
rect 32999 36768 33011 36771
rect 33045 36771 33103 36777
rect 33045 36768 33057 36771
rect 32999 36740 33057 36768
rect 32999 36737 33011 36740
rect 32953 36731 33011 36737
rect 33045 36737 33057 36740
rect 33091 36737 33103 36771
rect 33045 36731 33103 36737
rect 33597 36771 33655 36777
rect 33597 36737 33609 36771
rect 33643 36768 33655 36771
rect 33689 36771 33747 36777
rect 33689 36768 33701 36771
rect 33643 36740 33701 36768
rect 33643 36737 33655 36740
rect 33597 36731 33655 36737
rect 33689 36737 33701 36740
rect 33735 36737 33747 36771
rect 33689 36731 33747 36737
rect 34241 36771 34299 36777
rect 34241 36737 34253 36771
rect 34287 36768 34299 36771
rect 34333 36771 34391 36777
rect 34333 36768 34345 36771
rect 34287 36740 34345 36768
rect 34287 36737 34299 36740
rect 34241 36731 34299 36737
rect 34333 36737 34345 36740
rect 34379 36737 34391 36771
rect 34333 36731 34391 36737
rect 34885 36771 34943 36777
rect 34885 36737 34897 36771
rect 34931 36768 34943 36771
rect 34977 36771 35035 36777
rect 34977 36768 34989 36771
rect 34931 36740 34989 36768
rect 34931 36737 34943 36740
rect 34885 36731 34943 36737
rect 34977 36737 34989 36740
rect 35023 36737 35035 36771
rect 34977 36731 35035 36737
rect 35253 36771 35311 36777
rect 35253 36737 35265 36771
rect 35299 36768 35311 36771
rect 35342 36768 35348 36780
rect 35299 36740 35348 36768
rect 35299 36737 35311 36740
rect 35253 36731 35311 36737
rect 35342 36728 35348 36740
rect 35400 36728 35406 36780
rect 36081 36771 36139 36777
rect 36081 36737 36093 36771
rect 36127 36768 36139 36771
rect 36173 36771 36231 36777
rect 36173 36768 36185 36771
rect 36127 36740 36185 36768
rect 36127 36737 36139 36740
rect 36081 36731 36139 36737
rect 36173 36737 36185 36740
rect 36219 36737 36231 36771
rect 36173 36731 36231 36737
rect 36725 36771 36783 36777
rect 36725 36737 36737 36771
rect 36771 36768 36783 36771
rect 36817 36771 36875 36777
rect 36817 36768 36829 36771
rect 36771 36740 36829 36768
rect 36771 36737 36783 36740
rect 36725 36731 36783 36737
rect 36817 36737 36829 36740
rect 36863 36737 36875 36771
rect 36817 36731 36875 36737
rect 37277 36771 37335 36777
rect 37277 36737 37289 36771
rect 37323 36768 37335 36771
rect 37366 36768 37372 36780
rect 37323 36740 37372 36768
rect 37323 36737 37335 36740
rect 37277 36731 37335 36737
rect 37366 36728 37372 36740
rect 37424 36728 37430 36780
rect 38105 36771 38163 36777
rect 38105 36737 38117 36771
rect 38151 36768 38163 36771
rect 38197 36771 38255 36777
rect 38197 36768 38209 36771
rect 38151 36740 38209 36768
rect 38151 36737 38163 36740
rect 38105 36731 38163 36737
rect 38197 36737 38209 36740
rect 38243 36737 38255 36771
rect 38197 36731 38255 36737
rect 38749 36771 38807 36777
rect 38749 36737 38761 36771
rect 38795 36768 38807 36771
rect 38841 36771 38899 36777
rect 38841 36768 38853 36771
rect 38795 36740 38853 36768
rect 38795 36737 38807 36740
rect 38749 36731 38807 36737
rect 38841 36737 38853 36740
rect 38887 36737 38899 36771
rect 38841 36731 38899 36737
rect 39393 36771 39451 36777
rect 39393 36737 39405 36771
rect 39439 36768 39451 36771
rect 39485 36771 39543 36777
rect 39485 36768 39497 36771
rect 39439 36740 39497 36768
rect 39439 36737 39451 36740
rect 39393 36731 39451 36737
rect 39485 36737 39497 36740
rect 39531 36737 39543 36771
rect 39485 36731 39543 36737
rect 40037 36771 40095 36777
rect 40037 36737 40049 36771
rect 40083 36768 40095 36771
rect 40129 36771 40187 36777
rect 40129 36768 40141 36771
rect 40083 36740 40141 36768
rect 40083 36737 40095 36740
rect 40037 36731 40095 36737
rect 40129 36737 40141 36740
rect 40175 36737 40187 36771
rect 40129 36731 40187 36737
rect 40681 36771 40739 36777
rect 40681 36737 40693 36771
rect 40727 36768 40739 36771
rect 40773 36771 40831 36777
rect 40773 36768 40785 36771
rect 40727 36740 40785 36768
rect 40727 36737 40739 36740
rect 40681 36731 40739 36737
rect 40773 36737 40785 36740
rect 40819 36737 40831 36771
rect 40773 36731 40831 36737
rect 41325 36771 41383 36777
rect 41325 36737 41337 36771
rect 41371 36768 41383 36771
rect 41417 36771 41475 36777
rect 41417 36768 41429 36771
rect 41371 36740 41429 36768
rect 41371 36737 41383 36740
rect 41325 36731 41383 36737
rect 41417 36737 41429 36740
rect 41463 36737 41475 36771
rect 41417 36731 41475 36737
rect 41969 36771 42027 36777
rect 41969 36737 41981 36771
rect 42015 36768 42027 36771
rect 42061 36771 42119 36777
rect 42061 36768 42073 36771
rect 42015 36740 42073 36768
rect 42015 36737 42027 36740
rect 41969 36731 42027 36737
rect 42061 36737 42073 36740
rect 42107 36737 42119 36771
rect 42061 36731 42119 36737
rect 42429 36771 42487 36777
rect 42429 36737 42441 36771
rect 42475 36768 42487 36771
rect 42518 36768 42524 36780
rect 42475 36740 42524 36768
rect 42475 36737 42487 36740
rect 42429 36731 42487 36737
rect 42518 36728 42524 36740
rect 42576 36728 42582 36780
rect 43257 36771 43315 36777
rect 43257 36737 43269 36771
rect 43303 36768 43315 36771
rect 43349 36771 43407 36777
rect 43349 36768 43361 36771
rect 43303 36740 43361 36768
rect 43303 36737 43315 36740
rect 43257 36731 43315 36737
rect 43349 36737 43361 36740
rect 43395 36737 43407 36771
rect 43349 36731 43407 36737
rect 43901 36771 43959 36777
rect 43901 36737 43913 36771
rect 43947 36768 43959 36771
rect 43993 36771 44051 36777
rect 43993 36768 44005 36771
rect 43947 36740 44005 36768
rect 43947 36737 43959 36740
rect 43901 36731 43959 36737
rect 43993 36737 44005 36740
rect 44039 36737 44051 36771
rect 43993 36731 44051 36737
rect 44545 36771 44603 36777
rect 44545 36737 44557 36771
rect 44591 36768 44603 36771
rect 44637 36771 44695 36777
rect 44637 36768 44649 36771
rect 44591 36740 44649 36768
rect 44591 36737 44603 36740
rect 44545 36731 44603 36737
rect 44637 36737 44649 36740
rect 44683 36737 44695 36771
rect 44637 36731 44695 36737
rect 45189 36771 45247 36777
rect 45189 36737 45201 36771
rect 45235 36768 45247 36771
rect 45281 36771 45339 36777
rect 45281 36768 45293 36771
rect 45235 36740 45293 36768
rect 45235 36737 45247 36740
rect 45189 36731 45247 36737
rect 45281 36737 45293 36740
rect 45327 36737 45339 36771
rect 45281 36731 45339 36737
rect 45833 36771 45891 36777
rect 45833 36737 45845 36771
rect 45879 36768 45891 36771
rect 45925 36771 45983 36777
rect 45925 36768 45937 36771
rect 45879 36740 45937 36768
rect 45879 36737 45891 36740
rect 45833 36731 45891 36737
rect 45925 36737 45937 36740
rect 45971 36737 45983 36771
rect 45925 36731 45983 36737
rect 46198 36728 46204 36780
rect 46256 36728 46262 36780
rect 46937 36771 46995 36777
rect 46937 36737 46949 36771
rect 46983 36737 46995 36771
rect 46937 36731 46995 36737
rect 47305 36771 47363 36777
rect 47305 36737 47317 36771
rect 47351 36768 47363 36771
rect 47857 36771 47915 36777
rect 47857 36768 47869 36771
rect 47351 36740 47869 36768
rect 47351 36737 47363 36740
rect 47305 36731 47363 36737
rect 47857 36737 47869 36740
rect 47903 36737 47915 36771
rect 47857 36731 47915 36737
rect 46952 36700 46980 36731
rect 47581 36703 47639 36709
rect 47581 36700 47593 36703
rect 46952 36672 47593 36700
rect 47581 36669 47593 36672
rect 47627 36669 47639 36703
rect 47581 36663 47639 36669
rect 1104 36474 58880 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 58880 36474
rect 1104 36400 58880 36422
rect 24210 36320 24216 36372
rect 24268 36320 24274 36372
rect 25314 36320 25320 36372
rect 25372 36320 25378 36372
rect 32214 36320 32220 36372
rect 32272 36320 32278 36372
rect 35253 36363 35311 36369
rect 35253 36329 35265 36363
rect 35299 36360 35311 36363
rect 35342 36360 35348 36372
rect 35299 36332 35348 36360
rect 35299 36329 35311 36332
rect 35253 36323 35311 36329
rect 35342 36320 35348 36332
rect 35400 36320 35406 36372
rect 37366 36320 37372 36372
rect 37424 36320 37430 36372
rect 42518 36320 42524 36372
rect 42576 36320 42582 36372
rect 46198 36320 46204 36372
rect 46256 36320 46262 36372
rect 24228 36224 24256 36320
rect 24949 36227 25007 36233
rect 24949 36224 24961 36227
rect 24228 36196 24961 36224
rect 24949 36193 24961 36196
rect 24995 36193 25007 36227
rect 24949 36187 25007 36193
rect 22094 36116 22100 36168
rect 22152 36156 22158 36168
rect 22833 36159 22891 36165
rect 22833 36156 22845 36159
rect 22152 36128 22845 36156
rect 22152 36116 22158 36128
rect 22833 36125 22845 36128
rect 22879 36125 22891 36159
rect 22833 36119 22891 36125
rect 29365 36159 29423 36165
rect 29365 36125 29377 36159
rect 29411 36156 29423 36159
rect 29411 36128 30328 36156
rect 29411 36125 29423 36128
rect 29365 36119 29423 36125
rect 23100 36091 23158 36097
rect 23100 36057 23112 36091
rect 23146 36088 23158 36091
rect 23290 36088 23296 36100
rect 23146 36060 23296 36088
rect 23146 36057 23158 36060
rect 23100 36051 23158 36057
rect 23290 36048 23296 36060
rect 23348 36048 23354 36100
rect 23566 36048 23572 36100
rect 23624 36088 23630 36100
rect 24397 36091 24455 36097
rect 24397 36088 24409 36091
rect 23624 36060 24409 36088
rect 23624 36048 23630 36060
rect 24397 36057 24409 36060
rect 24443 36057 24455 36091
rect 24397 36051 24455 36057
rect 28810 36048 28816 36100
rect 28868 36088 28874 36100
rect 29089 36091 29147 36097
rect 29089 36088 29101 36091
rect 28868 36060 29101 36088
rect 28868 36048 28874 36060
rect 29089 36057 29101 36060
rect 29135 36088 29147 36091
rect 29135 36060 29684 36088
rect 29135 36057 29147 36060
rect 29089 36051 29147 36057
rect 29546 35980 29552 36032
rect 29604 35980 29610 36032
rect 29656 36020 29684 36060
rect 29730 36048 29736 36100
rect 29788 36048 29794 36100
rect 29917 36091 29975 36097
rect 29917 36057 29929 36091
rect 29963 36088 29975 36091
rect 30009 36091 30067 36097
rect 30009 36088 30021 36091
rect 29963 36060 30021 36088
rect 29963 36057 29975 36060
rect 29917 36051 29975 36057
rect 30009 36057 30021 36060
rect 30055 36057 30067 36091
rect 30009 36051 30067 36057
rect 29932 36020 29960 36051
rect 30300 36029 30328 36128
rect 29656 35992 29960 36020
rect 30285 36023 30343 36029
rect 30285 35989 30297 36023
rect 30331 36020 30343 36023
rect 33318 36020 33324 36032
rect 30331 35992 33324 36020
rect 30331 35989 30343 35992
rect 30285 35983 30343 35989
rect 33318 35980 33324 35992
rect 33376 35980 33382 36032
rect 1104 35930 58880 35952
rect 1104 35878 4874 35930
rect 4926 35878 4938 35930
rect 4990 35878 5002 35930
rect 5054 35878 5066 35930
rect 5118 35878 5130 35930
rect 5182 35878 35594 35930
rect 35646 35878 35658 35930
rect 35710 35878 35722 35930
rect 35774 35878 35786 35930
rect 35838 35878 35850 35930
rect 35902 35878 58880 35930
rect 1104 35856 58880 35878
rect 23014 35776 23020 35828
rect 23072 35816 23078 35828
rect 23201 35819 23259 35825
rect 23201 35816 23213 35819
rect 23072 35788 23213 35816
rect 23072 35776 23078 35788
rect 23201 35785 23213 35788
rect 23247 35785 23259 35819
rect 23201 35779 23259 35785
rect 23290 35776 23296 35828
rect 23348 35776 23354 35828
rect 24121 35819 24179 35825
rect 24121 35785 24133 35819
rect 24167 35816 24179 35819
rect 25222 35816 25228 35828
rect 24167 35788 25228 35816
rect 24167 35785 24179 35788
rect 24121 35779 24179 35785
rect 24136 35748 24164 35779
rect 25222 35776 25228 35788
rect 25280 35816 25286 35828
rect 28810 35816 28816 35828
rect 25280 35788 28816 35816
rect 25280 35776 25286 35788
rect 28810 35776 28816 35788
rect 28868 35776 28874 35828
rect 29730 35776 29736 35828
rect 29788 35816 29794 35828
rect 29917 35819 29975 35825
rect 29917 35816 29929 35819
rect 29788 35788 29929 35816
rect 29788 35776 29794 35788
rect 29917 35785 29929 35788
rect 29963 35785 29975 35819
rect 29917 35779 29975 35785
rect 26694 35748 26700 35760
rect 23676 35720 24164 35748
rect 26542 35720 26700 35748
rect 23676 35692 23704 35720
rect 26694 35708 26700 35720
rect 26752 35748 26758 35760
rect 29270 35748 29276 35760
rect 26752 35720 29276 35748
rect 26752 35708 26758 35720
rect 29270 35708 29276 35720
rect 29328 35708 29334 35760
rect 21910 35640 21916 35692
rect 21968 35680 21974 35692
rect 22077 35683 22135 35689
rect 22077 35680 22089 35683
rect 21968 35652 22089 35680
rect 21968 35640 21974 35652
rect 22077 35649 22089 35652
rect 22123 35649 22135 35683
rect 22077 35643 22135 35649
rect 23566 35640 23572 35692
rect 23624 35640 23630 35692
rect 23658 35640 23664 35692
rect 23716 35640 23722 35692
rect 23750 35640 23756 35692
rect 23808 35640 23814 35692
rect 28810 35689 28816 35692
rect 23937 35683 23995 35689
rect 23937 35649 23949 35683
rect 23983 35649 23995 35683
rect 23937 35643 23995 35649
rect 28804 35643 28816 35689
rect 21821 35615 21879 35621
rect 21821 35581 21833 35615
rect 21867 35581 21879 35615
rect 21821 35575 21879 35581
rect 21836 35476 21864 35575
rect 23952 35544 23980 35643
rect 28810 35640 28816 35643
rect 28868 35640 28874 35692
rect 25038 35572 25044 35624
rect 25096 35572 25102 35624
rect 25314 35572 25320 35624
rect 25372 35572 25378 35624
rect 27798 35572 27804 35624
rect 27856 35612 27862 35624
rect 28537 35615 28595 35621
rect 28537 35612 28549 35615
rect 27856 35584 28549 35612
rect 27856 35572 27862 35584
rect 28537 35581 28549 35584
rect 28583 35581 28595 35615
rect 28537 35575 28595 35581
rect 23952 35516 25176 35544
rect 25148 35488 25176 35516
rect 22094 35476 22100 35488
rect 21836 35448 22100 35476
rect 22094 35436 22100 35448
rect 22152 35436 22158 35488
rect 25130 35436 25136 35488
rect 25188 35436 25194 35488
rect 26786 35436 26792 35488
rect 26844 35436 26850 35488
rect 1104 35386 58880 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 58880 35386
rect 1104 35312 58880 35334
rect 21910 35232 21916 35284
rect 21968 35232 21974 35284
rect 22278 35232 22284 35284
rect 22336 35272 22342 35284
rect 23569 35275 23627 35281
rect 23569 35272 23581 35275
rect 22336 35244 23581 35272
rect 22336 35232 22342 35244
rect 23569 35241 23581 35244
rect 23615 35272 23627 35275
rect 23658 35272 23664 35284
rect 23615 35244 23664 35272
rect 23615 35241 23627 35244
rect 23569 35235 23627 35241
rect 23658 35232 23664 35244
rect 23716 35232 23722 35284
rect 25225 35275 25283 35281
rect 25225 35241 25237 35275
rect 25271 35272 25283 35275
rect 25314 35272 25320 35284
rect 25271 35244 25320 35272
rect 25271 35241 25283 35244
rect 25225 35235 25283 35241
rect 25314 35232 25320 35244
rect 25372 35232 25378 35284
rect 26053 35275 26111 35281
rect 26053 35241 26065 35275
rect 26099 35272 26111 35275
rect 28549 35275 28607 35281
rect 28549 35272 28561 35275
rect 26099 35244 28561 35272
rect 26099 35241 26111 35244
rect 26053 35235 26111 35241
rect 28549 35241 28561 35244
rect 28595 35241 28607 35275
rect 28549 35235 28607 35241
rect 28810 35232 28816 35284
rect 28868 35272 28874 35284
rect 28905 35275 28963 35281
rect 28905 35272 28917 35275
rect 28868 35244 28917 35272
rect 28868 35232 28874 35244
rect 28905 35241 28917 35244
rect 28951 35241 28963 35275
rect 28905 35235 28963 35241
rect 29089 35275 29147 35281
rect 29089 35241 29101 35275
rect 29135 35272 29147 35275
rect 29546 35272 29552 35284
rect 29135 35244 29552 35272
rect 29135 35241 29147 35244
rect 29089 35235 29147 35241
rect 29546 35232 29552 35244
rect 29604 35232 29610 35284
rect 31662 35232 31668 35284
rect 31720 35232 31726 35284
rect 22741 35139 22799 35145
rect 22741 35136 22753 35139
rect 22204 35108 22753 35136
rect 18598 35028 18604 35080
rect 18656 35028 18662 35080
rect 22204 35077 22232 35108
rect 22741 35105 22753 35108
rect 22787 35105 22799 35139
rect 22741 35099 22799 35105
rect 23014 35096 23020 35148
rect 23072 35136 23078 35148
rect 23293 35139 23351 35145
rect 23293 35136 23305 35139
rect 23072 35108 23305 35136
rect 23072 35096 23078 35108
rect 23293 35105 23305 35108
rect 23339 35105 23351 35139
rect 23293 35099 23351 35105
rect 25424 35108 25820 35136
rect 22189 35071 22247 35077
rect 22189 35037 22201 35071
rect 22235 35037 22247 35071
rect 22189 35031 22247 35037
rect 22278 35028 22284 35080
rect 22336 35028 22342 35080
rect 22373 35071 22431 35077
rect 22373 35037 22385 35071
rect 22419 35068 22431 35071
rect 22462 35068 22468 35080
rect 22419 35040 22468 35068
rect 22419 35037 22431 35040
rect 22373 35031 22431 35037
rect 21821 35003 21879 35009
rect 21821 34969 21833 35003
rect 21867 35000 21879 35003
rect 22388 35000 22416 35031
rect 22462 35028 22468 35040
rect 22520 35028 22526 35080
rect 22557 35071 22615 35077
rect 22557 35037 22569 35071
rect 22603 35068 22615 35071
rect 22646 35068 22652 35080
rect 22603 35040 22652 35068
rect 22603 35037 22615 35040
rect 22557 35031 22615 35037
rect 22646 35028 22652 35040
rect 22704 35028 22710 35080
rect 24854 35028 24860 35080
rect 24912 35068 24918 35080
rect 25424 35077 25452 35108
rect 24949 35071 25007 35077
rect 24949 35068 24961 35071
rect 24912 35040 24961 35068
rect 24912 35028 24918 35040
rect 24949 35037 24961 35040
rect 24995 35037 25007 35071
rect 24949 35031 25007 35037
rect 25133 35071 25191 35077
rect 25133 35037 25145 35071
rect 25179 35037 25191 35071
rect 25133 35031 25191 35037
rect 25409 35071 25467 35077
rect 25409 35037 25421 35071
rect 25455 35037 25467 35071
rect 25409 35031 25467 35037
rect 21867 34972 22416 35000
rect 25148 35000 25176 35031
rect 25682 35028 25688 35080
rect 25740 35028 25746 35080
rect 25792 35077 25820 35108
rect 27798 35096 27804 35148
rect 27856 35136 27862 35148
rect 28810 35136 28816 35148
rect 27856 35108 28816 35136
rect 27856 35096 27862 35108
rect 28810 35096 28816 35108
rect 28868 35096 28874 35148
rect 25777 35071 25835 35077
rect 25777 35037 25789 35071
rect 25823 35068 25835 35071
rect 25866 35068 25872 35080
rect 25823 35040 25872 35068
rect 25823 35037 25835 35040
rect 25777 35031 25835 35037
rect 25866 35028 25872 35040
rect 25924 35028 25930 35080
rect 26050 35028 26056 35080
rect 26108 35028 26114 35080
rect 26237 35071 26295 35077
rect 26237 35037 26249 35071
rect 26283 35068 26295 35071
rect 26326 35068 26332 35080
rect 26283 35040 26332 35068
rect 26283 35037 26295 35040
rect 26237 35031 26295 35037
rect 26326 35028 26332 35040
rect 26384 35028 26390 35080
rect 26973 35071 27031 35077
rect 26973 35037 26985 35071
rect 27019 35068 27031 35071
rect 30374 35068 30380 35080
rect 27019 35040 27108 35068
rect 27019 35037 27031 35040
rect 26973 35031 27031 35037
rect 26418 35000 26424 35012
rect 25148 34972 26424 35000
rect 21867 34969 21879 34972
rect 21821 34963 21879 34969
rect 26418 34960 26424 34972
rect 26476 35000 26482 35012
rect 26786 35000 26792 35012
rect 26476 34972 26792 35000
rect 26476 34960 26482 34972
rect 26786 34960 26792 34972
rect 26844 34960 26850 35012
rect 27080 34944 27108 35040
rect 29196 35040 30380 35068
rect 29196 35000 29224 35040
rect 30374 35028 30380 35040
rect 30432 35028 30438 35080
rect 30650 35028 30656 35080
rect 30708 35068 30714 35080
rect 31021 35071 31079 35077
rect 31021 35068 31033 35071
rect 30708 35040 31033 35068
rect 30708 35028 30714 35040
rect 31021 35037 31033 35040
rect 31067 35037 31079 35071
rect 31021 35031 31079 35037
rect 31846 35028 31852 35080
rect 31904 35028 31910 35080
rect 28106 34972 29224 35000
rect 29270 34960 29276 35012
rect 29328 34960 29334 35012
rect 16850 34892 16856 34944
rect 16908 34932 16914 34944
rect 17957 34935 18015 34941
rect 17957 34932 17969 34935
rect 16908 34904 17969 34932
rect 16908 34892 16914 34904
rect 17957 34901 17969 34904
rect 18003 34901 18015 34935
rect 17957 34895 18015 34901
rect 25041 34935 25099 34941
rect 25041 34901 25053 34935
rect 25087 34932 25099 34935
rect 25593 34935 25651 34941
rect 25593 34932 25605 34935
rect 25087 34904 25605 34932
rect 25087 34901 25099 34904
rect 25041 34895 25099 34901
rect 25593 34901 25605 34904
rect 25639 34901 25651 34935
rect 25593 34895 25651 34901
rect 26329 34935 26387 34941
rect 26329 34901 26341 34935
rect 26375 34932 26387 34935
rect 26602 34932 26608 34944
rect 26375 34904 26608 34932
rect 26375 34901 26387 34904
rect 26329 34895 26387 34901
rect 26602 34892 26608 34904
rect 26660 34892 26666 34944
rect 27062 34892 27068 34944
rect 27120 34892 27126 34944
rect 29073 34935 29131 34941
rect 29073 34901 29085 34935
rect 29119 34932 29131 34935
rect 29178 34932 29184 34944
rect 29119 34904 29184 34932
rect 29119 34901 29131 34904
rect 29073 34895 29131 34901
rect 29178 34892 29184 34904
rect 29236 34892 29242 34944
rect 31202 34892 31208 34944
rect 31260 34892 31266 34944
rect 1104 34842 58880 34864
rect 1104 34790 4874 34842
rect 4926 34790 4938 34842
rect 4990 34790 5002 34842
rect 5054 34790 5066 34842
rect 5118 34790 5130 34842
rect 5182 34790 35594 34842
rect 35646 34790 35658 34842
rect 35710 34790 35722 34842
rect 35774 34790 35786 34842
rect 35838 34790 35850 34842
rect 35902 34790 58880 34842
rect 1104 34768 58880 34790
rect 24854 34688 24860 34740
rect 24912 34688 24918 34740
rect 25038 34688 25044 34740
rect 25096 34728 25102 34740
rect 27798 34728 27804 34740
rect 25096 34700 27804 34728
rect 25096 34688 25102 34700
rect 27798 34688 27804 34700
rect 27856 34688 27862 34740
rect 30852 34700 33088 34728
rect 18046 34620 18052 34672
rect 18104 34620 18110 34672
rect 16850 34552 16856 34604
rect 16908 34552 16914 34604
rect 21266 34552 21272 34604
rect 21324 34552 21330 34604
rect 22646 34552 22652 34604
rect 22704 34552 22710 34604
rect 24872 34592 24900 34688
rect 25682 34620 25688 34672
rect 25740 34660 25746 34672
rect 26053 34663 26111 34669
rect 26053 34660 26065 34663
rect 25740 34632 26065 34660
rect 25740 34620 25746 34632
rect 26053 34629 26065 34632
rect 26099 34629 26111 34663
rect 26697 34663 26755 34669
rect 26697 34660 26709 34663
rect 26053 34623 26111 34629
rect 26252 34632 26709 34660
rect 26252 34601 26280 34632
rect 26697 34629 26709 34632
rect 26743 34660 26755 34663
rect 26973 34663 27031 34669
rect 26973 34660 26985 34663
rect 26743 34632 26985 34660
rect 26743 34629 26755 34632
rect 26697 34623 26755 34629
rect 26973 34629 26985 34632
rect 27019 34629 27031 34663
rect 26973 34623 27031 34629
rect 27062 34620 27068 34672
rect 27120 34660 27126 34672
rect 27173 34663 27231 34669
rect 27173 34660 27185 34663
rect 27120 34632 27185 34660
rect 27120 34620 27126 34632
rect 27173 34629 27185 34632
rect 27219 34629 27231 34663
rect 27173 34623 27231 34629
rect 30374 34620 30380 34672
rect 30432 34660 30438 34672
rect 30852 34660 30880 34700
rect 33060 34660 33088 34700
rect 30432 34632 30958 34660
rect 33060 34632 33718 34660
rect 30432 34620 30438 34632
rect 25501 34595 25559 34601
rect 25501 34592 25513 34595
rect 16942 34484 16948 34536
rect 17000 34484 17006 34536
rect 17218 34484 17224 34536
rect 17276 34524 17282 34536
rect 17313 34527 17371 34533
rect 17313 34524 17325 34527
rect 17276 34496 17325 34524
rect 17276 34484 17282 34496
rect 17313 34493 17325 34496
rect 17359 34493 17371 34527
rect 17589 34527 17647 34533
rect 17589 34524 17601 34527
rect 17313 34487 17371 34493
rect 17420 34496 17601 34524
rect 17221 34391 17279 34397
rect 17221 34357 17233 34391
rect 17267 34388 17279 34391
rect 17420 34388 17448 34496
rect 17589 34493 17601 34496
rect 17635 34493 17647 34527
rect 17589 34487 17647 34493
rect 18138 34484 18144 34536
rect 18196 34524 18202 34536
rect 18598 34524 18604 34536
rect 18196 34496 18604 34524
rect 18196 34484 18202 34496
rect 18598 34484 18604 34496
rect 18656 34524 18662 34536
rect 19061 34527 19119 34533
rect 19061 34524 19073 34527
rect 18656 34496 19073 34524
rect 18656 34484 18662 34496
rect 19061 34493 19073 34496
rect 19107 34493 19119 34527
rect 19061 34487 19119 34493
rect 22094 34484 22100 34536
rect 22152 34524 22158 34536
rect 23106 34524 23112 34536
rect 22152 34496 23112 34524
rect 22152 34484 22158 34496
rect 23106 34484 23112 34496
rect 23164 34484 23170 34536
rect 23382 34484 23388 34536
rect 23440 34484 23446 34536
rect 24504 34524 24532 34578
rect 24872 34564 25513 34592
rect 25501 34561 25513 34564
rect 25547 34592 25559 34595
rect 26237 34595 26295 34601
rect 26237 34592 26249 34595
rect 25547 34564 26249 34592
rect 25547 34561 25559 34564
rect 25501 34555 25559 34561
rect 26237 34561 26249 34564
rect 26283 34561 26295 34595
rect 26237 34555 26295 34561
rect 26418 34552 26424 34604
rect 26476 34552 26482 34604
rect 26513 34595 26571 34601
rect 26513 34561 26525 34595
rect 26559 34561 26571 34595
rect 26513 34555 26571 34561
rect 24504 34496 26004 34524
rect 25976 34456 26004 34496
rect 26050 34484 26056 34536
rect 26108 34524 26114 34536
rect 26528 34524 26556 34555
rect 26786 34552 26792 34604
rect 26844 34552 26850 34604
rect 28810 34552 28816 34604
rect 28868 34592 28874 34604
rect 30193 34595 30251 34601
rect 30193 34592 30205 34595
rect 28868 34564 30205 34592
rect 28868 34552 28874 34564
rect 30193 34561 30205 34564
rect 30239 34561 30251 34595
rect 30193 34555 30251 34561
rect 26602 34524 26608 34536
rect 26108 34496 26464 34524
rect 26528 34496 26608 34524
rect 26108 34484 26114 34496
rect 26436 34456 26464 34496
rect 26602 34484 26608 34496
rect 26660 34484 26666 34536
rect 30466 34484 30472 34536
rect 30524 34484 30530 34536
rect 32306 34484 32312 34536
rect 32364 34524 32370 34536
rect 32953 34527 33011 34533
rect 32953 34524 32965 34527
rect 32364 34496 32965 34524
rect 32364 34484 32370 34496
rect 32953 34493 32965 34496
rect 32999 34493 33011 34527
rect 32953 34487 33011 34493
rect 33226 34484 33232 34536
rect 33284 34484 33290 34536
rect 34422 34484 34428 34536
rect 34480 34524 34486 34536
rect 34701 34527 34759 34533
rect 34701 34524 34713 34527
rect 34480 34496 34713 34524
rect 34480 34484 34486 34496
rect 34701 34493 34713 34496
rect 34747 34493 34759 34527
rect 34701 34487 34759 34493
rect 26513 34459 26571 34465
rect 26513 34456 26525 34459
rect 25976 34428 26280 34456
rect 26436 34428 26525 34456
rect 17267 34360 17448 34388
rect 17267 34357 17279 34360
rect 17221 34351 17279 34357
rect 21174 34348 21180 34400
rect 21232 34348 21238 34400
rect 24946 34348 24952 34400
rect 25004 34348 25010 34400
rect 26252 34388 26280 34428
rect 26513 34425 26525 34428
rect 26559 34425 26571 34459
rect 26513 34419 26571 34425
rect 26694 34388 26700 34400
rect 26252 34360 26700 34388
rect 26694 34348 26700 34360
rect 26752 34348 26758 34400
rect 26786 34348 26792 34400
rect 26844 34388 26850 34400
rect 27157 34391 27215 34397
rect 27157 34388 27169 34391
rect 26844 34360 27169 34388
rect 26844 34348 26850 34360
rect 27157 34357 27169 34360
rect 27203 34357 27215 34391
rect 27157 34351 27215 34357
rect 27246 34348 27252 34400
rect 27304 34388 27310 34400
rect 27341 34391 27399 34397
rect 27341 34388 27353 34391
rect 27304 34360 27353 34388
rect 27304 34348 27310 34360
rect 27341 34357 27353 34360
rect 27387 34357 27399 34391
rect 27341 34351 27399 34357
rect 31941 34391 31999 34397
rect 31941 34357 31953 34391
rect 31987 34388 31999 34391
rect 32122 34388 32128 34400
rect 31987 34360 32128 34388
rect 31987 34357 31999 34360
rect 31941 34351 31999 34357
rect 32122 34348 32128 34360
rect 32180 34348 32186 34400
rect 1104 34298 58880 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 58880 34298
rect 1104 34224 58880 34246
rect 18138 34184 18144 34196
rect 17604 34156 18144 34184
rect 17126 33940 17132 33992
rect 17184 33980 17190 33992
rect 17604 33980 17632 34156
rect 18138 34144 18144 34156
rect 18196 34144 18202 34196
rect 21266 34144 21272 34196
rect 21324 34144 21330 34196
rect 21729 34187 21787 34193
rect 21729 34153 21741 34187
rect 21775 34153 21787 34187
rect 21729 34147 21787 34153
rect 20254 34076 20260 34128
rect 20312 34076 20318 34128
rect 21634 34116 21640 34128
rect 20640 34088 21640 34116
rect 17681 34051 17739 34057
rect 17681 34017 17693 34051
rect 17727 34048 17739 34051
rect 18046 34048 18052 34060
rect 17727 34020 18052 34048
rect 17727 34017 17739 34020
rect 17681 34011 17739 34017
rect 18046 34008 18052 34020
rect 18104 34008 18110 34060
rect 19794 34008 19800 34060
rect 19852 34048 19858 34060
rect 20640 34057 20668 34088
rect 21634 34076 21640 34088
rect 21692 34116 21698 34128
rect 21744 34116 21772 34147
rect 25774 34144 25780 34196
rect 25832 34184 25838 34196
rect 25832 34156 26740 34184
rect 25832 34144 25838 34156
rect 21692 34088 21772 34116
rect 21692 34076 21698 34088
rect 26234 34076 26240 34128
rect 26292 34116 26298 34128
rect 26605 34119 26663 34125
rect 26605 34116 26617 34119
rect 26292 34088 26617 34116
rect 26292 34076 26298 34088
rect 26605 34085 26617 34088
rect 26651 34085 26663 34119
rect 26712 34116 26740 34156
rect 30466 34144 30472 34196
rect 30524 34184 30530 34196
rect 30561 34187 30619 34193
rect 30561 34184 30573 34187
rect 30524 34156 30573 34184
rect 30524 34144 30530 34156
rect 30561 34153 30573 34156
rect 30607 34153 30619 34187
rect 30561 34147 30619 34153
rect 30745 34187 30803 34193
rect 30745 34153 30757 34187
rect 30791 34153 30803 34187
rect 30745 34147 30803 34153
rect 30650 34116 30656 34128
rect 26712 34088 30656 34116
rect 26605 34079 26663 34085
rect 30650 34076 30656 34088
rect 30708 34076 30714 34128
rect 20625 34051 20683 34057
rect 20625 34048 20637 34051
rect 19852 34020 20637 34048
rect 19852 34008 19858 34020
rect 20625 34017 20637 34020
rect 20671 34017 20683 34051
rect 26145 34051 26203 34057
rect 26145 34048 26157 34051
rect 20625 34011 20683 34017
rect 24688 34020 26157 34048
rect 17773 33983 17831 33989
rect 17773 33980 17785 33983
rect 17184 33952 17785 33980
rect 17184 33940 17190 33952
rect 17773 33949 17785 33952
rect 17819 33949 17831 33983
rect 17773 33943 17831 33949
rect 17862 33940 17868 33992
rect 17920 33940 17926 33992
rect 17957 33983 18015 33989
rect 17957 33949 17969 33983
rect 18003 33980 18015 33983
rect 20533 33983 20591 33989
rect 18003 33952 18276 33980
rect 18003 33949 18015 33952
rect 17957 33943 18015 33949
rect 16942 33804 16948 33856
rect 17000 33844 17006 33856
rect 17770 33844 17776 33856
rect 17000 33816 17776 33844
rect 17000 33804 17006 33816
rect 17770 33804 17776 33816
rect 17828 33844 17834 33856
rect 17972 33844 18000 33943
rect 18248 33912 18276 33952
rect 20533 33949 20545 33983
rect 20579 33980 20591 33983
rect 22002 33980 22008 33992
rect 20579 33952 22008 33980
rect 20579 33949 20591 33952
rect 20533 33943 20591 33949
rect 22002 33940 22008 33952
rect 22060 33940 22066 33992
rect 23106 33940 23112 33992
rect 23164 33980 23170 33992
rect 24688 33989 24716 34020
rect 26145 34017 26157 34020
rect 26191 34048 26203 34051
rect 30282 34048 30288 34060
rect 26191 34020 30288 34048
rect 26191 34017 26203 34020
rect 26145 34011 26203 34017
rect 30282 34008 30288 34020
rect 30340 34008 30346 34060
rect 30760 34048 30788 34147
rect 31846 34144 31852 34196
rect 31904 34184 31910 34196
rect 31941 34187 31999 34193
rect 31941 34184 31953 34187
rect 31904 34156 31953 34184
rect 31904 34144 31910 34156
rect 31941 34153 31953 34156
rect 31987 34153 31999 34187
rect 31941 34147 31999 34153
rect 32674 34144 32680 34196
rect 32732 34184 32738 34196
rect 33045 34187 33103 34193
rect 33045 34184 33057 34187
rect 32732 34156 33057 34184
rect 32732 34144 32738 34156
rect 33045 34153 33057 34156
rect 33091 34153 33103 34187
rect 33045 34147 33103 34153
rect 31110 34076 31116 34128
rect 31168 34116 31174 34128
rect 32861 34119 32919 34125
rect 32861 34116 32873 34119
rect 31168 34088 32873 34116
rect 31168 34076 31174 34088
rect 32861 34085 32873 34088
rect 32907 34085 32919 34119
rect 33060 34116 33088 34147
rect 33226 34144 33232 34196
rect 33284 34184 33290 34196
rect 33965 34187 34023 34193
rect 33965 34184 33977 34187
rect 33284 34156 33977 34184
rect 33284 34144 33290 34156
rect 33965 34153 33977 34156
rect 34011 34153 34023 34187
rect 33965 34147 34023 34153
rect 33778 34116 33784 34128
rect 33060 34088 33784 34116
rect 32861 34079 32919 34085
rect 33778 34076 33784 34088
rect 33836 34076 33842 34128
rect 34333 34119 34391 34125
rect 34333 34116 34345 34119
rect 33980 34088 34345 34116
rect 31202 34048 31208 34060
rect 30760 34020 31208 34048
rect 31202 34008 31208 34020
rect 31260 34048 31266 34060
rect 32030 34048 32036 34060
rect 31260 34020 32036 34048
rect 31260 34008 31266 34020
rect 32030 34008 32036 34020
rect 32088 34008 32094 34060
rect 33042 34048 33048 34060
rect 32140 34020 33048 34048
rect 32140 33992 32168 34020
rect 23937 33983 23995 33989
rect 23937 33980 23949 33983
rect 23164 33952 23949 33980
rect 23164 33940 23170 33952
rect 23937 33949 23949 33952
rect 23983 33949 23995 33983
rect 23937 33943 23995 33949
rect 24673 33983 24731 33989
rect 24673 33949 24685 33983
rect 24719 33949 24731 33983
rect 24673 33943 24731 33949
rect 20257 33915 20315 33921
rect 20257 33912 20269 33915
rect 18248 33884 20269 33912
rect 20257 33881 20269 33884
rect 20303 33881 20315 33915
rect 20257 33875 20315 33881
rect 20441 33915 20499 33921
rect 20441 33881 20453 33915
rect 20487 33912 20499 33915
rect 21174 33912 21180 33924
rect 20487 33884 21180 33912
rect 20487 33881 20499 33884
rect 20441 33875 20499 33881
rect 17828 33816 18000 33844
rect 18141 33847 18199 33853
rect 17828 33804 17834 33816
rect 18141 33813 18153 33847
rect 18187 33844 18199 33847
rect 18322 33844 18328 33856
rect 18187 33816 18328 33844
rect 18187 33813 18199 33816
rect 18141 33807 18199 33813
rect 18322 33804 18328 33816
rect 18380 33804 18386 33856
rect 20272 33844 20300 33875
rect 21174 33872 21180 33884
rect 21232 33872 21238 33924
rect 21913 33915 21971 33921
rect 21913 33881 21925 33915
rect 21959 33912 21971 33915
rect 22554 33912 22560 33924
rect 21959 33884 22560 33912
rect 21959 33881 21971 33884
rect 21913 33875 21971 33881
rect 22554 33872 22560 33884
rect 22612 33872 22618 33924
rect 23952 33912 23980 33943
rect 25774 33940 25780 33992
rect 25832 33940 25838 33992
rect 26326 33940 26332 33992
rect 26384 33980 26390 33992
rect 26510 33980 26516 33992
rect 26384 33952 26516 33980
rect 26384 33940 26390 33952
rect 26510 33940 26516 33952
rect 26568 33940 26574 33992
rect 27154 33940 27160 33992
rect 27212 33980 27218 33992
rect 27341 33983 27399 33989
rect 27341 33980 27353 33983
rect 27212 33952 27353 33980
rect 27212 33940 27218 33952
rect 27341 33949 27353 33952
rect 27387 33949 27399 33983
rect 27341 33943 27399 33949
rect 30650 33940 30656 33992
rect 30708 33980 30714 33992
rect 31110 33980 31116 33992
rect 30708 33952 31116 33980
rect 30708 33940 30714 33952
rect 31110 33940 31116 33952
rect 31168 33940 31174 33992
rect 32122 33940 32128 33992
rect 32180 33940 32186 33992
rect 32508 33989 32536 34020
rect 33042 34008 33048 34020
rect 33100 34048 33106 34060
rect 33100 34020 33272 34048
rect 33100 34008 33106 34020
rect 32217 33983 32275 33989
rect 32217 33949 32229 33983
rect 32263 33980 32275 33983
rect 32493 33983 32551 33989
rect 32263 33952 32444 33980
rect 32263 33949 32275 33952
rect 32217 33943 32275 33949
rect 25038 33912 25044 33924
rect 23952 33884 25044 33912
rect 25038 33872 25044 33884
rect 25096 33912 25102 33924
rect 25409 33915 25467 33921
rect 25409 33912 25421 33915
rect 25096 33884 25421 33912
rect 25096 33872 25102 33884
rect 25409 33881 25421 33884
rect 25455 33881 25467 33915
rect 25409 33875 25467 33881
rect 26605 33915 26663 33921
rect 26605 33881 26617 33915
rect 26651 33912 26663 33915
rect 26789 33915 26847 33921
rect 26789 33912 26801 33915
rect 26651 33884 26801 33912
rect 26651 33881 26663 33884
rect 26605 33875 26663 33881
rect 26789 33881 26801 33884
rect 26835 33881 26847 33915
rect 26789 33875 26847 33881
rect 31662 33872 31668 33924
rect 31720 33912 31726 33924
rect 31941 33915 31999 33921
rect 31941 33912 31953 33915
rect 31720 33884 31953 33912
rect 31720 33872 31726 33884
rect 31941 33881 31953 33884
rect 31987 33881 31999 33915
rect 32309 33915 32367 33921
rect 32309 33912 32321 33915
rect 31941 33875 31999 33881
rect 32048 33884 32321 33912
rect 21545 33847 21603 33853
rect 21545 33844 21557 33847
rect 20272 33816 21557 33844
rect 21545 33813 21557 33816
rect 21591 33813 21603 33847
rect 21545 33807 21603 33813
rect 21713 33847 21771 33853
rect 21713 33813 21725 33847
rect 21759 33844 21771 33847
rect 22186 33844 22192 33856
rect 21759 33816 22192 33844
rect 21759 33813 21771 33816
rect 21713 33807 21771 33813
rect 22186 33804 22192 33816
rect 22244 33804 22250 33856
rect 25866 33804 25872 33856
rect 25924 33804 25930 33856
rect 26326 33804 26332 33856
rect 26384 33844 26390 33856
rect 26421 33847 26479 33853
rect 26421 33844 26433 33847
rect 26384 33816 26433 33844
rect 26384 33804 26390 33816
rect 26421 33813 26433 33816
rect 26467 33844 26479 33847
rect 27338 33844 27344 33856
rect 26467 33816 27344 33844
rect 26467 33813 26479 33816
rect 26421 33807 26479 33813
rect 27338 33804 27344 33816
rect 27396 33804 27402 33856
rect 30745 33847 30803 33853
rect 30745 33813 30757 33847
rect 30791 33844 30803 33847
rect 32048 33844 32076 33884
rect 32309 33881 32321 33884
rect 32355 33881 32367 33915
rect 32416 33912 32444 33952
rect 32493 33949 32505 33983
rect 32539 33949 32551 33983
rect 32493 33943 32551 33949
rect 32674 33940 32680 33992
rect 32732 33940 32738 33992
rect 32766 33940 32772 33992
rect 32824 33940 32830 33992
rect 33134 33912 33140 33924
rect 32416 33884 33140 33912
rect 32309 33875 32367 33881
rect 33134 33872 33140 33884
rect 33192 33872 33198 33924
rect 33244 33921 33272 34020
rect 33410 33940 33416 33992
rect 33468 33940 33474 33992
rect 33873 33983 33931 33989
rect 33873 33980 33885 33983
rect 33520 33952 33885 33980
rect 33229 33915 33287 33921
rect 33229 33881 33241 33915
rect 33275 33881 33287 33915
rect 33229 33875 33287 33881
rect 30791 33816 32076 33844
rect 30791 33813 30803 33816
rect 30745 33807 30803 33813
rect 32766 33804 32772 33856
rect 32824 33844 32830 33856
rect 33019 33847 33077 33853
rect 33019 33844 33031 33847
rect 32824 33816 33031 33844
rect 32824 33804 32830 33816
rect 33019 33813 33031 33816
rect 33065 33844 33077 33847
rect 33520 33844 33548 33952
rect 33873 33949 33885 33952
rect 33919 33980 33931 33983
rect 33980 33980 34008 34088
rect 34333 34085 34345 34088
rect 34379 34085 34391 34119
rect 34333 34079 34391 34085
rect 34422 34048 34428 34060
rect 33919 33952 34008 33980
rect 34072 34020 34428 34048
rect 33919 33949 33931 33952
rect 33873 33943 33931 33949
rect 33778 33872 33784 33924
rect 33836 33912 33842 33924
rect 34072 33912 34100 34020
rect 34422 34008 34428 34020
rect 34480 34008 34486 34060
rect 34149 33983 34207 33989
rect 34149 33949 34161 33983
rect 34195 33949 34207 33983
rect 34149 33943 34207 33949
rect 33836 33884 34100 33912
rect 33836 33872 33842 33884
rect 33065 33816 33548 33844
rect 33689 33847 33747 33853
rect 33065 33813 33077 33816
rect 33019 33807 33077 33813
rect 33689 33813 33701 33847
rect 33735 33844 33747 33847
rect 34164 33844 34192 33943
rect 33735 33816 34192 33844
rect 33735 33813 33747 33816
rect 33689 33807 33747 33813
rect 37090 33804 37096 33856
rect 37148 33804 37154 33856
rect 1104 33754 58880 33776
rect 1104 33702 4874 33754
rect 4926 33702 4938 33754
rect 4990 33702 5002 33754
rect 5054 33702 5066 33754
rect 5118 33702 5130 33754
rect 5182 33702 35594 33754
rect 35646 33702 35658 33754
rect 35710 33702 35722 33754
rect 35774 33702 35786 33754
rect 35838 33702 35850 33754
rect 35902 33702 58880 33754
rect 1104 33680 58880 33702
rect 17880 33612 21496 33640
rect 15930 33532 15936 33584
rect 15988 33572 15994 33584
rect 17880 33572 17908 33612
rect 17954 33572 17960 33584
rect 15988 33544 17960 33572
rect 15988 33532 15994 33544
rect 17954 33532 17960 33544
rect 18012 33532 18018 33584
rect 20165 33575 20223 33581
rect 20165 33541 20177 33575
rect 20211 33572 20223 33575
rect 20254 33572 20260 33584
rect 20211 33544 20260 33572
rect 20211 33541 20223 33544
rect 20165 33535 20223 33541
rect 20254 33532 20260 33544
rect 20312 33532 20318 33584
rect 21468 33572 21496 33612
rect 21634 33600 21640 33652
rect 21692 33600 21698 33652
rect 23382 33600 23388 33652
rect 23440 33640 23446 33652
rect 24397 33643 24455 33649
rect 24397 33640 24409 33643
rect 23440 33612 24409 33640
rect 23440 33600 23446 33612
rect 24397 33609 24409 33612
rect 24443 33609 24455 33643
rect 24397 33603 24455 33609
rect 26602 33600 26608 33652
rect 26660 33640 26666 33652
rect 27131 33643 27189 33649
rect 27131 33640 27143 33643
rect 26660 33612 27143 33640
rect 26660 33600 26666 33612
rect 27131 33609 27143 33612
rect 27177 33640 27189 33643
rect 27246 33640 27252 33652
rect 27177 33612 27252 33640
rect 27177 33609 27189 33612
rect 27131 33603 27189 33609
rect 27246 33600 27252 33612
rect 27304 33600 27310 33652
rect 32030 33600 32036 33652
rect 32088 33640 32094 33652
rect 33410 33640 33416 33652
rect 32088 33612 33416 33640
rect 32088 33600 32094 33612
rect 33410 33600 33416 33612
rect 33468 33640 33474 33652
rect 37093 33643 37151 33649
rect 33468 33612 35480 33640
rect 33468 33600 33474 33612
rect 22278 33572 22284 33584
rect 21390 33544 22284 33572
rect 22278 33532 22284 33544
rect 22336 33532 22342 33584
rect 24946 33572 24952 33584
rect 24688 33544 24952 33572
rect 16942 33464 16948 33516
rect 17000 33464 17006 33516
rect 17126 33464 17132 33516
rect 17184 33464 17190 33516
rect 22002 33464 22008 33516
rect 22060 33464 22066 33516
rect 22186 33464 22192 33516
rect 22244 33504 22250 33516
rect 24688 33513 24716 33544
rect 24946 33532 24952 33544
rect 25004 33532 25010 33584
rect 26694 33572 26700 33584
rect 26542 33544 26700 33572
rect 26694 33532 26700 33544
rect 26752 33532 26758 33584
rect 27338 33532 27344 33584
rect 27396 33532 27402 33584
rect 30374 33532 30380 33584
rect 30432 33532 30438 33584
rect 32784 33544 33640 33572
rect 23385 33507 23443 33513
rect 23385 33504 23397 33507
rect 22244 33476 23397 33504
rect 22244 33464 22250 33476
rect 23385 33473 23397 33476
rect 23431 33504 23443 33507
rect 24672 33507 24730 33513
rect 23431 33476 24164 33504
rect 23431 33473 23443 33476
rect 23385 33467 23443 33473
rect 17218 33396 17224 33448
rect 17276 33396 17282 33448
rect 17497 33439 17555 33445
rect 17497 33405 17509 33439
rect 17543 33436 17555 33439
rect 18230 33436 18236 33448
rect 17543 33408 18236 33436
rect 17543 33405 17555 33408
rect 17497 33399 17555 33405
rect 18230 33396 18236 33408
rect 18288 33396 18294 33448
rect 19889 33439 19947 33445
rect 19889 33405 19901 33439
rect 19935 33436 19947 33439
rect 20622 33436 20628 33448
rect 19935 33408 20628 33436
rect 19935 33405 19947 33408
rect 19889 33399 19947 33405
rect 20622 33396 20628 33408
rect 20680 33396 20686 33448
rect 22281 33439 22339 33445
rect 22281 33405 22293 33439
rect 22327 33436 22339 33439
rect 22465 33439 22523 33445
rect 22465 33436 22477 33439
rect 22327 33408 22477 33436
rect 22327 33405 22339 33408
rect 22281 33399 22339 33405
rect 22465 33405 22477 33408
rect 22511 33405 22523 33439
rect 22465 33399 22523 33405
rect 22554 33396 22560 33448
rect 22612 33436 22618 33448
rect 23017 33439 23075 33445
rect 23017 33436 23029 33439
rect 22612 33408 23029 33436
rect 22612 33396 22618 33408
rect 23017 33405 23029 33408
rect 23063 33436 23075 33439
rect 23201 33439 23259 33445
rect 23201 33436 23213 33439
rect 23063 33408 23213 33436
rect 23063 33405 23075 33408
rect 23017 33399 23075 33405
rect 23201 33405 23213 33408
rect 23247 33405 23259 33439
rect 23201 33399 23259 33405
rect 17034 33260 17040 33312
rect 17092 33260 17098 33312
rect 18046 33260 18052 33312
rect 18104 33300 18110 33312
rect 18966 33300 18972 33312
rect 18104 33272 18972 33300
rect 18104 33260 18110 33272
rect 18966 33260 18972 33272
rect 19024 33260 19030 33312
rect 21818 33260 21824 33312
rect 21876 33260 21882 33312
rect 23566 33260 23572 33312
rect 23624 33260 23630 33312
rect 24136 33300 24164 33476
rect 24672 33473 24684 33507
rect 24718 33473 24730 33507
rect 24672 33467 24730 33473
rect 24765 33507 24823 33513
rect 24765 33473 24777 33507
rect 24811 33504 24823 33507
rect 24854 33504 24860 33516
rect 24811 33476 24860 33504
rect 24811 33473 24823 33476
rect 24765 33467 24823 33473
rect 24854 33464 24860 33476
rect 24912 33464 24918 33516
rect 25038 33464 25044 33516
rect 25096 33464 25102 33516
rect 27798 33464 27804 33516
rect 27856 33504 27862 33516
rect 29089 33507 29147 33513
rect 29089 33504 29101 33507
rect 27856 33476 29101 33504
rect 27856 33464 27862 33476
rect 29089 33473 29101 33476
rect 29135 33473 29147 33507
rect 29089 33467 29147 33473
rect 31110 33464 31116 33516
rect 31168 33464 31174 33516
rect 32784 33513 32812 33544
rect 32769 33507 32827 33513
rect 32769 33473 32781 33507
rect 32815 33473 32827 33507
rect 32769 33467 32827 33473
rect 25314 33396 25320 33448
rect 25372 33396 25378 33448
rect 29365 33439 29423 33445
rect 29365 33405 29377 33439
rect 29411 33436 29423 33439
rect 30929 33439 30987 33445
rect 30929 33436 30941 33439
rect 29411 33408 30941 33436
rect 29411 33405 29423 33408
rect 29365 33399 29423 33405
rect 30929 33405 30941 33408
rect 30975 33405 30987 33439
rect 30929 33399 30987 33405
rect 31389 33439 31447 33445
rect 31389 33405 31401 33439
rect 31435 33436 31447 33439
rect 31662 33436 31668 33448
rect 31435 33408 31668 33436
rect 31435 33405 31447 33408
rect 31389 33399 31447 33405
rect 26789 33371 26847 33377
rect 26789 33337 26801 33371
rect 26835 33368 26847 33371
rect 26835 33340 27200 33368
rect 26835 33337 26847 33340
rect 26789 33331 26847 33337
rect 27172 33312 27200 33340
rect 30650 33328 30656 33380
rect 30708 33368 30714 33380
rect 31297 33371 31355 33377
rect 31297 33368 31309 33371
rect 30708 33340 31309 33368
rect 30708 33328 30714 33340
rect 31297 33337 31309 33340
rect 31343 33337 31355 33371
rect 31297 33331 31355 33337
rect 25958 33300 25964 33312
rect 24136 33272 25964 33300
rect 25958 33260 25964 33272
rect 26016 33300 26022 33312
rect 26973 33303 27031 33309
rect 26973 33300 26985 33303
rect 26016 33272 26985 33300
rect 26016 33260 26022 33272
rect 26973 33269 26985 33272
rect 27019 33269 27031 33303
rect 26973 33263 27031 33269
rect 27154 33260 27160 33312
rect 27212 33260 27218 33312
rect 30558 33260 30564 33312
rect 30616 33300 30622 33312
rect 30837 33303 30895 33309
rect 30837 33300 30849 33303
rect 30616 33272 30849 33300
rect 30616 33260 30622 33272
rect 30837 33269 30849 33272
rect 30883 33300 30895 33303
rect 31404 33300 31432 33399
rect 31662 33396 31668 33408
rect 31720 33436 31726 33448
rect 32784 33436 32812 33467
rect 32950 33464 32956 33516
rect 33008 33504 33014 33516
rect 33229 33507 33287 33513
rect 33229 33504 33241 33507
rect 33008 33476 33241 33504
rect 33008 33464 33014 33476
rect 33229 33473 33241 33476
rect 33275 33473 33287 33507
rect 33229 33467 33287 33473
rect 33505 33507 33563 33513
rect 33505 33473 33517 33507
rect 33551 33502 33563 33507
rect 33612 33502 33640 33544
rect 33551 33474 33640 33502
rect 33551 33473 33563 33474
rect 33505 33467 33563 33473
rect 31720 33408 32812 33436
rect 33137 33439 33195 33445
rect 31720 33396 31726 33408
rect 33137 33405 33149 33439
rect 33183 33436 33195 33439
rect 33686 33436 33692 33448
rect 33183 33408 33692 33436
rect 33183 33405 33195 33408
rect 33137 33399 33195 33405
rect 33686 33396 33692 33408
rect 33744 33396 33750 33448
rect 33781 33439 33839 33445
rect 33781 33405 33793 33439
rect 33827 33405 33839 33439
rect 33781 33399 33839 33405
rect 33796 33368 33824 33399
rect 33060 33340 33824 33368
rect 33060 33312 33088 33340
rect 30883 33272 31432 33300
rect 30883 33269 30895 33272
rect 30837 33263 30895 33269
rect 33042 33260 33048 33312
rect 33100 33260 33106 33312
rect 33410 33260 33416 33312
rect 33468 33260 33474 33312
rect 33778 33260 33784 33312
rect 33836 33260 33842 33312
rect 34054 33260 34060 33312
rect 34112 33260 34118 33312
rect 35452 33300 35480 33612
rect 37093 33609 37105 33643
rect 37139 33640 37151 33643
rect 37139 33612 37596 33640
rect 37139 33609 37151 33612
rect 37093 33603 37151 33609
rect 36909 33575 36967 33581
rect 36909 33541 36921 33575
rect 36955 33572 36967 33575
rect 37458 33572 37464 33584
rect 36955 33544 37464 33572
rect 36955 33541 36967 33544
rect 36909 33535 36967 33541
rect 37458 33532 37464 33544
rect 37516 33532 37522 33584
rect 37568 33581 37596 33612
rect 37553 33575 37611 33581
rect 37553 33541 37565 33575
rect 37599 33541 37611 33575
rect 37553 33535 37611 33541
rect 38654 33464 38660 33516
rect 38712 33464 38718 33516
rect 37274 33396 37280 33448
rect 37332 33396 37338 33448
rect 36541 33371 36599 33377
rect 36541 33337 36553 33371
rect 36587 33368 36599 33371
rect 36630 33368 36636 33380
rect 36587 33340 36636 33368
rect 36587 33337 36599 33340
rect 36541 33331 36599 33337
rect 36630 33328 36636 33340
rect 36688 33328 36694 33380
rect 36909 33303 36967 33309
rect 36909 33300 36921 33303
rect 35452 33272 36921 33300
rect 36909 33269 36921 33272
rect 36955 33300 36967 33303
rect 37366 33300 37372 33312
rect 36955 33272 37372 33300
rect 36955 33269 36967 33272
rect 36909 33263 36967 33269
rect 37366 33260 37372 33272
rect 37424 33260 37430 33312
rect 39022 33260 39028 33312
rect 39080 33260 39086 33312
rect 1104 33210 58880 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 58880 33210
rect 1104 33136 58880 33158
rect 18230 33056 18236 33108
rect 18288 33056 18294 33108
rect 19794 33056 19800 33108
rect 19852 33056 19858 33108
rect 22554 33056 22560 33108
rect 22612 33056 22618 33108
rect 23750 33096 23756 33108
rect 22664 33068 23756 33096
rect 18322 32988 18328 33040
rect 18380 32988 18386 33040
rect 16117 32963 16175 32969
rect 16117 32929 16129 32963
rect 16163 32929 16175 32963
rect 16117 32923 16175 32929
rect 13906 32852 13912 32904
rect 13964 32892 13970 32904
rect 14369 32895 14427 32901
rect 14369 32892 14381 32895
rect 13964 32864 14381 32892
rect 13964 32852 13970 32864
rect 14369 32861 14381 32864
rect 14415 32861 14427 32895
rect 16132 32892 16160 32923
rect 18966 32920 18972 32972
rect 19024 32960 19030 32972
rect 19521 32963 19579 32969
rect 19521 32960 19533 32963
rect 19024 32932 19533 32960
rect 19024 32920 19030 32932
rect 19521 32929 19533 32932
rect 19567 32929 19579 32963
rect 19521 32923 19579 32929
rect 21085 32963 21143 32969
rect 21085 32929 21097 32963
rect 21131 32960 21143 32963
rect 21818 32960 21824 32972
rect 21131 32932 21824 32960
rect 21131 32929 21143 32932
rect 21085 32923 21143 32929
rect 21818 32920 21824 32932
rect 21876 32920 21882 32972
rect 22278 32960 22284 32972
rect 22204 32932 22284 32960
rect 17037 32895 17095 32901
rect 17037 32892 17049 32895
rect 16132 32864 17049 32892
rect 14369 32855 14427 32861
rect 17037 32861 17049 32864
rect 17083 32892 17095 32895
rect 17862 32892 17868 32904
rect 17083 32864 17868 32892
rect 17083 32861 17095 32864
rect 17037 32855 17095 32861
rect 17862 32852 17868 32864
rect 17920 32852 17926 32904
rect 17957 32895 18015 32901
rect 17957 32861 17969 32895
rect 18003 32892 18015 32895
rect 18046 32892 18052 32904
rect 18003 32864 18052 32892
rect 18003 32861 18015 32864
rect 17957 32855 18015 32861
rect 18046 32852 18052 32864
rect 18104 32852 18110 32904
rect 18138 32852 18144 32904
rect 18196 32892 18202 32904
rect 19429 32895 19487 32901
rect 19429 32892 19441 32895
rect 18196 32864 19441 32892
rect 18196 32852 18202 32864
rect 19429 32861 19441 32864
rect 19475 32861 19487 32895
rect 19429 32855 19487 32861
rect 20622 32852 20628 32904
rect 20680 32892 20686 32904
rect 20809 32895 20867 32901
rect 20809 32892 20821 32895
rect 20680 32864 20821 32892
rect 20680 32852 20686 32864
rect 20809 32861 20821 32864
rect 20855 32861 20867 32895
rect 22204 32878 22232 32932
rect 22278 32920 22284 32932
rect 22336 32960 22342 32972
rect 22664 32960 22692 33068
rect 23750 33056 23756 33068
rect 23808 33056 23814 33108
rect 24121 33099 24179 33105
rect 24121 33065 24133 33099
rect 24167 33096 24179 33099
rect 24949 33099 25007 33105
rect 24167 33068 24716 33096
rect 24167 33065 24179 33068
rect 24121 33059 24179 33065
rect 23566 32988 23572 33040
rect 23624 33028 23630 33040
rect 23937 33031 23995 33037
rect 23937 33028 23949 33031
rect 23624 33000 23949 33028
rect 23624 32988 23630 33000
rect 23937 32997 23949 33000
rect 23983 33028 23995 33031
rect 24688 33028 24716 33068
rect 24949 33065 24961 33099
rect 24995 33096 25007 33099
rect 25133 33099 25191 33105
rect 25133 33096 25145 33099
rect 24995 33068 25145 33096
rect 24995 33065 25007 33068
rect 24949 33059 25007 33065
rect 25133 33065 25145 33068
rect 25179 33096 25191 33099
rect 25222 33096 25228 33108
rect 25179 33068 25228 33096
rect 25179 33065 25191 33068
rect 25133 33059 25191 33065
rect 25222 33056 25228 33068
rect 25280 33056 25286 33108
rect 25314 33056 25320 33108
rect 25372 33096 25378 33108
rect 25777 33099 25835 33105
rect 25777 33096 25789 33099
rect 25372 33068 25789 33096
rect 25372 33056 25378 33068
rect 25777 33065 25789 33068
rect 25823 33065 25835 33099
rect 25777 33059 25835 33065
rect 26053 33099 26111 33105
rect 26053 33065 26065 33099
rect 26099 33096 26111 33099
rect 26326 33096 26332 33108
rect 26099 33068 26332 33096
rect 26099 33065 26111 33068
rect 26053 33059 26111 33065
rect 26326 33056 26332 33068
rect 26384 33056 26390 33108
rect 30377 33099 30435 33105
rect 30377 33065 30389 33099
rect 30423 33096 30435 33099
rect 31110 33096 31116 33108
rect 30423 33068 31116 33096
rect 30423 33065 30435 33068
rect 30377 33059 30435 33065
rect 31110 33056 31116 33068
rect 31168 33056 31174 33108
rect 33134 33056 33140 33108
rect 33192 33096 33198 33108
rect 33229 33099 33287 33105
rect 33229 33096 33241 33099
rect 33192 33068 33241 33096
rect 33192 33056 33198 33068
rect 33229 33065 33241 33068
rect 33275 33065 33287 33099
rect 33229 33059 33287 33065
rect 33962 33056 33968 33108
rect 34020 33096 34026 33108
rect 34057 33099 34115 33105
rect 34057 33096 34069 33099
rect 34020 33068 34069 33096
rect 34020 33056 34026 33068
rect 34057 33065 34069 33068
rect 34103 33065 34115 33099
rect 34057 33059 34115 33065
rect 37458 33056 37464 33108
rect 37516 33096 37522 33108
rect 38013 33099 38071 33105
rect 38013 33096 38025 33099
rect 37516 33068 38025 33096
rect 37516 33056 37522 33068
rect 38013 33065 38025 33068
rect 38059 33065 38071 33099
rect 38013 33059 38071 33065
rect 25682 33028 25688 33040
rect 23983 33000 24440 33028
rect 24688 33000 25688 33028
rect 23983 32997 23995 33000
rect 23937 32991 23995 32997
rect 24412 32969 24440 33000
rect 25682 32988 25688 33000
rect 25740 32988 25746 33040
rect 32766 32988 32772 33040
rect 32824 33028 32830 33040
rect 34241 33031 34299 33037
rect 34241 33028 34253 33031
rect 32824 33000 34253 33028
rect 32824 32988 32830 33000
rect 34241 32997 34253 33000
rect 34287 32997 34299 33031
rect 34241 32991 34299 32997
rect 37182 32988 37188 33040
rect 37240 32988 37246 33040
rect 24397 32963 24455 32969
rect 22336 32932 22692 32960
rect 23216 32932 23704 32960
rect 22336 32920 22342 32932
rect 23216 32901 23244 32932
rect 23201 32895 23259 32901
rect 20809 32855 20867 32861
rect 23201 32861 23213 32895
rect 23247 32861 23259 32895
rect 23201 32855 23259 32861
rect 23385 32895 23443 32901
rect 23385 32861 23397 32895
rect 23431 32892 23443 32895
rect 23566 32892 23572 32904
rect 23431 32864 23572 32892
rect 23431 32861 23443 32864
rect 23385 32855 23443 32861
rect 23566 32852 23572 32864
rect 23624 32852 23630 32904
rect 23676 32901 23704 32932
rect 24397 32929 24409 32963
rect 24443 32929 24455 32963
rect 26234 32960 26240 32972
rect 24397 32923 24455 32929
rect 25792 32932 26240 32960
rect 23661 32895 23719 32901
rect 23661 32861 23673 32895
rect 23707 32892 23719 32895
rect 23842 32892 23848 32904
rect 23707 32864 23848 32892
rect 23707 32861 23719 32864
rect 23661 32855 23719 32861
rect 23842 32852 23848 32864
rect 23900 32892 23906 32904
rect 24765 32895 24823 32901
rect 24765 32892 24777 32895
rect 23900 32864 24777 32892
rect 23900 32852 23906 32864
rect 24765 32861 24777 32864
rect 24811 32861 24823 32895
rect 24765 32855 24823 32861
rect 24854 32852 24860 32904
rect 24912 32892 24918 32904
rect 25792 32901 25820 32932
rect 26234 32920 26240 32932
rect 26292 32920 26298 32972
rect 27798 32920 27804 32972
rect 27856 32920 27862 32972
rect 35805 32963 35863 32969
rect 32876 32932 34376 32960
rect 25501 32895 25559 32901
rect 25501 32892 25513 32895
rect 24912 32864 25513 32892
rect 24912 32852 24918 32864
rect 25501 32861 25513 32864
rect 25547 32861 25559 32895
rect 25501 32855 25559 32861
rect 25777 32895 25835 32901
rect 25777 32861 25789 32895
rect 25823 32861 25835 32895
rect 25777 32855 25835 32861
rect 14642 32784 14648 32836
rect 14700 32784 14706 32836
rect 15930 32824 15936 32836
rect 15870 32796 15936 32824
rect 15930 32784 15936 32796
rect 15988 32784 15994 32836
rect 17770 32784 17776 32836
rect 17828 32784 17834 32836
rect 16298 32716 16304 32768
rect 16356 32756 16362 32768
rect 16393 32759 16451 32765
rect 16393 32756 16405 32759
rect 16356 32728 16405 32756
rect 16356 32716 16362 32728
rect 16393 32725 16405 32728
rect 16439 32725 16451 32759
rect 16393 32719 16451 32725
rect 16482 32716 16488 32768
rect 16540 32756 16546 32768
rect 17880 32765 17908 32852
rect 18230 32784 18236 32836
rect 18288 32824 18294 32836
rect 18693 32827 18751 32833
rect 18693 32824 18705 32827
rect 18288 32796 18705 32824
rect 18288 32784 18294 32796
rect 18693 32793 18705 32796
rect 18739 32793 18751 32827
rect 19889 32827 19947 32833
rect 19889 32824 19901 32827
rect 18693 32787 18751 32793
rect 18800 32796 19901 32824
rect 17589 32759 17647 32765
rect 17589 32756 17601 32759
rect 16540 32728 17601 32756
rect 16540 32716 16546 32728
rect 17589 32725 17601 32728
rect 17635 32725 17647 32759
rect 17589 32719 17647 32725
rect 17865 32759 17923 32765
rect 17865 32725 17877 32759
rect 17911 32756 17923 32759
rect 18800 32756 18828 32796
rect 19889 32793 19901 32796
rect 19935 32793 19947 32827
rect 23293 32827 23351 32833
rect 23293 32824 23305 32827
rect 19889 32787 19947 32793
rect 22480 32796 23305 32824
rect 17911 32728 18828 32756
rect 17911 32725 17923 32728
rect 17865 32719 17923 32725
rect 19242 32716 19248 32768
rect 19300 32716 19306 32768
rect 22002 32716 22008 32768
rect 22060 32756 22066 32768
rect 22480 32756 22508 32796
rect 23293 32793 23305 32796
rect 23339 32793 23351 32827
rect 23293 32787 23351 32793
rect 22060 32728 22508 32756
rect 22060 32716 22066 32728
rect 24578 32716 24584 32768
rect 24636 32716 24642 32768
rect 25516 32756 25544 32855
rect 25958 32852 25964 32904
rect 26016 32852 26022 32904
rect 30558 32852 30564 32904
rect 30616 32852 30622 32904
rect 30650 32852 30656 32904
rect 30708 32852 30714 32904
rect 30745 32895 30803 32901
rect 30745 32861 30757 32895
rect 30791 32861 30803 32895
rect 30745 32855 30803 32861
rect 30929 32895 30987 32901
rect 30929 32861 30941 32895
rect 30975 32892 30987 32895
rect 32766 32892 32772 32904
rect 30975 32864 32772 32892
rect 30975 32861 30987 32864
rect 30929 32855 30987 32861
rect 26786 32784 26792 32836
rect 26844 32784 26850 32836
rect 27522 32784 27528 32836
rect 27580 32784 27586 32836
rect 28902 32784 28908 32836
rect 28960 32824 28966 32836
rect 30377 32827 30435 32833
rect 30377 32824 30389 32827
rect 28960 32796 30389 32824
rect 28960 32784 28966 32796
rect 30377 32793 30389 32796
rect 30423 32824 30435 32827
rect 30760 32824 30788 32855
rect 32766 32852 32772 32864
rect 32824 32852 32830 32904
rect 32582 32824 32588 32836
rect 30423 32796 32588 32824
rect 30423 32793 30435 32796
rect 30377 32787 30435 32793
rect 32582 32784 32588 32796
rect 32640 32824 32646 32836
rect 32876 32824 32904 32932
rect 33413 32895 33471 32901
rect 33413 32886 33425 32895
rect 32640 32796 32904 32824
rect 33336 32861 33425 32886
rect 33459 32861 33471 32895
rect 33336 32858 33471 32861
rect 32640 32784 32646 32796
rect 25866 32756 25872 32768
rect 25516 32728 25872 32756
rect 25866 32716 25872 32728
rect 25924 32756 25930 32768
rect 27154 32756 27160 32768
rect 25924 32728 27160 32756
rect 25924 32716 25930 32728
rect 27154 32716 27160 32728
rect 27212 32716 27218 32768
rect 30834 32716 30840 32768
rect 30892 32716 30898 32768
rect 33336 32756 33364 32858
rect 33413 32855 33471 32858
rect 33502 32852 33508 32904
rect 33560 32852 33566 32904
rect 33594 32852 33600 32904
rect 33652 32892 33658 32904
rect 33689 32895 33747 32901
rect 33689 32892 33701 32895
rect 33652 32864 33701 32892
rect 33652 32852 33658 32864
rect 33689 32861 33701 32864
rect 33735 32861 33747 32895
rect 33689 32855 33747 32861
rect 33778 32852 33784 32904
rect 33836 32852 33842 32904
rect 34238 32892 34244 32904
rect 33888 32864 34244 32892
rect 33888 32833 33916 32864
rect 34238 32852 34244 32864
rect 34296 32852 34302 32904
rect 34348 32901 34376 32932
rect 35805 32929 35817 32963
rect 35851 32960 35863 32963
rect 36814 32960 36820 32972
rect 35851 32932 36820 32960
rect 35851 32929 35863 32932
rect 35805 32923 35863 32929
rect 36814 32920 36820 32932
rect 36872 32960 36878 32972
rect 37200 32960 37228 32988
rect 36872 32932 37228 32960
rect 36872 32920 36878 32932
rect 34333 32895 34391 32901
rect 34333 32861 34345 32895
rect 34379 32861 34391 32895
rect 34333 32855 34391 32861
rect 34514 32852 34520 32904
rect 34572 32852 34578 32904
rect 37090 32852 37096 32904
rect 37148 32892 37154 32904
rect 37148 32864 37780 32892
rect 37148 32852 37154 32864
rect 33873 32827 33931 32833
rect 33873 32793 33885 32827
rect 33919 32793 33931 32827
rect 33873 32787 33931 32793
rect 34089 32827 34147 32833
rect 34089 32793 34101 32827
rect 34135 32824 34147 32827
rect 35986 32824 35992 32836
rect 34135 32796 35992 32824
rect 34135 32793 34147 32796
rect 34089 32787 34147 32793
rect 35986 32784 35992 32796
rect 36044 32784 36050 32836
rect 36078 32784 36084 32836
rect 36136 32784 36142 32836
rect 37645 32827 37703 32833
rect 37645 32824 37657 32827
rect 37384 32796 37657 32824
rect 33686 32756 33692 32768
rect 33336 32728 33692 32756
rect 33686 32716 33692 32728
rect 33744 32716 33750 32768
rect 34425 32759 34483 32765
rect 34425 32725 34437 32759
rect 34471 32756 34483 32759
rect 36262 32756 36268 32768
rect 34471 32728 36268 32756
rect 34471 32725 34483 32728
rect 34425 32719 34483 32725
rect 36262 32716 36268 32728
rect 36320 32716 36326 32768
rect 36722 32716 36728 32768
rect 36780 32756 36786 32768
rect 37384 32756 37412 32796
rect 37645 32793 37657 32796
rect 37691 32793 37703 32827
rect 37645 32787 37703 32793
rect 36780 32728 37412 32756
rect 36780 32716 36786 32728
rect 37550 32716 37556 32768
rect 37608 32716 37614 32768
rect 37752 32756 37780 32864
rect 37826 32784 37832 32836
rect 37884 32824 37890 32836
rect 39022 32824 39028 32836
rect 37884 32796 39028 32824
rect 37884 32784 37890 32796
rect 39022 32784 39028 32796
rect 39080 32784 39086 32836
rect 38197 32759 38255 32765
rect 38197 32756 38209 32759
rect 37752 32728 38209 32756
rect 38197 32725 38209 32728
rect 38243 32756 38255 32759
rect 38562 32756 38568 32768
rect 38243 32728 38568 32756
rect 38243 32725 38255 32728
rect 38197 32719 38255 32725
rect 38562 32716 38568 32728
rect 38620 32716 38626 32768
rect 1104 32666 58880 32688
rect 1104 32614 4874 32666
rect 4926 32614 4938 32666
rect 4990 32614 5002 32666
rect 5054 32614 5066 32666
rect 5118 32614 5130 32666
rect 5182 32614 35594 32666
rect 35646 32614 35658 32666
rect 35710 32614 35722 32666
rect 35774 32614 35786 32666
rect 35838 32614 35850 32666
rect 35902 32614 58880 32666
rect 1104 32592 58880 32614
rect 14642 32512 14648 32564
rect 14700 32552 14706 32564
rect 15933 32555 15991 32561
rect 15933 32552 15945 32555
rect 14700 32524 15945 32552
rect 14700 32512 14706 32524
rect 15933 32521 15945 32524
rect 15979 32521 15991 32555
rect 15933 32515 15991 32521
rect 26786 32512 26792 32564
rect 26844 32552 26850 32564
rect 27246 32552 27252 32564
rect 26844 32524 27252 32552
rect 26844 32512 26850 32524
rect 27246 32512 27252 32524
rect 27304 32512 27310 32564
rect 27341 32555 27399 32561
rect 27341 32521 27353 32555
rect 27387 32552 27399 32555
rect 27522 32552 27528 32564
rect 27387 32524 27528 32552
rect 27387 32521 27399 32524
rect 27341 32515 27399 32521
rect 27522 32512 27528 32524
rect 27580 32512 27586 32564
rect 30466 32512 30472 32564
rect 30524 32552 30530 32564
rect 34238 32552 34244 32564
rect 30524 32524 31754 32552
rect 30524 32512 30530 32524
rect 13906 32444 13912 32496
rect 13964 32484 13970 32496
rect 30834 32484 30840 32496
rect 13964 32456 16804 32484
rect 13964 32444 13970 32456
rect 16298 32376 16304 32428
rect 16356 32376 16362 32428
rect 16776 32425 16804 32456
rect 30116 32456 30840 32484
rect 16761 32419 16819 32425
rect 16761 32385 16773 32419
rect 16807 32416 16819 32419
rect 17310 32416 17316 32428
rect 16807 32388 17316 32416
rect 16807 32385 16819 32388
rect 16761 32379 16819 32385
rect 17310 32376 17316 32388
rect 17368 32376 17374 32428
rect 26326 32376 26332 32428
rect 26384 32416 26390 32428
rect 26421 32419 26479 32425
rect 26421 32416 26433 32419
rect 26384 32388 26433 32416
rect 26384 32376 26390 32388
rect 26421 32385 26433 32388
rect 26467 32385 26479 32419
rect 26973 32419 27031 32425
rect 26973 32416 26985 32419
rect 26421 32379 26479 32385
rect 26804 32388 26985 32416
rect 16393 32351 16451 32357
rect 16393 32317 16405 32351
rect 16439 32348 16451 32351
rect 17034 32348 17040 32360
rect 16439 32320 17040 32348
rect 16439 32317 16451 32320
rect 16393 32311 16451 32317
rect 17034 32308 17040 32320
rect 17092 32308 17098 32360
rect 26510 32308 26516 32360
rect 26568 32308 26574 32360
rect 26804 32357 26832 32388
rect 26973 32385 26985 32388
rect 27019 32385 27031 32419
rect 26973 32379 27031 32385
rect 27154 32376 27160 32428
rect 27212 32376 27218 32428
rect 30116 32425 30144 32456
rect 30834 32444 30840 32456
rect 30892 32444 30898 32496
rect 30101 32419 30159 32425
rect 30101 32385 30113 32419
rect 30147 32385 30159 32419
rect 30101 32379 30159 32385
rect 30466 32376 30472 32428
rect 30524 32376 30530 32428
rect 30558 32376 30564 32428
rect 30616 32416 30622 32428
rect 30653 32419 30711 32425
rect 30653 32416 30665 32419
rect 30616 32388 30665 32416
rect 30616 32376 30622 32388
rect 30653 32385 30665 32388
rect 30699 32385 30711 32419
rect 30653 32379 30711 32385
rect 26789 32351 26847 32357
rect 26789 32317 26801 32351
rect 26835 32317 26847 32351
rect 26789 32311 26847 32317
rect 30377 32351 30435 32357
rect 30377 32317 30389 32351
rect 30423 32348 30435 32351
rect 31294 32348 31300 32360
rect 30423 32320 31300 32348
rect 30423 32317 30435 32320
rect 30377 32311 30435 32317
rect 31294 32308 31300 32320
rect 31352 32308 31358 32360
rect 31726 32348 31754 32524
rect 33248 32524 34244 32552
rect 32950 32444 32956 32496
rect 33008 32484 33014 32496
rect 33137 32487 33195 32493
rect 33137 32484 33149 32487
rect 33008 32456 33149 32484
rect 33008 32444 33014 32456
rect 33137 32453 33149 32456
rect 33183 32484 33195 32487
rect 33248 32484 33276 32524
rect 34238 32512 34244 32524
rect 34296 32552 34302 32564
rect 34777 32555 34835 32561
rect 34296 32524 34652 32552
rect 34296 32512 34302 32524
rect 33183 32456 33276 32484
rect 33183 32453 33195 32456
rect 33137 32447 33195 32453
rect 33367 32453 33425 32459
rect 32858 32376 32864 32428
rect 32916 32416 32922 32428
rect 33367 32419 33379 32453
rect 33413 32419 33425 32453
rect 33778 32444 33784 32496
rect 33836 32484 33842 32496
rect 33873 32487 33931 32493
rect 33873 32484 33885 32487
rect 33836 32456 33885 32484
rect 33836 32444 33842 32456
rect 33873 32453 33885 32456
rect 33919 32453 33931 32487
rect 33873 32447 33931 32453
rect 34057 32487 34115 32493
rect 34057 32453 34069 32487
rect 34103 32484 34115 32487
rect 34146 32484 34152 32496
rect 34103 32456 34152 32484
rect 34103 32453 34115 32456
rect 34057 32447 34115 32453
rect 34146 32444 34152 32456
rect 34204 32444 34210 32496
rect 34517 32487 34575 32493
rect 34287 32453 34345 32459
rect 34287 32450 34299 32453
rect 33367 32416 33425 32419
rect 34275 32419 34299 32450
rect 34333 32428 34345 32453
rect 34517 32453 34529 32487
rect 34563 32453 34575 32487
rect 34624 32484 34652 32524
rect 34777 32521 34789 32555
rect 34823 32552 34835 32555
rect 35986 32552 35992 32564
rect 34823 32524 35992 32552
rect 34823 32521 34835 32524
rect 34777 32515 34835 32521
rect 35986 32512 35992 32524
rect 36044 32512 36050 32564
rect 36078 32512 36084 32564
rect 36136 32512 36142 32564
rect 36630 32552 36636 32564
rect 36464 32524 36636 32552
rect 34977 32487 35035 32493
rect 34977 32484 34989 32487
rect 34624 32456 34989 32484
rect 34517 32447 34575 32453
rect 34977 32453 34989 32456
rect 35023 32484 35035 32487
rect 35434 32484 35440 32496
rect 35023 32456 35440 32484
rect 35023 32453 35035 32456
rect 34977 32447 35035 32453
rect 34333 32419 34336 32428
rect 34275 32416 34336 32419
rect 32916 32388 34336 32416
rect 32916 32376 32922 32388
rect 34330 32376 34336 32388
rect 34388 32376 34394 32428
rect 34422 32376 34428 32428
rect 34480 32416 34486 32428
rect 34532 32416 34560 32447
rect 35434 32444 35440 32456
rect 35492 32444 35498 32496
rect 34480 32388 34836 32416
rect 34480 32376 34486 32388
rect 34514 32348 34520 32360
rect 31726 32320 34520 32348
rect 34514 32308 34520 32320
rect 34572 32348 34578 32360
rect 34808 32348 34836 32388
rect 34882 32376 34888 32428
rect 34940 32416 34946 32428
rect 35069 32419 35127 32425
rect 35069 32416 35081 32419
rect 34940 32388 35081 32416
rect 34940 32376 34946 32388
rect 35069 32385 35081 32388
rect 35115 32385 35127 32419
rect 35069 32379 35127 32385
rect 36262 32376 36268 32428
rect 36320 32376 36326 32428
rect 36464 32425 36492 32524
rect 36630 32512 36636 32524
rect 36688 32512 36694 32564
rect 37550 32484 37556 32496
rect 36556 32456 37556 32484
rect 36556 32425 36584 32456
rect 37550 32444 37556 32456
rect 37608 32444 37614 32496
rect 36449 32419 36507 32425
rect 36449 32385 36461 32419
rect 36495 32385 36507 32419
rect 36449 32379 36507 32385
rect 36541 32419 36599 32425
rect 36541 32385 36553 32419
rect 36587 32385 36599 32419
rect 36541 32379 36599 32385
rect 36817 32419 36875 32425
rect 36817 32385 36829 32419
rect 36863 32385 36875 32419
rect 36817 32379 36875 32385
rect 37001 32419 37059 32425
rect 37001 32385 37013 32419
rect 37047 32416 37059 32419
rect 37826 32416 37832 32428
rect 37047 32388 37832 32416
rect 37047 32385 37059 32388
rect 37001 32379 37059 32385
rect 36556 32348 36584 32379
rect 34572 32320 34652 32348
rect 34572 32308 34578 32320
rect 29362 32240 29368 32292
rect 29420 32280 29426 32292
rect 30469 32283 30527 32289
rect 30469 32280 30481 32283
rect 29420 32252 30481 32280
rect 29420 32240 29426 32252
rect 30469 32249 30481 32252
rect 30515 32249 30527 32283
rect 30469 32243 30527 32249
rect 33042 32240 33048 32292
rect 33100 32280 33106 32292
rect 34624 32289 34652 32320
rect 34808 32320 36584 32348
rect 33505 32283 33563 32289
rect 33505 32280 33517 32283
rect 33100 32252 33517 32280
rect 33100 32240 33106 32252
rect 33505 32249 33517 32252
rect 33551 32249 33563 32283
rect 34149 32283 34207 32289
rect 34149 32280 34161 32283
rect 33505 32243 33563 32249
rect 34072 32252 34161 32280
rect 17954 32172 17960 32224
rect 18012 32212 18018 32224
rect 18322 32212 18328 32224
rect 18012 32184 18328 32212
rect 18012 32172 18018 32184
rect 18322 32172 18328 32184
rect 18380 32172 18386 32224
rect 29914 32172 29920 32224
rect 29972 32172 29978 32224
rect 30098 32172 30104 32224
rect 30156 32212 30162 32224
rect 30285 32215 30343 32221
rect 30285 32212 30297 32215
rect 30156 32184 30297 32212
rect 30156 32172 30162 32184
rect 30285 32181 30297 32184
rect 30331 32181 30343 32215
rect 30285 32175 30343 32181
rect 33318 32172 33324 32224
rect 33376 32172 33382 32224
rect 33594 32172 33600 32224
rect 33652 32212 33658 32224
rect 33689 32215 33747 32221
rect 33689 32212 33701 32215
rect 33652 32184 33701 32212
rect 33652 32172 33658 32184
rect 33689 32181 33701 32184
rect 33735 32181 33747 32215
rect 33689 32175 33747 32181
rect 33870 32172 33876 32224
rect 33928 32212 33934 32224
rect 34072 32212 34100 32252
rect 34149 32249 34161 32252
rect 34195 32249 34207 32283
rect 34149 32243 34207 32249
rect 34609 32283 34667 32289
rect 34609 32249 34621 32283
rect 34655 32249 34667 32283
rect 34609 32243 34667 32249
rect 33928 32184 34100 32212
rect 33928 32172 33934 32184
rect 34238 32172 34244 32224
rect 34296 32212 34302 32224
rect 34808 32221 34836 32320
rect 35986 32240 35992 32292
rect 36044 32280 36050 32292
rect 36722 32280 36728 32292
rect 36044 32252 36728 32280
rect 36044 32240 36050 32252
rect 36722 32240 36728 32252
rect 36780 32280 36786 32292
rect 36832 32280 36860 32379
rect 36780 32252 36860 32280
rect 36780 32240 36786 32252
rect 34333 32215 34391 32221
rect 34333 32212 34345 32215
rect 34296 32184 34345 32212
rect 34296 32172 34302 32184
rect 34333 32181 34345 32184
rect 34379 32181 34391 32215
rect 34333 32175 34391 32181
rect 34793 32215 34851 32221
rect 34793 32181 34805 32215
rect 34839 32181 34851 32215
rect 34793 32175 34851 32181
rect 35434 32172 35440 32224
rect 35492 32212 35498 32224
rect 37016 32212 37044 32379
rect 37826 32376 37832 32388
rect 37884 32376 37890 32428
rect 35492 32184 37044 32212
rect 35492 32172 35498 32184
rect 1104 32122 58880 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 58880 32122
rect 1104 32048 58880 32070
rect 16482 32008 16488 32020
rect 15304 31980 16488 32008
rect 15304 31813 15332 31980
rect 16482 31968 16488 31980
rect 16540 32008 16546 32020
rect 18138 32008 18144 32020
rect 16540 31980 18144 32008
rect 16540 31968 16546 31980
rect 18138 31968 18144 31980
rect 18196 31968 18202 32020
rect 19426 31968 19432 32020
rect 19484 31968 19490 32020
rect 22094 31968 22100 32020
rect 22152 31968 22158 32020
rect 24578 31968 24584 32020
rect 24636 32008 24642 32020
rect 28902 32008 28908 32020
rect 24636 31980 28908 32008
rect 24636 31968 24642 31980
rect 28902 31968 28908 31980
rect 28960 31968 28966 32020
rect 29812 32011 29870 32017
rect 29812 31977 29824 32011
rect 29858 32008 29870 32011
rect 29914 32008 29920 32020
rect 29858 31980 29920 32008
rect 29858 31977 29870 31980
rect 29812 31971 29870 31977
rect 29914 31968 29920 31980
rect 29972 31968 29978 32020
rect 31294 31968 31300 32020
rect 31352 31968 31358 32020
rect 33778 31968 33784 32020
rect 33836 31968 33842 32020
rect 34149 32011 34207 32017
rect 34149 32008 34161 32011
rect 33888 31980 34161 32008
rect 15565 31943 15623 31949
rect 15565 31909 15577 31943
rect 15611 31940 15623 31943
rect 22112 31940 22140 31968
rect 15611 31912 17540 31940
rect 15611 31909 15623 31912
rect 15565 31903 15623 31909
rect 17512 31881 17540 31912
rect 22066 31912 22140 31940
rect 26053 31943 26111 31949
rect 17497 31875 17555 31881
rect 17497 31841 17509 31875
rect 17543 31841 17555 31875
rect 17497 31835 17555 31841
rect 18598 31832 18604 31884
rect 18656 31872 18662 31884
rect 19337 31875 19395 31881
rect 19337 31872 19349 31875
rect 18656 31844 19349 31872
rect 18656 31832 18662 31844
rect 19337 31841 19349 31844
rect 19383 31841 19395 31875
rect 19337 31835 19395 31841
rect 20257 31875 20315 31881
rect 20257 31841 20269 31875
rect 20303 31872 20315 31875
rect 20622 31872 20628 31884
rect 20303 31844 20628 31872
rect 20303 31841 20315 31844
rect 20257 31835 20315 31841
rect 20622 31832 20628 31844
rect 20680 31872 20686 31884
rect 22066 31872 22094 31912
rect 26053 31909 26065 31943
rect 26099 31940 26111 31943
rect 26099 31912 26372 31940
rect 26099 31909 26111 31912
rect 26053 31903 26111 31909
rect 20680 31844 22094 31872
rect 20680 31832 20686 31844
rect 15289 31807 15347 31813
rect 15289 31773 15301 31807
rect 15335 31773 15347 31807
rect 15289 31767 15347 31773
rect 15562 31764 15568 31816
rect 15620 31764 15626 31816
rect 15749 31807 15807 31813
rect 15749 31773 15761 31807
rect 15795 31804 15807 31807
rect 15838 31804 15844 31816
rect 15795 31776 15844 31804
rect 15795 31773 15807 31776
rect 15749 31767 15807 31773
rect 15381 31739 15439 31745
rect 15381 31705 15393 31739
rect 15427 31736 15439 31739
rect 15764 31736 15792 31767
rect 15838 31764 15844 31776
rect 15896 31764 15902 31816
rect 16393 31807 16451 31813
rect 16393 31773 16405 31807
rect 16439 31804 16451 31807
rect 17954 31804 17960 31816
rect 16439 31776 17960 31804
rect 16439 31773 16451 31776
rect 16393 31767 16451 31773
rect 17954 31764 17960 31776
rect 18012 31764 18018 31816
rect 18049 31807 18107 31813
rect 18049 31773 18061 31807
rect 18095 31804 18107 31807
rect 18141 31807 18199 31813
rect 18141 31804 18153 31807
rect 18095 31776 18153 31804
rect 18095 31773 18107 31776
rect 18049 31767 18107 31773
rect 18141 31773 18153 31776
rect 18187 31773 18199 31807
rect 18141 31767 18199 31773
rect 18325 31807 18383 31813
rect 18325 31773 18337 31807
rect 18371 31804 18383 31807
rect 18414 31804 18420 31816
rect 18371 31776 18420 31804
rect 18371 31773 18383 31776
rect 18325 31767 18383 31773
rect 18414 31764 18420 31776
rect 18472 31764 18478 31816
rect 19242 31764 19248 31816
rect 19300 31764 19306 31816
rect 22066 31813 22094 31844
rect 23658 31832 23664 31884
rect 23716 31872 23722 31884
rect 23845 31875 23903 31881
rect 23845 31872 23857 31875
rect 23716 31844 23857 31872
rect 23716 31832 23722 31844
rect 23845 31841 23857 31844
rect 23891 31872 23903 31875
rect 24949 31875 25007 31881
rect 24949 31872 24961 31875
rect 23891 31844 24961 31872
rect 23891 31841 23903 31844
rect 23845 31835 23903 31841
rect 24949 31841 24961 31844
rect 24995 31841 25007 31875
rect 24949 31835 25007 31841
rect 25590 31832 25596 31884
rect 25648 31872 25654 31884
rect 25648 31844 26188 31872
rect 25648 31832 25654 31844
rect 19521 31807 19579 31813
rect 19521 31773 19533 31807
rect 19567 31773 19579 31807
rect 22066 31807 22144 31813
rect 22066 31776 22098 31807
rect 19521 31767 19579 31773
rect 22086 31773 22098 31776
rect 22132 31773 22144 31807
rect 22086 31767 22144 31773
rect 15427 31708 15792 31736
rect 17221 31739 17279 31745
rect 15427 31705 15439 31708
rect 15381 31699 15439 31705
rect 17221 31705 17233 31739
rect 17267 31736 17279 31739
rect 17310 31736 17316 31748
rect 17267 31708 17316 31736
rect 17267 31705 17279 31708
rect 17221 31699 17279 31705
rect 17310 31696 17316 31708
rect 17368 31696 17374 31748
rect 19536 31736 19564 31767
rect 25406 31764 25412 31816
rect 25464 31764 25470 31816
rect 26160 31813 26188 31844
rect 26145 31807 26203 31813
rect 26145 31773 26157 31807
rect 26191 31773 26203 31807
rect 26145 31767 26203 31773
rect 26234 31764 26240 31816
rect 26292 31764 26298 31816
rect 26344 31813 26372 31912
rect 26329 31807 26387 31813
rect 26329 31773 26341 31807
rect 26375 31773 26387 31807
rect 28920 31804 28948 31968
rect 31312 31940 31340 31968
rect 33502 31940 33508 31952
rect 31312 31912 33508 31940
rect 28994 31832 29000 31884
rect 29052 31872 29058 31884
rect 29549 31875 29607 31881
rect 29549 31872 29561 31875
rect 29052 31844 29561 31872
rect 29052 31832 29058 31844
rect 29549 31841 29561 31844
rect 29595 31872 29607 31875
rect 29595 31844 31064 31872
rect 29595 31841 29607 31844
rect 29549 31835 29607 31841
rect 29089 31807 29147 31813
rect 29089 31804 29101 31807
rect 28920 31776 29101 31804
rect 26329 31767 26387 31773
rect 29089 31773 29101 31776
rect 29135 31773 29147 31807
rect 29273 31807 29331 31813
rect 29273 31804 29285 31807
rect 29251 31776 29285 31804
rect 29089 31767 29147 31773
rect 29273 31773 29285 31776
rect 29319 31773 29331 31807
rect 29273 31767 29331 31773
rect 19536 31708 20484 31736
rect 16114 31628 16120 31680
rect 16172 31668 16178 31680
rect 16301 31671 16359 31677
rect 16301 31668 16313 31671
rect 16172 31640 16313 31668
rect 16172 31628 16178 31640
rect 16301 31637 16313 31640
rect 16347 31637 16359 31671
rect 16301 31631 16359 31637
rect 18230 31628 18236 31680
rect 18288 31628 18294 31680
rect 19702 31628 19708 31680
rect 19760 31628 19766 31680
rect 20456 31668 20484 31708
rect 20530 31696 20536 31748
rect 20588 31696 20594 31748
rect 22278 31736 22284 31748
rect 21758 31708 22284 31736
rect 22278 31696 22284 31708
rect 22336 31696 22342 31748
rect 22370 31696 22376 31748
rect 22428 31696 22434 31748
rect 23750 31736 23756 31748
rect 23598 31708 23756 31736
rect 23750 31696 23756 31708
rect 23808 31696 23814 31748
rect 29288 31736 29316 31767
rect 29362 31764 29368 31816
rect 29420 31764 29426 31816
rect 31036 31804 31064 31844
rect 33244 31816 33272 31912
rect 33502 31900 33508 31912
rect 33560 31900 33566 31952
rect 33594 31900 33600 31952
rect 33652 31940 33658 31952
rect 33888 31940 33916 31980
rect 34149 31977 34161 31980
rect 34195 31977 34207 32011
rect 34149 31971 34207 31977
rect 37366 31968 37372 32020
rect 37424 32008 37430 32020
rect 37461 32011 37519 32017
rect 37461 32008 37473 32011
rect 37424 31980 37473 32008
rect 37424 31968 37430 31980
rect 37461 31977 37473 31980
rect 37507 32008 37519 32011
rect 37550 32008 37556 32020
rect 37507 31980 37556 32008
rect 37507 31977 37519 31980
rect 37461 31971 37519 31977
rect 37550 31968 37556 31980
rect 37608 31968 37614 32020
rect 34238 31940 34244 31952
rect 33652 31912 33916 31940
rect 33996 31912 34244 31940
rect 33652 31900 33658 31912
rect 33520 31872 33548 31900
rect 33996 31872 34024 31912
rect 34238 31900 34244 31912
rect 34296 31900 34302 31952
rect 36722 31900 36728 31952
rect 36780 31940 36786 31952
rect 37093 31943 37151 31949
rect 37093 31940 37105 31943
rect 36780 31912 37105 31940
rect 36780 31900 36786 31912
rect 37093 31909 37105 31912
rect 37139 31909 37151 31943
rect 37093 31903 37151 31909
rect 37645 31943 37703 31949
rect 37645 31909 37657 31943
rect 37691 31940 37703 31943
rect 38746 31940 38752 31952
rect 37691 31912 38752 31940
rect 37691 31909 37703 31912
rect 37645 31903 37703 31909
rect 38746 31900 38752 31912
rect 38804 31900 38810 31952
rect 33520 31844 34024 31872
rect 34790 31832 34796 31884
rect 34848 31872 34854 31884
rect 38378 31872 38384 31884
rect 34848 31844 38384 31872
rect 34848 31832 34854 31844
rect 38378 31832 38384 31844
rect 38436 31832 38442 31884
rect 32306 31804 32312 31816
rect 31036 31776 32312 31804
rect 32306 31764 32312 31776
rect 32364 31764 32370 31816
rect 32950 31764 32956 31816
rect 33008 31804 33014 31816
rect 33045 31807 33103 31813
rect 33045 31804 33057 31807
rect 33008 31776 33057 31804
rect 33008 31764 33014 31776
rect 33045 31773 33057 31776
rect 33091 31773 33103 31807
rect 33045 31767 33103 31773
rect 33137 31785 33195 31791
rect 33137 31751 33149 31785
rect 33183 31751 33195 31785
rect 33226 31764 33232 31816
rect 33284 31764 33290 31816
rect 33410 31764 33416 31816
rect 33468 31804 33474 31816
rect 33597 31807 33655 31813
rect 33597 31804 33609 31807
rect 33468 31776 33609 31804
rect 33468 31764 33474 31776
rect 33597 31773 33609 31776
rect 33643 31773 33655 31807
rect 33597 31767 33655 31773
rect 33781 31807 33839 31813
rect 33781 31773 33793 31807
rect 33827 31804 33839 31807
rect 33870 31804 33876 31816
rect 33827 31776 33876 31804
rect 33827 31773 33839 31776
rect 33781 31767 33839 31773
rect 33870 31764 33876 31776
rect 33928 31764 33934 31816
rect 33962 31764 33968 31816
rect 34020 31804 34026 31816
rect 34149 31807 34207 31813
rect 34149 31804 34161 31807
rect 34020 31776 34161 31804
rect 34020 31764 34026 31776
rect 34149 31773 34161 31776
rect 34195 31773 34207 31807
rect 34149 31767 34207 31773
rect 34241 31807 34299 31813
rect 34241 31773 34253 31807
rect 34287 31804 34299 31807
rect 34698 31804 34704 31816
rect 34287 31776 34704 31804
rect 34287 31773 34299 31776
rect 34241 31767 34299 31773
rect 34698 31764 34704 31776
rect 34756 31764 34762 31816
rect 37826 31764 37832 31816
rect 37884 31804 37890 31816
rect 38105 31807 38163 31813
rect 38105 31804 38117 31807
rect 37884 31776 38117 31804
rect 37884 31764 37890 31776
rect 38105 31773 38117 31776
rect 38151 31773 38163 31807
rect 38105 31767 38163 31773
rect 30098 31736 30104 31748
rect 29288 31708 30104 31736
rect 30098 31696 30104 31708
rect 30156 31696 30162 31748
rect 31570 31736 31576 31748
rect 31050 31708 31576 31736
rect 31570 31696 31576 31708
rect 31628 31696 31634 31748
rect 33137 31745 33195 31751
rect 21450 31668 21456 31680
rect 20456 31640 21456 31668
rect 21450 31628 21456 31640
rect 21508 31668 21514 31680
rect 22005 31671 22063 31677
rect 22005 31668 22017 31671
rect 21508 31640 22017 31668
rect 21508 31628 21514 31640
rect 22005 31637 22017 31640
rect 22051 31668 22063 31671
rect 22554 31668 22560 31680
rect 22051 31640 22560 31668
rect 22051 31637 22063 31640
rect 22005 31631 22063 31637
rect 22554 31628 22560 31640
rect 22612 31628 22618 31680
rect 24394 31628 24400 31680
rect 24452 31628 24458 31680
rect 29362 31628 29368 31680
rect 29420 31628 29426 31680
rect 30558 31628 30564 31680
rect 30616 31668 30622 31680
rect 32858 31668 32864 31680
rect 30616 31640 32864 31668
rect 30616 31628 30622 31640
rect 32858 31628 32864 31640
rect 32916 31668 32922 31680
rect 33152 31668 33180 31745
rect 33318 31696 33324 31748
rect 33376 31736 33382 31748
rect 34425 31739 34483 31745
rect 33376 31708 34100 31736
rect 33376 31696 33382 31708
rect 32916 31640 33180 31668
rect 32916 31628 32922 31640
rect 33502 31628 33508 31680
rect 33560 31628 33566 31680
rect 33686 31628 33692 31680
rect 33744 31668 33750 31680
rect 33965 31671 34023 31677
rect 33965 31668 33977 31671
rect 33744 31640 33977 31668
rect 33744 31628 33750 31640
rect 33965 31637 33977 31640
rect 34011 31637 34023 31671
rect 34072 31668 34100 31708
rect 34425 31705 34437 31739
rect 34471 31736 34483 31739
rect 34606 31736 34612 31748
rect 34471 31708 34612 31736
rect 34471 31705 34483 31708
rect 34425 31699 34483 31705
rect 34606 31696 34612 31708
rect 34664 31696 34670 31748
rect 37918 31696 37924 31748
rect 37976 31696 37982 31748
rect 34514 31668 34520 31680
rect 34072 31640 34520 31668
rect 33965 31631 34023 31637
rect 34514 31628 34520 31640
rect 34572 31628 34578 31680
rect 37461 31671 37519 31677
rect 37461 31637 37473 31671
rect 37507 31668 37519 31671
rect 37737 31671 37795 31677
rect 37737 31668 37749 31671
rect 37507 31640 37749 31668
rect 37507 31637 37519 31640
rect 37461 31631 37519 31637
rect 37737 31637 37749 31640
rect 37783 31637 37795 31671
rect 37737 31631 37795 31637
rect 1104 31578 58880 31600
rect 1104 31526 4874 31578
rect 4926 31526 4938 31578
rect 4990 31526 5002 31578
rect 5054 31526 5066 31578
rect 5118 31526 5130 31578
rect 5182 31526 35594 31578
rect 35646 31526 35658 31578
rect 35710 31526 35722 31578
rect 35774 31526 35786 31578
rect 35838 31526 35850 31578
rect 35902 31526 58880 31578
rect 1104 31504 58880 31526
rect 15562 31424 15568 31476
rect 15620 31464 15626 31476
rect 16669 31467 16727 31473
rect 16669 31464 16681 31467
rect 15620 31436 16681 31464
rect 15620 31424 15626 31436
rect 16669 31433 16681 31436
rect 16715 31433 16727 31467
rect 16669 31427 16727 31433
rect 18138 31424 18144 31476
rect 18196 31473 18202 31476
rect 18196 31467 18215 31473
rect 18203 31433 18215 31467
rect 18196 31427 18215 31433
rect 18325 31467 18383 31473
rect 18325 31433 18337 31467
rect 18371 31464 18383 31467
rect 18414 31464 18420 31476
rect 18371 31436 18420 31464
rect 18371 31433 18383 31436
rect 18325 31427 18383 31433
rect 18196 31424 18202 31427
rect 18414 31424 18420 31436
rect 18472 31424 18478 31476
rect 21913 31467 21971 31473
rect 21913 31433 21925 31467
rect 21959 31464 21971 31467
rect 22370 31464 22376 31476
rect 21959 31436 22376 31464
rect 21959 31433 21971 31436
rect 21913 31427 21971 31433
rect 22370 31424 22376 31436
rect 22428 31424 22434 31476
rect 23842 31424 23848 31476
rect 23900 31424 23906 31476
rect 24765 31467 24823 31473
rect 24765 31464 24777 31467
rect 24504 31436 24777 31464
rect 15930 31396 15936 31408
rect 15410 31368 15936 31396
rect 15930 31356 15936 31368
rect 15988 31356 15994 31408
rect 17773 31399 17831 31405
rect 17773 31365 17785 31399
rect 17819 31396 17831 31399
rect 17862 31396 17868 31408
rect 17819 31368 17868 31396
rect 17819 31365 17831 31368
rect 17773 31359 17831 31365
rect 17862 31356 17868 31368
rect 17920 31356 17926 31408
rect 17957 31399 18015 31405
rect 17957 31365 17969 31399
rect 18003 31365 18015 31399
rect 17957 31359 18015 31365
rect 18432 31396 18460 31424
rect 22278 31405 22284 31408
rect 22265 31399 22284 31405
rect 18432 31368 19012 31396
rect 13906 31288 13912 31340
rect 13964 31288 13970 31340
rect 16114 31288 16120 31340
rect 16172 31288 16178 31340
rect 14185 31263 14243 31269
rect 14185 31229 14197 31263
rect 14231 31260 14243 31263
rect 15749 31263 15807 31269
rect 15749 31260 15761 31263
rect 14231 31232 15761 31260
rect 14231 31229 14243 31232
rect 14185 31223 14243 31229
rect 15749 31229 15761 31232
rect 15795 31229 15807 31263
rect 15749 31223 15807 31229
rect 16209 31263 16267 31269
rect 16209 31229 16221 31263
rect 16255 31260 16267 31263
rect 16482 31260 16488 31272
rect 16255 31232 16488 31260
rect 16255 31229 16267 31232
rect 16209 31223 16267 31229
rect 16482 31220 16488 31232
rect 16540 31220 16546 31272
rect 17218 31220 17224 31272
rect 17276 31260 17282 31272
rect 17972 31260 18000 31359
rect 18432 31328 18460 31368
rect 18984 31337 19012 31368
rect 22265 31365 22277 31399
rect 22265 31359 22284 31365
rect 22278 31356 22284 31359
rect 22336 31356 22342 31408
rect 22465 31399 22523 31405
rect 22465 31365 22477 31399
rect 22511 31396 22523 31399
rect 22554 31396 22560 31408
rect 22511 31368 22560 31396
rect 22511 31365 22523 31368
rect 22465 31359 22523 31365
rect 22554 31356 22560 31368
rect 22612 31396 22618 31408
rect 22612 31368 22692 31396
rect 22612 31356 22618 31368
rect 18509 31331 18567 31337
rect 18509 31328 18521 31331
rect 18432 31300 18521 31328
rect 18509 31297 18521 31300
rect 18555 31297 18567 31331
rect 18705 31331 18763 31337
rect 18705 31326 18717 31331
rect 18509 31291 18567 31297
rect 18616 31298 18717 31326
rect 17276 31232 18000 31260
rect 17276 31220 17282 31232
rect 15657 31195 15715 31201
rect 15657 31161 15669 31195
rect 15703 31192 15715 31195
rect 15838 31192 15844 31204
rect 15703 31164 15844 31192
rect 15703 31161 15715 31164
rect 15657 31155 15715 31161
rect 15838 31152 15844 31164
rect 15896 31192 15902 31204
rect 15896 31164 17816 31192
rect 15896 31152 15902 31164
rect 17788 31136 17816 31164
rect 15930 31084 15936 31136
rect 15988 31124 15994 31136
rect 16482 31124 16488 31136
rect 15988 31096 16488 31124
rect 15988 31084 15994 31096
rect 16482 31084 16488 31096
rect 16540 31124 16546 31136
rect 17497 31127 17555 31133
rect 17497 31124 17509 31127
rect 16540 31096 17509 31124
rect 16540 31084 16546 31096
rect 17497 31093 17509 31096
rect 17543 31093 17555 31127
rect 17497 31087 17555 31093
rect 17770 31084 17776 31136
rect 17828 31124 17834 31136
rect 18141 31127 18199 31133
rect 18141 31124 18153 31127
rect 17828 31096 18153 31124
rect 17828 31084 17834 31096
rect 18141 31093 18153 31096
rect 18187 31093 18199 31127
rect 18141 31087 18199 31093
rect 18506 31084 18512 31136
rect 18564 31084 18570 31136
rect 18616 31124 18644 31298
rect 18705 31297 18717 31298
rect 18751 31297 18763 31331
rect 18705 31291 18763 31297
rect 18969 31331 19027 31337
rect 18969 31297 18981 31331
rect 19015 31297 19027 31331
rect 18969 31291 19027 31297
rect 20165 31331 20223 31337
rect 20165 31297 20177 31331
rect 20211 31328 20223 31331
rect 20901 31331 20959 31337
rect 20901 31328 20913 31331
rect 20211 31300 20913 31328
rect 20211 31297 20223 31300
rect 20165 31291 20223 31297
rect 20901 31297 20913 31300
rect 20947 31297 20959 31331
rect 20901 31291 20959 31297
rect 21450 31288 21456 31340
rect 21508 31288 21514 31340
rect 21821 31331 21879 31337
rect 21821 31297 21833 31331
rect 21867 31297 21879 31331
rect 21821 31291 21879 31297
rect 18785 31263 18843 31269
rect 18785 31229 18797 31263
rect 18831 31260 18843 31263
rect 19426 31260 19432 31272
rect 18831 31232 19432 31260
rect 18831 31229 18843 31232
rect 18785 31223 18843 31229
rect 19426 31220 19432 31232
rect 19484 31260 19490 31272
rect 19794 31260 19800 31272
rect 19484 31232 19800 31260
rect 19484 31220 19490 31232
rect 19794 31220 19800 31232
rect 19852 31220 19858 31272
rect 20257 31263 20315 31269
rect 20257 31229 20269 31263
rect 20303 31229 20315 31263
rect 20257 31223 20315 31229
rect 19153 31195 19211 31201
rect 19153 31161 19165 31195
rect 19199 31192 19211 31195
rect 20272 31192 20300 31223
rect 20530 31220 20536 31272
rect 20588 31220 20594 31272
rect 21836 31260 21864 31291
rect 22002 31288 22008 31340
rect 22060 31288 22066 31340
rect 22664 31337 22692 31368
rect 23382 31356 23388 31408
rect 23440 31356 23446 31408
rect 22649 31331 22707 31337
rect 22649 31297 22661 31331
rect 22695 31297 22707 31331
rect 22649 31291 22707 31297
rect 23661 31331 23719 31337
rect 23661 31297 23673 31331
rect 23707 31328 23719 31331
rect 24504 31328 24532 31436
rect 24765 31433 24777 31436
rect 24811 31464 24823 31467
rect 24854 31464 24860 31476
rect 24811 31436 24860 31464
rect 24811 31433 24823 31436
rect 24765 31427 24823 31433
rect 24854 31424 24860 31436
rect 24912 31424 24918 31476
rect 27430 31424 27436 31476
rect 27488 31464 27494 31476
rect 27488 31436 29132 31464
rect 27488 31424 27494 31436
rect 28994 31396 29000 31408
rect 28460 31368 29000 31396
rect 23707 31300 24532 31328
rect 23707 31297 23719 31300
rect 23661 31291 23719 31297
rect 24670 31288 24676 31340
rect 24728 31288 24734 31340
rect 24949 31331 25007 31337
rect 24949 31297 24961 31331
rect 24995 31328 25007 31331
rect 25041 31331 25099 31337
rect 25041 31328 25053 31331
rect 24995 31300 25053 31328
rect 24995 31297 25007 31300
rect 24949 31291 25007 31297
rect 25041 31297 25053 31300
rect 25087 31297 25099 31331
rect 25041 31291 25099 31297
rect 25682 31288 25688 31340
rect 25740 31328 25746 31340
rect 28460 31337 28488 31368
rect 28994 31356 29000 31368
rect 29052 31356 29058 31408
rect 29104 31396 29132 31436
rect 29546 31424 29552 31476
rect 29604 31464 29610 31476
rect 30190 31464 30196 31476
rect 29604 31436 30196 31464
rect 29604 31424 29610 31436
rect 30190 31424 30196 31436
rect 30248 31464 30254 31476
rect 30469 31467 30527 31473
rect 30469 31464 30481 31467
rect 30248 31436 30481 31464
rect 30248 31424 30254 31436
rect 30469 31433 30481 31436
rect 30515 31433 30527 31467
rect 30469 31427 30527 31433
rect 30484 31396 30512 31427
rect 36722 31424 36728 31476
rect 36780 31424 36786 31476
rect 37277 31467 37335 31473
rect 37277 31433 37289 31467
rect 37323 31464 37335 31467
rect 37918 31464 37924 31476
rect 37323 31436 37924 31464
rect 37323 31433 37335 31436
rect 37277 31427 37335 31433
rect 30653 31399 30711 31405
rect 30653 31396 30665 31399
rect 29104 31368 29210 31396
rect 30484 31368 30665 31396
rect 30653 31365 30665 31368
rect 30699 31365 30711 31399
rect 30653 31359 30711 31365
rect 31481 31399 31539 31405
rect 31481 31365 31493 31399
rect 31527 31396 31539 31399
rect 32030 31396 32036 31408
rect 31527 31368 32036 31396
rect 31527 31365 31539 31368
rect 31481 31359 31539 31365
rect 32030 31356 32036 31368
rect 32088 31396 32094 31408
rect 32306 31396 32312 31408
rect 32088 31368 32312 31396
rect 32088 31356 32094 31368
rect 32306 31356 32312 31368
rect 32364 31356 32370 31408
rect 36630 31356 36636 31408
rect 36688 31396 36694 31408
rect 36877 31399 36935 31405
rect 36877 31396 36889 31399
rect 36688 31368 36889 31396
rect 36688 31356 36694 31368
rect 36877 31365 36889 31368
rect 36923 31365 36935 31399
rect 36877 31359 36935 31365
rect 37093 31399 37151 31405
rect 37093 31365 37105 31399
rect 37139 31396 37151 31399
rect 37292 31396 37320 31427
rect 37918 31424 37924 31436
rect 37976 31424 37982 31476
rect 38654 31396 38660 31408
rect 37139 31368 37320 31396
rect 38318 31368 38660 31396
rect 37139 31365 37151 31368
rect 37093 31359 37151 31365
rect 26513 31331 26571 31337
rect 26513 31328 26525 31331
rect 25740 31300 26525 31328
rect 25740 31288 25746 31300
rect 26513 31297 26525 31300
rect 26559 31297 26571 31331
rect 26513 31291 26571 31297
rect 26697 31331 26755 31337
rect 26697 31297 26709 31331
rect 26743 31297 26755 31331
rect 26697 31291 26755 31297
rect 28445 31331 28503 31337
rect 28445 31297 28457 31331
rect 28491 31297 28503 31331
rect 28445 31291 28503 31297
rect 21744 31232 21864 31260
rect 23569 31263 23627 31269
rect 21634 31192 21640 31204
rect 19199 31164 21640 31192
rect 19199 31161 19211 31164
rect 19153 31155 19211 31161
rect 19444 31136 19472 31164
rect 21634 31152 21640 31164
rect 21692 31152 21698 31204
rect 19245 31127 19303 31133
rect 19245 31124 19257 31127
rect 18616 31096 19257 31124
rect 19245 31093 19257 31096
rect 19291 31093 19303 31127
rect 19245 31087 19303 31093
rect 19426 31084 19432 31136
rect 19484 31084 19490 31136
rect 21744 31124 21772 31232
rect 23569 31229 23581 31263
rect 23615 31260 23627 31263
rect 23615 31232 25544 31260
rect 23615 31229 23627 31232
rect 23569 31223 23627 31229
rect 21818 31152 21824 31204
rect 21876 31192 21882 31204
rect 22186 31192 22192 31204
rect 21876 31164 22192 31192
rect 21876 31152 21882 31164
rect 22186 31152 22192 31164
rect 22244 31152 22250 31204
rect 24949 31195 25007 31201
rect 22848 31164 23704 31192
rect 21910 31124 21916 31136
rect 21744 31096 21916 31124
rect 21910 31084 21916 31096
rect 21968 31124 21974 31136
rect 22097 31127 22155 31133
rect 22097 31124 22109 31127
rect 21968 31096 22109 31124
rect 21968 31084 21974 31096
rect 22097 31093 22109 31096
rect 22143 31093 22155 31127
rect 22097 31087 22155 31093
rect 22281 31127 22339 31133
rect 22281 31093 22293 31127
rect 22327 31124 22339 31127
rect 22848 31124 22876 31164
rect 23676 31136 23704 31164
rect 24949 31161 24961 31195
rect 24995 31192 25007 31195
rect 25406 31192 25412 31204
rect 24995 31164 25412 31192
rect 24995 31161 25007 31164
rect 24949 31155 25007 31161
rect 25406 31152 25412 31164
rect 25464 31152 25470 31204
rect 25516 31192 25544 31232
rect 26326 31220 26332 31272
rect 26384 31260 26390 31272
rect 26712 31260 26740 31291
rect 30374 31288 30380 31340
rect 30432 31328 30438 31340
rect 31570 31328 31576 31340
rect 30432 31300 31576 31328
rect 30432 31288 30438 31300
rect 31570 31288 31576 31300
rect 31628 31288 31634 31340
rect 33226 31288 33232 31340
rect 33284 31328 33290 31340
rect 33413 31331 33471 31337
rect 33413 31328 33425 31331
rect 33284 31300 33425 31328
rect 33284 31288 33290 31300
rect 33413 31297 33425 31300
rect 33459 31297 33471 31331
rect 33413 31291 33471 31297
rect 33505 31331 33563 31337
rect 33505 31297 33517 31331
rect 33551 31328 33563 31331
rect 33594 31328 33600 31340
rect 33551 31300 33600 31328
rect 33551 31297 33563 31300
rect 33505 31291 33563 31297
rect 33594 31288 33600 31300
rect 33652 31288 33658 31340
rect 33873 31331 33931 31337
rect 33873 31297 33885 31331
rect 33919 31328 33931 31331
rect 33962 31328 33968 31340
rect 33919 31300 33968 31328
rect 33919 31297 33931 31300
rect 33873 31291 33931 31297
rect 33962 31288 33968 31300
rect 34020 31288 34026 31340
rect 34330 31288 34336 31340
rect 34388 31288 34394 31340
rect 34698 31288 34704 31340
rect 34756 31328 34762 31340
rect 37108 31328 37136 31359
rect 38654 31356 38660 31368
rect 38712 31356 38718 31408
rect 38746 31356 38752 31408
rect 38804 31356 38810 31408
rect 34756 31300 37136 31328
rect 34756 31288 34762 31300
rect 26384 31232 26740 31260
rect 28721 31263 28779 31269
rect 26384 31220 26390 31232
rect 28721 31229 28733 31263
rect 28767 31260 28779 31263
rect 29362 31260 29368 31272
rect 28767 31232 29368 31260
rect 28767 31229 28779 31232
rect 28721 31223 28779 31229
rect 29362 31220 29368 31232
rect 29420 31220 29426 31272
rect 34241 31263 34299 31269
rect 34241 31229 34253 31263
rect 34287 31260 34299 31263
rect 34422 31260 34428 31272
rect 34287 31232 34428 31260
rect 34287 31229 34299 31232
rect 34241 31223 34299 31229
rect 34422 31220 34428 31232
rect 34480 31220 34486 31272
rect 36354 31220 36360 31272
rect 36412 31260 36418 31272
rect 36633 31263 36691 31269
rect 36633 31260 36645 31263
rect 36412 31232 36645 31260
rect 36412 31220 36418 31232
rect 36633 31229 36645 31232
rect 36679 31260 36691 31263
rect 38654 31260 38660 31272
rect 36679 31232 38660 31260
rect 36679 31229 36691 31232
rect 36633 31223 36691 31229
rect 38654 31220 38660 31232
rect 38712 31220 38718 31272
rect 39025 31263 39083 31269
rect 39025 31229 39037 31263
rect 39071 31229 39083 31263
rect 39025 31223 39083 31229
rect 26605 31195 26663 31201
rect 26605 31192 26617 31195
rect 25516 31164 26617 31192
rect 26605 31161 26617 31164
rect 26651 31161 26663 31195
rect 26605 31155 26663 31161
rect 22327 31096 22876 31124
rect 22327 31093 22339 31096
rect 22281 31087 22339 31093
rect 22922 31084 22928 31136
rect 22980 31124 22986 31136
rect 23201 31127 23259 31133
rect 23201 31124 23213 31127
rect 22980 31096 23213 31124
rect 22980 31084 22986 31096
rect 23201 31093 23213 31096
rect 23247 31093 23259 31127
rect 23201 31087 23259 31093
rect 23658 31084 23664 31136
rect 23716 31084 23722 31136
rect 25498 31084 25504 31136
rect 25556 31124 25562 31136
rect 25777 31127 25835 31133
rect 25777 31124 25789 31127
rect 25556 31096 25789 31124
rect 25556 31084 25562 31096
rect 25777 31093 25789 31096
rect 25823 31093 25835 31127
rect 25777 31087 25835 31093
rect 30193 31127 30251 31133
rect 30193 31093 30205 31127
rect 30239 31124 30251 31127
rect 30558 31124 30564 31136
rect 30239 31096 30564 31124
rect 30239 31093 30251 31096
rect 30193 31087 30251 31093
rect 30558 31084 30564 31096
rect 30616 31084 30622 31136
rect 32950 31084 32956 31136
rect 33008 31124 33014 31136
rect 33781 31127 33839 31133
rect 33781 31124 33793 31127
rect 33008 31096 33793 31124
rect 33008 31084 33014 31096
rect 33781 31093 33793 31096
rect 33827 31093 33839 31127
rect 33781 31087 33839 31093
rect 34054 31084 34060 31136
rect 34112 31084 34118 31136
rect 34606 31084 34612 31136
rect 34664 31084 34670 31136
rect 34698 31084 34704 31136
rect 34756 31124 34762 31136
rect 34885 31127 34943 31133
rect 34885 31124 34897 31127
rect 34756 31096 34897 31124
rect 34756 31084 34762 31096
rect 34885 31093 34897 31096
rect 34931 31093 34943 31127
rect 34885 31087 34943 31093
rect 36814 31084 36820 31136
rect 36872 31124 36878 31136
rect 36909 31127 36967 31133
rect 36909 31124 36921 31127
rect 36872 31096 36921 31124
rect 36872 31084 36878 31096
rect 36909 31093 36921 31096
rect 36955 31093 36967 31127
rect 36909 31087 36967 31093
rect 38746 31084 38752 31136
rect 38804 31124 38810 31136
rect 39040 31124 39068 31223
rect 38804 31096 39068 31124
rect 38804 31084 38810 31096
rect 1104 31034 58880 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 58880 31034
rect 1104 30960 58880 30982
rect 15565 30923 15623 30929
rect 15565 30889 15577 30923
rect 15611 30920 15623 30923
rect 17218 30920 17224 30932
rect 15611 30892 17224 30920
rect 15611 30889 15623 30892
rect 15565 30883 15623 30889
rect 17218 30880 17224 30892
rect 17276 30880 17282 30932
rect 17865 30923 17923 30929
rect 17865 30889 17877 30923
rect 17911 30920 17923 30923
rect 18598 30920 18604 30932
rect 17911 30892 18604 30920
rect 17911 30889 17923 30892
rect 17865 30883 17923 30889
rect 18598 30880 18604 30892
rect 18656 30880 18662 30932
rect 22002 30880 22008 30932
rect 22060 30920 22066 30932
rect 23109 30923 23167 30929
rect 23109 30920 23121 30923
rect 22060 30892 23121 30920
rect 22060 30880 22066 30892
rect 23109 30889 23121 30892
rect 23155 30889 23167 30923
rect 23109 30883 23167 30889
rect 25038 30880 25044 30932
rect 25096 30920 25102 30932
rect 25682 30920 25688 30932
rect 25096 30892 25688 30920
rect 25096 30880 25102 30892
rect 25682 30880 25688 30892
rect 25740 30880 25746 30932
rect 25961 30923 26019 30929
rect 25961 30889 25973 30923
rect 26007 30920 26019 30923
rect 26326 30920 26332 30932
rect 26007 30892 26332 30920
rect 26007 30889 26019 30892
rect 25961 30883 26019 30889
rect 26326 30880 26332 30892
rect 26384 30880 26390 30932
rect 30098 30880 30104 30932
rect 30156 30920 30162 30932
rect 30285 30923 30343 30929
rect 30285 30920 30297 30923
rect 30156 30892 30297 30920
rect 30156 30880 30162 30892
rect 30285 30889 30297 30892
rect 30331 30889 30343 30923
rect 30285 30883 30343 30889
rect 33597 30923 33655 30929
rect 33597 30889 33609 30923
rect 33643 30920 33655 30923
rect 33870 30920 33876 30932
rect 33643 30892 33876 30920
rect 33643 30889 33655 30892
rect 33597 30883 33655 30889
rect 33870 30880 33876 30892
rect 33928 30880 33934 30932
rect 34054 30880 34060 30932
rect 34112 30920 34118 30932
rect 34260 30923 34318 30929
rect 34260 30920 34272 30923
rect 34112 30892 34272 30920
rect 34112 30880 34118 30892
rect 34260 30889 34272 30892
rect 34306 30889 34318 30923
rect 34260 30883 34318 30889
rect 34790 30880 34796 30932
rect 34848 30920 34854 30932
rect 34885 30923 34943 30929
rect 34885 30920 34897 30923
rect 34848 30892 34897 30920
rect 34848 30880 34854 30892
rect 34885 30889 34897 30892
rect 34931 30889 34943 30923
rect 34885 30883 34943 30889
rect 36354 30880 36360 30932
rect 36412 30880 36418 30932
rect 36817 30923 36875 30929
rect 36817 30889 36829 30923
rect 36863 30920 36875 30923
rect 37826 30920 37832 30932
rect 36863 30892 37832 30920
rect 36863 30889 36875 30892
rect 36817 30883 36875 30889
rect 37826 30880 37832 30892
rect 37884 30880 37890 30932
rect 17236 30852 17264 30880
rect 17236 30824 18000 30852
rect 17310 30676 17316 30728
rect 17368 30676 17374 30728
rect 17770 30676 17776 30728
rect 17828 30676 17834 30728
rect 17972 30725 18000 30824
rect 18414 30812 18420 30864
rect 18472 30852 18478 30864
rect 19245 30855 19303 30861
rect 19245 30852 19257 30855
rect 18472 30824 19257 30852
rect 18472 30812 18478 30824
rect 19245 30821 19257 30824
rect 19291 30821 19303 30855
rect 19245 30815 19303 30821
rect 21910 30812 21916 30864
rect 21968 30852 21974 30864
rect 22738 30852 22744 30864
rect 21968 30824 22744 30852
rect 21968 30812 21974 30824
rect 22738 30812 22744 30824
rect 22796 30812 22802 30864
rect 25225 30855 25283 30861
rect 25225 30821 25237 30855
rect 25271 30821 25283 30855
rect 25225 30815 25283 30821
rect 33336 30824 34100 30852
rect 25240 30784 25268 30815
rect 25590 30784 25596 30796
rect 25240 30756 25596 30784
rect 25590 30744 25596 30756
rect 25648 30744 25654 30796
rect 25869 30787 25927 30793
rect 25869 30753 25881 30787
rect 25915 30784 25927 30787
rect 27433 30787 27491 30793
rect 27433 30784 27445 30787
rect 25915 30756 27445 30784
rect 25915 30753 25927 30756
rect 25869 30747 25927 30753
rect 27433 30753 27445 30756
rect 27479 30753 27491 30787
rect 27433 30747 27491 30753
rect 27709 30787 27767 30793
rect 27709 30753 27721 30787
rect 27755 30784 27767 30787
rect 28994 30784 29000 30796
rect 27755 30756 29000 30784
rect 27755 30753 27767 30756
rect 27709 30747 27767 30753
rect 28994 30744 29000 30756
rect 29052 30744 29058 30796
rect 31021 30787 31079 30793
rect 31021 30753 31033 30787
rect 31067 30784 31079 30787
rect 32030 30784 32036 30796
rect 31067 30756 32036 30784
rect 31067 30753 31079 30756
rect 31021 30747 31079 30753
rect 32030 30744 32036 30756
rect 32088 30744 32094 30796
rect 17957 30719 18015 30725
rect 17957 30685 17969 30719
rect 18003 30685 18015 30719
rect 17957 30679 18015 30685
rect 18506 30676 18512 30728
rect 18564 30716 18570 30728
rect 19245 30719 19303 30725
rect 19245 30716 19257 30719
rect 18564 30688 19257 30716
rect 18564 30676 18570 30688
rect 19245 30685 19257 30688
rect 19291 30685 19303 30719
rect 19245 30679 19303 30685
rect 19426 30676 19432 30728
rect 19484 30676 19490 30728
rect 22186 30676 22192 30728
rect 22244 30716 22250 30728
rect 22833 30719 22891 30725
rect 22833 30716 22845 30719
rect 22244 30688 22845 30716
rect 22244 30676 22250 30688
rect 22833 30685 22845 30688
rect 22879 30685 22891 30719
rect 22833 30679 22891 30685
rect 22922 30676 22928 30728
rect 22980 30676 22986 30728
rect 23109 30719 23167 30725
rect 23109 30685 23121 30719
rect 23155 30716 23167 30719
rect 24394 30716 24400 30728
rect 23155 30688 24400 30716
rect 23155 30685 23167 30688
rect 23109 30679 23167 30685
rect 24394 30676 24400 30688
rect 24452 30676 24458 30728
rect 25498 30676 25504 30728
rect 25556 30676 25562 30728
rect 30466 30676 30472 30728
rect 30524 30676 30530 30728
rect 30558 30676 30564 30728
rect 30616 30676 30622 30728
rect 32766 30676 32772 30728
rect 32824 30716 32830 30728
rect 33336 30725 33364 30824
rect 33502 30744 33508 30796
rect 33560 30744 33566 30796
rect 34072 30793 34100 30824
rect 34146 30812 34152 30864
rect 34204 30852 34210 30864
rect 34204 30824 34284 30852
rect 34204 30812 34210 30824
rect 34059 30787 34117 30793
rect 34059 30753 34071 30787
rect 34105 30753 34117 30787
rect 34059 30747 34117 30753
rect 33321 30719 33379 30725
rect 33321 30716 33333 30719
rect 32824 30688 33333 30716
rect 32824 30676 32830 30688
rect 33321 30685 33333 30688
rect 33367 30685 33379 30719
rect 33321 30679 33379 30685
rect 33597 30719 33655 30725
rect 33597 30685 33609 30719
rect 33643 30716 33655 30719
rect 34256 30716 34284 30824
rect 34606 30744 34612 30796
rect 34664 30784 34670 30796
rect 34664 30756 35112 30784
rect 34664 30744 34670 30756
rect 33643 30688 34284 30716
rect 34425 30719 34483 30725
rect 33643 30685 33655 30688
rect 33597 30679 33655 30685
rect 34425 30685 34437 30719
rect 34471 30716 34483 30719
rect 34698 30716 34704 30728
rect 34471 30688 34704 30716
rect 34471 30685 34483 30688
rect 34425 30679 34483 30685
rect 34698 30676 34704 30688
rect 34756 30676 34762 30728
rect 35084 30725 35112 30756
rect 34885 30719 34943 30725
rect 34885 30685 34897 30719
rect 34931 30685 34943 30719
rect 34885 30679 34943 30685
rect 35069 30719 35127 30725
rect 35069 30685 35081 30719
rect 35115 30716 35127 30719
rect 36541 30719 36599 30725
rect 36541 30716 36553 30719
rect 35115 30688 36553 30716
rect 35115 30685 35127 30688
rect 35069 30679 35127 30685
rect 36541 30685 36553 30688
rect 36587 30685 36599 30719
rect 36541 30679 36599 30685
rect 16482 30608 16488 30660
rect 16540 30608 16546 30660
rect 17037 30651 17095 30657
rect 17037 30617 17049 30651
rect 17083 30648 17095 30651
rect 18230 30648 18236 30660
rect 17083 30620 18236 30648
rect 17083 30617 17095 30620
rect 17037 30611 17095 30617
rect 18230 30608 18236 30620
rect 18288 30608 18294 30660
rect 24854 30608 24860 30660
rect 24912 30608 24918 30660
rect 27430 30648 27436 30660
rect 27002 30620 27436 30648
rect 27430 30608 27436 30620
rect 27488 30608 27494 30660
rect 31297 30651 31355 30657
rect 31297 30617 31309 30651
rect 31343 30617 31355 30651
rect 31297 30611 31355 30617
rect 17954 30540 17960 30592
rect 18012 30580 18018 30592
rect 18141 30583 18199 30589
rect 18141 30580 18153 30583
rect 18012 30552 18153 30580
rect 18012 30540 18018 30552
rect 18141 30549 18153 30552
rect 18187 30580 18199 30583
rect 18690 30580 18696 30592
rect 18187 30552 18696 30580
rect 18187 30549 18199 30552
rect 18141 30543 18199 30549
rect 18690 30540 18696 30552
rect 18748 30540 18754 30592
rect 22738 30540 22744 30592
rect 22796 30580 22802 30592
rect 24670 30580 24676 30592
rect 22796 30552 24676 30580
rect 22796 30540 22802 30552
rect 24670 30540 24676 30552
rect 24728 30580 24734 30592
rect 25057 30583 25115 30589
rect 25057 30580 25069 30583
rect 24728 30552 25069 30580
rect 24728 30540 24734 30552
rect 25057 30549 25069 30552
rect 25103 30549 25115 30583
rect 31312 30580 31340 30611
rect 31570 30608 31576 30660
rect 31628 30648 31634 30660
rect 33962 30648 33968 30660
rect 31628 30620 31786 30648
rect 32784 30620 33968 30648
rect 31628 30608 31634 30620
rect 32214 30580 32220 30592
rect 31312 30552 32220 30580
rect 25057 30543 25115 30549
rect 32214 30540 32220 30552
rect 32272 30540 32278 30592
rect 32784 30589 32812 30620
rect 33962 30608 33968 30620
rect 34020 30648 34026 30660
rect 34900 30648 34928 30679
rect 34020 30620 34928 30648
rect 34020 30608 34026 30620
rect 35342 30608 35348 30660
rect 35400 30608 35406 30660
rect 32769 30583 32827 30589
rect 32769 30549 32781 30583
rect 32815 30549 32827 30583
rect 32769 30543 32827 30549
rect 33137 30583 33195 30589
rect 33137 30549 33149 30583
rect 33183 30580 33195 30583
rect 33226 30580 33232 30592
rect 33183 30552 33232 30580
rect 33183 30549 33195 30552
rect 33137 30543 33195 30549
rect 33226 30540 33232 30552
rect 33284 30540 33290 30592
rect 33778 30540 33784 30592
rect 33836 30540 33842 30592
rect 33870 30540 33876 30592
rect 33928 30580 33934 30592
rect 34701 30583 34759 30589
rect 34701 30580 34713 30583
rect 33928 30552 34713 30580
rect 33928 30540 33934 30552
rect 34701 30549 34713 30552
rect 34747 30549 34759 30583
rect 36556 30580 36584 30679
rect 36630 30676 36636 30728
rect 36688 30676 36694 30728
rect 36906 30676 36912 30728
rect 36964 30676 36970 30728
rect 37185 30651 37243 30657
rect 37185 30617 37197 30651
rect 37231 30648 37243 30651
rect 37274 30648 37280 30660
rect 37231 30620 37280 30648
rect 37231 30617 37243 30620
rect 37185 30611 37243 30617
rect 37274 30608 37280 30620
rect 37332 30608 37338 30660
rect 38562 30648 38568 30660
rect 38410 30620 38568 30648
rect 38562 30608 38568 30620
rect 38620 30608 38626 30660
rect 38746 30608 38752 30660
rect 38804 30608 38810 30660
rect 36814 30580 36820 30592
rect 36556 30552 36820 30580
rect 34701 30543 34759 30549
rect 36814 30540 36820 30552
rect 36872 30580 36878 30592
rect 38657 30583 38715 30589
rect 38657 30580 38669 30583
rect 36872 30552 38669 30580
rect 36872 30540 36878 30552
rect 38657 30549 38669 30552
rect 38703 30580 38715 30583
rect 38838 30580 38844 30592
rect 38703 30552 38844 30580
rect 38703 30549 38715 30552
rect 38657 30543 38715 30549
rect 38838 30540 38844 30552
rect 38896 30540 38902 30592
rect 1104 30490 58880 30512
rect 1104 30438 4874 30490
rect 4926 30438 4938 30490
rect 4990 30438 5002 30490
rect 5054 30438 5066 30490
rect 5118 30438 5130 30490
rect 5182 30438 35594 30490
rect 35646 30438 35658 30490
rect 35710 30438 35722 30490
rect 35774 30438 35786 30490
rect 35838 30438 35850 30490
rect 35902 30438 58880 30490
rect 1104 30416 58880 30438
rect 19794 30336 19800 30388
rect 19852 30336 19858 30388
rect 24305 30379 24363 30385
rect 24305 30345 24317 30379
rect 24351 30376 24363 30379
rect 24854 30376 24860 30388
rect 24351 30348 24860 30376
rect 24351 30345 24363 30348
rect 24305 30339 24363 30345
rect 24854 30336 24860 30348
rect 24912 30336 24918 30388
rect 25038 30336 25044 30388
rect 25096 30336 25102 30388
rect 27430 30376 27436 30388
rect 26160 30348 27436 30376
rect 18325 30311 18383 30317
rect 18325 30277 18337 30311
rect 18371 30308 18383 30311
rect 18414 30308 18420 30320
rect 18371 30280 18420 30308
rect 18371 30277 18383 30280
rect 18325 30271 18383 30277
rect 18414 30268 18420 30280
rect 18472 30268 18478 30320
rect 19981 30311 20039 30317
rect 19981 30308 19993 30311
rect 19550 30294 19993 30308
rect 19536 30280 19993 30294
rect 17310 30200 17316 30252
rect 17368 30240 17374 30252
rect 18049 30243 18107 30249
rect 18049 30240 18061 30243
rect 17368 30212 18061 30240
rect 17368 30200 17374 30212
rect 18049 30209 18061 30212
rect 18095 30209 18107 30243
rect 18049 30203 18107 30209
rect 18690 30132 18696 30184
rect 18748 30172 18754 30184
rect 19536 30172 19564 30280
rect 19981 30277 19993 30280
rect 20027 30308 20039 30311
rect 22462 30308 22468 30320
rect 20027 30280 22468 30308
rect 20027 30277 20039 30280
rect 19981 30271 20039 30277
rect 22462 30268 22468 30280
rect 22520 30308 22526 30320
rect 26160 30308 26188 30348
rect 27430 30336 27436 30348
rect 27488 30336 27494 30388
rect 32214 30336 32220 30388
rect 32272 30376 32278 30388
rect 32953 30379 33011 30385
rect 32953 30376 32965 30379
rect 32272 30348 32965 30376
rect 32272 30336 32278 30348
rect 32953 30345 32965 30348
rect 32999 30345 33011 30379
rect 32953 30339 33011 30345
rect 33505 30379 33563 30385
rect 33505 30345 33517 30379
rect 33551 30376 33563 30379
rect 33594 30376 33600 30388
rect 33551 30348 33600 30376
rect 33551 30345 33563 30348
rect 33505 30339 33563 30345
rect 33594 30336 33600 30348
rect 33652 30376 33658 30388
rect 35342 30376 35348 30388
rect 33652 30348 35348 30376
rect 33652 30336 33658 30348
rect 35342 30336 35348 30348
rect 35400 30336 35406 30388
rect 22520 30280 23322 30308
rect 26082 30280 26188 30308
rect 22520 30268 22526 30280
rect 26234 30268 26240 30320
rect 26292 30308 26298 30320
rect 26513 30311 26571 30317
rect 26513 30308 26525 30311
rect 26292 30280 26525 30308
rect 26292 30268 26298 30280
rect 26513 30277 26525 30280
rect 26559 30277 26571 30311
rect 26513 30271 26571 30277
rect 32582 30268 32588 30320
rect 32640 30308 32646 30320
rect 32677 30311 32735 30317
rect 32677 30308 32689 30311
rect 32640 30280 32689 30308
rect 32640 30268 32646 30280
rect 32677 30277 32689 30280
rect 32723 30277 32735 30311
rect 32677 30271 32735 30277
rect 33321 30311 33379 30317
rect 33321 30277 33333 30311
rect 33367 30308 33379 30311
rect 33781 30311 33839 30317
rect 33781 30308 33793 30311
rect 33367 30280 33793 30308
rect 33367 30277 33379 30280
rect 33321 30271 33379 30277
rect 33781 30277 33793 30280
rect 33827 30308 33839 30311
rect 33870 30308 33876 30320
rect 33827 30280 33876 30308
rect 33827 30277 33839 30280
rect 33781 30271 33839 30277
rect 33870 30268 33876 30280
rect 33928 30268 33934 30320
rect 33981 30311 34039 30317
rect 33981 30308 33993 30311
rect 33980 30277 33993 30308
rect 34027 30277 34039 30311
rect 33980 30271 34039 30277
rect 22094 30200 22100 30252
rect 22152 30240 22158 30252
rect 22557 30243 22615 30249
rect 22557 30240 22569 30243
rect 22152 30212 22569 30240
rect 22152 30200 22158 30212
rect 22557 30209 22569 30212
rect 22603 30209 22615 30243
rect 22557 30203 22615 30209
rect 32953 30243 33011 30249
rect 32953 30209 32965 30243
rect 32999 30209 33011 30243
rect 32953 30203 33011 30209
rect 33597 30243 33655 30249
rect 33597 30209 33609 30243
rect 33643 30240 33655 30243
rect 33980 30240 34008 30271
rect 36630 30268 36636 30320
rect 36688 30308 36694 30320
rect 38657 30311 38715 30317
rect 38657 30308 38669 30311
rect 36688 30280 38669 30308
rect 36688 30268 36694 30280
rect 38657 30277 38669 30280
rect 38703 30277 38715 30311
rect 38657 30271 38715 30277
rect 38838 30268 38844 30320
rect 38896 30268 38902 30320
rect 42245 30311 42303 30317
rect 42245 30277 42257 30311
rect 42291 30308 42303 30311
rect 42291 30280 42564 30308
rect 42291 30277 42303 30280
rect 42245 30271 42303 30277
rect 42536 30252 42564 30280
rect 43346 30268 43352 30320
rect 43404 30308 43410 30320
rect 43404 30280 43562 30308
rect 43404 30268 43410 30280
rect 34146 30240 34152 30252
rect 33643 30212 34152 30240
rect 33643 30209 33655 30212
rect 33597 30203 33655 30209
rect 18748 30144 19564 30172
rect 18748 30132 18754 30144
rect 22830 30132 22836 30184
rect 22888 30132 22894 30184
rect 26789 30175 26847 30181
rect 26789 30141 26801 30175
rect 26835 30172 26847 30175
rect 28258 30172 28264 30184
rect 26835 30144 28264 30172
rect 26835 30141 26847 30144
rect 26789 30135 26847 30141
rect 28258 30132 28264 30144
rect 28316 30132 28322 30184
rect 32968 30172 32996 30203
rect 33796 30184 33824 30212
rect 34146 30200 34152 30212
rect 34204 30200 34210 30252
rect 38562 30200 38568 30252
rect 38620 30200 38626 30252
rect 42426 30200 42432 30252
rect 42484 30200 42490 30252
rect 42518 30200 42524 30252
rect 42576 30200 42582 30252
rect 42702 30200 42708 30252
rect 42760 30200 42766 30252
rect 32968 30144 33364 30172
rect 33336 30113 33364 30144
rect 33778 30132 33784 30184
rect 33836 30132 33842 30184
rect 36906 30132 36912 30184
rect 36964 30172 36970 30184
rect 37829 30175 37887 30181
rect 37829 30172 37841 30175
rect 36964 30144 37841 30172
rect 36964 30132 36970 30144
rect 37829 30141 37841 30144
rect 37875 30172 37887 30175
rect 38746 30172 38752 30184
rect 37875 30144 38752 30172
rect 37875 30141 37887 30144
rect 37829 30135 37887 30141
rect 38746 30132 38752 30144
rect 38804 30172 38810 30184
rect 42797 30175 42855 30181
rect 42797 30172 42809 30175
rect 38804 30144 42809 30172
rect 38804 30132 38810 30144
rect 42797 30141 42809 30144
rect 42843 30141 42855 30175
rect 43073 30175 43131 30181
rect 43073 30172 43085 30175
rect 42797 30135 42855 30141
rect 42904 30144 43085 30172
rect 32861 30107 32919 30113
rect 32861 30073 32873 30107
rect 32907 30073 32919 30107
rect 32861 30067 32919 30073
rect 33321 30107 33379 30113
rect 33321 30073 33333 30107
rect 33367 30073 33379 30107
rect 34149 30107 34207 30113
rect 34149 30104 34161 30107
rect 33321 30067 33379 30073
rect 33520 30076 34161 30104
rect 25222 29996 25228 30048
rect 25280 30036 25286 30048
rect 29638 30036 29644 30048
rect 25280 30008 29644 30036
rect 25280 29996 25286 30008
rect 29638 29996 29644 30008
rect 29696 29996 29702 30048
rect 32876 30036 32904 30067
rect 33520 30036 33548 30076
rect 34149 30073 34161 30076
rect 34195 30104 34207 30107
rect 36630 30104 36636 30116
rect 34195 30076 36636 30104
rect 34195 30073 34207 30076
rect 34149 30067 34207 30073
rect 36630 30064 36636 30076
rect 36688 30064 36694 30116
rect 38562 30064 38568 30116
rect 38620 30104 38626 30116
rect 39117 30107 39175 30113
rect 39117 30104 39129 30107
rect 38620 30076 39129 30104
rect 38620 30064 38626 30076
rect 39117 30073 39129 30076
rect 39163 30073 39175 30107
rect 39117 30067 39175 30073
rect 42705 30107 42763 30113
rect 42705 30073 42717 30107
rect 42751 30104 42763 30107
rect 42904 30104 42932 30144
rect 43073 30141 43085 30144
rect 43119 30141 43131 30175
rect 43073 30135 43131 30141
rect 44726 30132 44732 30184
rect 44784 30172 44790 30184
rect 44821 30175 44879 30181
rect 44821 30172 44833 30175
rect 44784 30144 44833 30172
rect 44784 30132 44790 30144
rect 44821 30141 44833 30144
rect 44867 30141 44879 30175
rect 44821 30135 44879 30141
rect 42751 30076 42932 30104
rect 42751 30073 42763 30076
rect 42705 30067 42763 30073
rect 32876 30008 33548 30036
rect 33594 29996 33600 30048
rect 33652 30036 33658 30048
rect 33962 30036 33968 30048
rect 33652 30008 33968 30036
rect 33652 29996 33658 30008
rect 33962 29996 33968 30008
rect 34020 29996 34026 30048
rect 34606 29996 34612 30048
rect 34664 30036 34670 30048
rect 36538 30036 36544 30048
rect 34664 30008 36544 30036
rect 34664 29996 34670 30008
rect 36538 29996 36544 30008
rect 36596 29996 36602 30048
rect 37458 29996 37464 30048
rect 37516 30036 37522 30048
rect 39025 30039 39083 30045
rect 39025 30036 39037 30039
rect 37516 30008 39037 30036
rect 37516 29996 37522 30008
rect 39025 30005 39037 30008
rect 39071 30005 39083 30039
rect 39025 29999 39083 30005
rect 1104 29946 58880 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 58880 29946
rect 1104 29872 58880 29894
rect 22557 29835 22615 29841
rect 22557 29801 22569 29835
rect 22603 29832 22615 29835
rect 22830 29832 22836 29844
rect 22603 29804 22836 29832
rect 22603 29801 22615 29804
rect 22557 29795 22615 29801
rect 22830 29792 22836 29804
rect 22888 29792 22894 29844
rect 28810 29792 28816 29844
rect 28868 29792 28874 29844
rect 32122 29832 32128 29844
rect 28920 29804 32128 29832
rect 16850 29724 16856 29776
rect 16908 29764 16914 29776
rect 25222 29764 25228 29776
rect 16908 29736 25228 29764
rect 16908 29724 16914 29736
rect 25222 29724 25228 29736
rect 25280 29724 25286 29776
rect 22738 29656 22744 29708
rect 22796 29696 22802 29708
rect 22833 29699 22891 29705
rect 22833 29696 22845 29699
rect 22796 29668 22845 29696
rect 22796 29656 22802 29668
rect 22833 29665 22845 29668
rect 22879 29665 22891 29699
rect 22833 29659 22891 29665
rect 24854 29656 24860 29708
rect 24912 29696 24918 29708
rect 24949 29699 25007 29705
rect 24949 29696 24961 29699
rect 24912 29668 24961 29696
rect 24912 29656 24918 29668
rect 24949 29665 24961 29668
rect 24995 29665 25007 29699
rect 24949 29659 25007 29665
rect 22925 29631 22983 29637
rect 22925 29597 22937 29631
rect 22971 29628 22983 29631
rect 24397 29631 24455 29637
rect 24397 29628 24409 29631
rect 22971 29600 24409 29628
rect 22971 29597 22983 29600
rect 22925 29591 22983 29597
rect 24397 29597 24409 29600
rect 24443 29597 24455 29631
rect 24397 29591 24455 29597
rect 27154 29520 27160 29572
rect 27212 29560 27218 29572
rect 28920 29560 28948 29804
rect 32122 29792 32128 29804
rect 32180 29832 32186 29844
rect 32950 29832 32956 29844
rect 32180 29804 32956 29832
rect 32180 29792 32186 29804
rect 32950 29792 32956 29804
rect 33008 29792 33014 29844
rect 34241 29835 34299 29841
rect 34241 29801 34253 29835
rect 34287 29832 34299 29835
rect 35069 29835 35127 29841
rect 35069 29832 35081 29835
rect 34287 29804 35081 29832
rect 34287 29801 34299 29804
rect 34241 29795 34299 29801
rect 35069 29801 35081 29804
rect 35115 29801 35127 29835
rect 35069 29795 35127 29801
rect 37274 29792 37280 29844
rect 37332 29792 37338 29844
rect 37461 29835 37519 29841
rect 37461 29801 37473 29835
rect 37507 29832 37519 29835
rect 37550 29832 37556 29844
rect 37507 29804 37556 29832
rect 37507 29801 37519 29804
rect 37461 29795 37519 29801
rect 37550 29792 37556 29804
rect 37608 29792 37614 29844
rect 42518 29832 42524 29844
rect 40420 29804 42524 29832
rect 29086 29724 29092 29776
rect 29144 29764 29150 29776
rect 29733 29767 29791 29773
rect 29733 29764 29745 29767
rect 29144 29736 29745 29764
rect 29144 29724 29150 29736
rect 29733 29733 29745 29736
rect 29779 29764 29791 29767
rect 32490 29764 32496 29776
rect 29779 29736 32496 29764
rect 29779 29733 29791 29736
rect 29733 29727 29791 29733
rect 32490 29724 32496 29736
rect 32548 29724 32554 29776
rect 33226 29724 33232 29776
rect 33284 29764 33290 29776
rect 33284 29736 35204 29764
rect 33284 29724 33290 29736
rect 29104 29668 29592 29696
rect 29104 29637 29132 29668
rect 29089 29631 29147 29637
rect 29089 29597 29101 29631
rect 29135 29597 29147 29631
rect 29089 29591 29147 29597
rect 29270 29588 29276 29640
rect 29328 29588 29334 29640
rect 29564 29637 29592 29668
rect 29638 29656 29644 29708
rect 29696 29696 29702 29708
rect 29696 29668 35020 29696
rect 29696 29656 29702 29668
rect 29549 29631 29607 29637
rect 29549 29597 29561 29631
rect 29595 29628 29607 29631
rect 30006 29628 30012 29640
rect 29595 29600 30012 29628
rect 29595 29597 29607 29600
rect 29549 29591 29607 29597
rect 30006 29588 30012 29600
rect 30064 29588 30070 29640
rect 33778 29588 33784 29640
rect 33836 29588 33842 29640
rect 33962 29588 33968 29640
rect 34020 29628 34026 29640
rect 34885 29631 34943 29637
rect 34885 29628 34897 29631
rect 34020 29600 34897 29628
rect 34020 29588 34026 29600
rect 34885 29597 34897 29600
rect 34931 29597 34943 29631
rect 34885 29591 34943 29597
rect 28997 29563 29055 29569
rect 28997 29560 29009 29563
rect 27212 29532 29009 29560
rect 27212 29520 27218 29532
rect 28997 29529 29009 29532
rect 29043 29529 29055 29563
rect 29288 29560 29316 29588
rect 29641 29563 29699 29569
rect 29641 29560 29653 29563
rect 29288 29532 29653 29560
rect 28997 29523 29055 29529
rect 29641 29529 29653 29532
rect 29687 29529 29699 29563
rect 29641 29523 29699 29529
rect 29825 29563 29883 29569
rect 29825 29529 29837 29563
rect 29871 29560 29883 29563
rect 30466 29560 30472 29572
rect 29871 29532 30472 29560
rect 29871 29529 29883 29532
rect 29825 29523 29883 29529
rect 30466 29520 30472 29532
rect 30524 29520 30530 29572
rect 32401 29563 32459 29569
rect 32401 29529 32413 29563
rect 32447 29560 32459 29563
rect 32490 29560 32496 29572
rect 32447 29532 32496 29560
rect 32447 29529 32459 29532
rect 32401 29523 32459 29529
rect 32490 29520 32496 29532
rect 32548 29520 32554 29572
rect 32585 29563 32643 29569
rect 32585 29529 32597 29563
rect 32631 29560 32643 29563
rect 32858 29560 32864 29572
rect 32631 29532 32864 29560
rect 32631 29529 32643 29532
rect 32585 29523 32643 29529
rect 32858 29520 32864 29532
rect 32916 29520 32922 29572
rect 32950 29520 32956 29572
rect 33008 29560 33014 29572
rect 34057 29563 34115 29569
rect 34057 29560 34069 29563
rect 33008 29532 34069 29560
rect 33008 29520 33014 29532
rect 34057 29529 34069 29532
rect 34103 29529 34115 29563
rect 34057 29523 34115 29529
rect 34146 29520 34152 29572
rect 34204 29560 34210 29572
rect 34701 29563 34759 29569
rect 34701 29560 34713 29563
rect 34204 29532 34713 29560
rect 34204 29520 34210 29532
rect 34701 29529 34713 29532
rect 34747 29529 34759 29563
rect 34992 29560 35020 29668
rect 35176 29628 35204 29736
rect 37826 29724 37832 29776
rect 37884 29724 37890 29776
rect 38013 29767 38071 29773
rect 38013 29733 38025 29767
rect 38059 29764 38071 29767
rect 40310 29764 40316 29776
rect 38059 29736 40316 29764
rect 38059 29733 38071 29736
rect 38013 29727 38071 29733
rect 40310 29724 40316 29736
rect 40368 29724 40374 29776
rect 38194 29656 38200 29708
rect 38252 29656 38258 29708
rect 40420 29696 40448 29804
rect 42518 29792 42524 29804
rect 42576 29792 42582 29844
rect 42702 29792 42708 29844
rect 42760 29832 42766 29844
rect 43441 29835 43499 29841
rect 43441 29832 43453 29835
rect 42760 29804 43453 29832
rect 42760 29792 42766 29804
rect 43441 29801 43453 29804
rect 43487 29801 43499 29835
rect 43441 29795 43499 29801
rect 40770 29724 40776 29776
rect 40828 29764 40834 29776
rect 40865 29767 40923 29773
rect 40865 29764 40877 29767
rect 40828 29736 40877 29764
rect 40828 29724 40834 29736
rect 40865 29733 40877 29736
rect 40911 29733 40923 29767
rect 40865 29727 40923 29733
rect 38304 29668 40448 29696
rect 40497 29699 40555 29705
rect 37921 29631 37979 29637
rect 37921 29628 37933 29631
rect 35176 29600 37933 29628
rect 37921 29597 37933 29600
rect 37967 29597 37979 29631
rect 37921 29591 37979 29597
rect 34992 29532 35112 29560
rect 34701 29523 34759 29529
rect 28626 29452 28632 29504
rect 28684 29452 28690 29504
rect 28797 29495 28855 29501
rect 28797 29461 28809 29495
rect 28843 29492 28855 29495
rect 29089 29495 29147 29501
rect 29089 29492 29101 29495
rect 28843 29464 29101 29492
rect 28843 29461 28855 29464
rect 28797 29455 28855 29461
rect 29089 29461 29101 29464
rect 29135 29461 29147 29495
rect 29089 29455 29147 29461
rect 32766 29452 32772 29504
rect 32824 29452 32830 29504
rect 33965 29495 34023 29501
rect 33965 29461 33977 29495
rect 34011 29492 34023 29495
rect 34257 29495 34315 29501
rect 34257 29492 34269 29495
rect 34011 29464 34269 29492
rect 34011 29461 34023 29464
rect 33965 29455 34023 29461
rect 34257 29461 34269 29464
rect 34303 29461 34315 29495
rect 34257 29455 34315 29461
rect 34425 29495 34483 29501
rect 34425 29461 34437 29495
rect 34471 29492 34483 29495
rect 34974 29492 34980 29504
rect 34471 29464 34980 29492
rect 34471 29461 34483 29464
rect 34425 29455 34483 29461
rect 34974 29452 34980 29464
rect 35032 29452 35038 29504
rect 35084 29492 35112 29532
rect 37458 29520 37464 29572
rect 37516 29520 37522 29572
rect 38304 29560 38332 29668
rect 40497 29665 40509 29699
rect 40543 29665 40555 29699
rect 40497 29659 40555 29665
rect 41386 29668 44036 29696
rect 39666 29588 39672 29640
rect 39724 29628 39730 29640
rect 40221 29631 40279 29637
rect 40221 29628 40233 29631
rect 39724 29600 40233 29628
rect 39724 29588 39730 29600
rect 40221 29597 40233 29600
rect 40267 29597 40279 29631
rect 40221 29591 40279 29597
rect 40313 29631 40371 29637
rect 40313 29597 40325 29631
rect 40359 29597 40371 29631
rect 40512 29628 40540 29659
rect 40586 29628 40592 29640
rect 40512 29600 40592 29628
rect 40313 29591 40371 29597
rect 37568 29532 38332 29560
rect 40328 29560 40356 29591
rect 40586 29588 40592 29600
rect 40644 29588 40650 29640
rect 41386 29572 41414 29668
rect 42518 29588 42524 29640
rect 42576 29628 42582 29640
rect 43257 29631 43315 29637
rect 43257 29628 43269 29631
rect 42576 29600 43269 29628
rect 42576 29588 42582 29600
rect 43257 29597 43269 29600
rect 43303 29628 43315 29631
rect 43441 29631 43499 29637
rect 43441 29628 43453 29631
rect 43303 29600 43453 29628
rect 43303 29597 43315 29600
rect 43257 29591 43315 29597
rect 43441 29597 43453 29600
rect 43487 29597 43499 29631
rect 43441 29591 43499 29597
rect 43625 29631 43683 29637
rect 43625 29597 43637 29631
rect 43671 29597 43683 29631
rect 43625 29591 43683 29597
rect 40865 29563 40923 29569
rect 40328 29532 40724 29560
rect 37568 29492 37596 29532
rect 35084 29464 37596 29492
rect 37642 29452 37648 29504
rect 37700 29492 37706 29504
rect 38197 29495 38255 29501
rect 38197 29492 38209 29495
rect 37700 29464 38209 29492
rect 37700 29452 37706 29464
rect 38197 29461 38209 29464
rect 38243 29461 38255 29495
rect 38197 29455 38255 29461
rect 40494 29452 40500 29504
rect 40552 29452 40558 29504
rect 40696 29501 40724 29532
rect 40865 29529 40877 29563
rect 40911 29560 40923 29563
rect 41386 29560 41420 29572
rect 40911 29532 41420 29560
rect 40911 29529 40923 29532
rect 40865 29523 40923 29529
rect 41414 29520 41420 29532
rect 41472 29520 41478 29572
rect 42794 29520 42800 29572
rect 42852 29560 42858 29572
rect 43640 29560 43668 29591
rect 44008 29572 44036 29668
rect 44174 29656 44180 29708
rect 44232 29696 44238 29708
rect 44545 29699 44603 29705
rect 44545 29696 44557 29699
rect 44232 29668 44557 29696
rect 44232 29656 44238 29668
rect 44545 29665 44557 29668
rect 44591 29665 44603 29699
rect 44545 29659 44603 29665
rect 44358 29588 44364 29640
rect 44416 29588 44422 29640
rect 47397 29631 47455 29637
rect 47397 29597 47409 29631
rect 47443 29628 47455 29631
rect 49694 29628 49700 29640
rect 47443 29600 49700 29628
rect 47443 29597 47455 29600
rect 47397 29591 47455 29597
rect 49694 29588 49700 29600
rect 49752 29588 49758 29640
rect 42852 29532 43668 29560
rect 42852 29520 42858 29532
rect 40681 29495 40739 29501
rect 40681 29461 40693 29495
rect 40727 29492 40739 29495
rect 41138 29492 41144 29504
rect 40727 29464 41144 29492
rect 40727 29461 40739 29464
rect 40681 29455 40739 29461
rect 41138 29452 41144 29464
rect 41196 29452 41202 29504
rect 41230 29452 41236 29504
rect 41288 29492 41294 29504
rect 42705 29495 42763 29501
rect 42705 29492 42717 29495
rect 41288 29464 42717 29492
rect 41288 29452 41294 29464
rect 42705 29461 42717 29464
rect 42751 29492 42763 29495
rect 43346 29492 43352 29504
rect 42751 29464 43352 29492
rect 42751 29461 42763 29464
rect 42705 29455 42763 29461
rect 43346 29452 43352 29464
rect 43404 29452 43410 29504
rect 43640 29492 43668 29532
rect 43990 29520 43996 29572
rect 44048 29520 44054 29572
rect 44376 29560 44404 29588
rect 45370 29560 45376 29572
rect 44376 29532 45376 29560
rect 45370 29520 45376 29532
rect 45428 29520 45434 29572
rect 46690 29532 47072 29560
rect 44174 29492 44180 29504
rect 43640 29464 44180 29492
rect 44174 29452 44180 29464
rect 44232 29452 44238 29504
rect 47044 29492 47072 29532
rect 47118 29520 47124 29572
rect 47176 29520 47182 29572
rect 47394 29492 47400 29504
rect 47044 29464 47400 29492
rect 47394 29452 47400 29464
rect 47452 29492 47458 29504
rect 47489 29495 47547 29501
rect 47489 29492 47501 29495
rect 47452 29464 47501 29492
rect 47452 29452 47458 29464
rect 47489 29461 47501 29464
rect 47535 29461 47547 29495
rect 47489 29455 47547 29461
rect 1104 29402 58880 29424
rect 1104 29350 4874 29402
rect 4926 29350 4938 29402
rect 4990 29350 5002 29402
rect 5054 29350 5066 29402
rect 5118 29350 5130 29402
rect 5182 29350 35594 29402
rect 35646 29350 35658 29402
rect 35710 29350 35722 29402
rect 35774 29350 35786 29402
rect 35838 29350 35850 29402
rect 35902 29350 58880 29402
rect 1104 29328 58880 29350
rect 27154 29248 27160 29300
rect 27212 29288 27218 29300
rect 27212 29260 28304 29288
rect 27212 29248 27218 29260
rect 27172 29152 27200 29248
rect 28276 29229 28304 29260
rect 28368 29260 30420 29288
rect 27341 29223 27399 29229
rect 27341 29189 27353 29223
rect 27387 29220 27399 29223
rect 27525 29223 27583 29229
rect 27525 29220 27537 29223
rect 27387 29192 27537 29220
rect 27387 29189 27399 29192
rect 27341 29183 27399 29189
rect 27525 29189 27537 29192
rect 27571 29220 27583 29223
rect 28261 29223 28319 29229
rect 27571 29192 28212 29220
rect 27571 29189 27583 29192
rect 27525 29183 27583 29189
rect 26252 29124 27200 29152
rect 27893 29155 27951 29161
rect 26252 29025 26280 29124
rect 27893 29121 27905 29155
rect 27939 29152 27951 29155
rect 28184 29152 28212 29192
rect 28261 29189 28273 29223
rect 28307 29189 28319 29223
rect 28261 29183 28319 29189
rect 28368 29152 28396 29260
rect 28477 29223 28535 29229
rect 28477 29189 28489 29223
rect 28523 29220 28535 29223
rect 29086 29220 29092 29232
rect 28523 29192 29092 29220
rect 28523 29189 28535 29192
rect 28477 29183 28535 29189
rect 29086 29180 29092 29192
rect 29144 29180 29150 29232
rect 29380 29220 29408 29260
rect 30392 29220 30420 29260
rect 30466 29248 30472 29300
rect 30524 29248 30530 29300
rect 31726 29260 33732 29288
rect 31570 29220 31576 29232
rect 29380 29192 29486 29220
rect 30392 29192 31576 29220
rect 31570 29180 31576 29192
rect 31628 29220 31634 29232
rect 31726 29220 31754 29260
rect 32490 29220 32496 29232
rect 31628 29192 31754 29220
rect 31864 29192 32496 29220
rect 31628 29180 31634 29192
rect 27939 29124 28120 29152
rect 28184 29124 28396 29152
rect 31757 29155 31815 29161
rect 27939 29121 27951 29124
rect 27893 29115 27951 29121
rect 26510 29044 26516 29096
rect 26568 29044 26574 29096
rect 28092 29028 28120 29124
rect 31757 29121 31769 29155
rect 31803 29152 31815 29155
rect 31864 29152 31892 29192
rect 32490 29180 32496 29192
rect 32548 29180 32554 29232
rect 33704 29220 33732 29260
rect 33962 29248 33968 29300
rect 34020 29248 34026 29300
rect 37093 29291 37151 29297
rect 37093 29257 37105 29291
rect 37139 29288 37151 29291
rect 38010 29288 38016 29300
rect 37139 29260 38016 29288
rect 37139 29257 37151 29260
rect 37093 29251 37151 29257
rect 38010 29248 38016 29260
rect 38068 29288 38074 29300
rect 38654 29288 38660 29300
rect 38068 29260 38660 29288
rect 38068 29248 38074 29260
rect 38654 29248 38660 29260
rect 38712 29288 38718 29300
rect 40405 29291 40463 29297
rect 38712 29260 38976 29288
rect 38712 29248 38718 29260
rect 33626 29192 34270 29220
rect 37642 29180 37648 29232
rect 37700 29180 37706 29232
rect 38948 29220 38976 29260
rect 40405 29257 40417 29291
rect 40451 29288 40463 29291
rect 41138 29288 41144 29300
rect 40451 29260 41144 29288
rect 40451 29257 40463 29260
rect 40405 29251 40463 29257
rect 41138 29248 41144 29260
rect 41196 29248 41202 29300
rect 42886 29288 42892 29300
rect 41386 29260 42892 29288
rect 41046 29220 41052 29232
rect 38870 29192 41052 29220
rect 41046 29180 41052 29192
rect 41104 29180 41110 29232
rect 41386 29220 41414 29260
rect 42886 29248 42892 29260
rect 42944 29288 42950 29300
rect 43809 29291 43867 29297
rect 43809 29288 43821 29291
rect 42944 29260 43821 29288
rect 42944 29248 42950 29260
rect 43809 29257 43821 29260
rect 43855 29257 43867 29291
rect 43809 29251 43867 29257
rect 45370 29248 45376 29300
rect 45428 29288 45434 29300
rect 46017 29291 46075 29297
rect 46017 29288 46029 29291
rect 45428 29260 46029 29288
rect 45428 29248 45434 29260
rect 46017 29257 46029 29260
rect 46063 29257 46075 29291
rect 46017 29251 46075 29257
rect 46477 29291 46535 29297
rect 46477 29257 46489 29291
rect 46523 29288 46535 29291
rect 47118 29288 47124 29300
rect 46523 29260 47124 29288
rect 46523 29257 46535 29260
rect 46477 29251 46535 29257
rect 47118 29248 47124 29260
rect 47176 29248 47182 29300
rect 41156 29192 41414 29220
rect 31803 29124 31892 29152
rect 31941 29155 31999 29161
rect 31803 29121 31815 29124
rect 31757 29115 31815 29121
rect 31941 29121 31953 29155
rect 31987 29121 31999 29155
rect 31941 29115 31999 29121
rect 28258 29044 28264 29096
rect 28316 29084 28322 29096
rect 28721 29087 28779 29093
rect 28721 29084 28733 29087
rect 28316 29056 28733 29084
rect 28316 29044 28322 29056
rect 28721 29053 28733 29056
rect 28767 29053 28779 29087
rect 28997 29087 29055 29093
rect 28997 29084 29009 29087
rect 28721 29047 28779 29053
rect 28828 29056 29009 29084
rect 26237 29019 26295 29025
rect 26237 28985 26249 29019
rect 26283 28985 26295 29019
rect 26237 28979 26295 28985
rect 27157 29019 27215 29025
rect 27157 28985 27169 29019
rect 27203 29016 27215 29019
rect 27430 29016 27436 29028
rect 27203 28988 27436 29016
rect 27203 28985 27215 28988
rect 27157 28979 27215 28985
rect 27430 28976 27436 28988
rect 27488 28976 27494 29028
rect 28074 28976 28080 29028
rect 28132 28976 28138 29028
rect 28629 29019 28687 29025
rect 28629 28985 28641 29019
rect 28675 29016 28687 29019
rect 28828 29016 28856 29056
rect 28997 29053 29009 29056
rect 29043 29053 29055 29087
rect 31956 29084 31984 29115
rect 32030 29112 32036 29164
rect 32088 29152 32094 29164
rect 32125 29155 32183 29161
rect 32125 29152 32137 29155
rect 32088 29124 32137 29152
rect 32088 29112 32094 29124
rect 32125 29121 32137 29124
rect 32171 29121 32183 29155
rect 32125 29115 32183 29121
rect 35713 29155 35771 29161
rect 35713 29121 35725 29155
rect 35759 29152 35771 29155
rect 35986 29152 35992 29164
rect 35759 29124 35992 29152
rect 35759 29121 35771 29124
rect 35713 29115 35771 29121
rect 35986 29112 35992 29124
rect 36044 29152 36050 29164
rect 36906 29152 36912 29164
rect 36044 29124 36912 29152
rect 36044 29112 36050 29124
rect 36906 29112 36912 29124
rect 36964 29152 36970 29164
rect 37369 29155 37427 29161
rect 37369 29152 37381 29155
rect 36964 29124 37381 29152
rect 36964 29112 36970 29124
rect 37369 29121 37381 29124
rect 37415 29121 37427 29155
rect 37369 29115 37427 29121
rect 39393 29155 39451 29161
rect 39393 29121 39405 29155
rect 39439 29152 39451 29155
rect 39761 29155 39819 29161
rect 39761 29152 39773 29155
rect 39439 29124 39773 29152
rect 39439 29121 39451 29124
rect 39393 29115 39451 29121
rect 39761 29121 39773 29124
rect 39807 29152 39819 29155
rect 39942 29152 39948 29164
rect 39807 29124 39948 29152
rect 39807 29121 39819 29124
rect 39761 29115 39819 29121
rect 39942 29112 39948 29124
rect 40000 29112 40006 29164
rect 40218 29161 40224 29164
rect 40037 29155 40095 29161
rect 40037 29121 40049 29155
rect 40083 29121 40095 29155
rect 40037 29115 40095 29121
rect 40191 29155 40224 29161
rect 40191 29121 40203 29155
rect 40191 29115 40224 29121
rect 31956 29056 32076 29084
rect 28997 29047 29055 29053
rect 28675 28988 28856 29016
rect 28675 28985 28687 28988
rect 28629 28979 28687 28985
rect 25958 28908 25964 28960
rect 26016 28948 26022 28960
rect 26053 28951 26111 28957
rect 26053 28948 26065 28951
rect 26016 28920 26065 28948
rect 26016 28908 26022 28920
rect 26053 28917 26065 28920
rect 26099 28917 26111 28951
rect 26053 28911 26111 28917
rect 28445 28951 28503 28957
rect 28445 28917 28457 28951
rect 28491 28948 28503 28951
rect 30650 28948 30656 28960
rect 28491 28920 30656 28948
rect 28491 28917 28503 28920
rect 28445 28911 28503 28917
rect 30650 28908 30656 28920
rect 30708 28908 30714 28960
rect 31846 28908 31852 28960
rect 31904 28908 31910 28960
rect 32048 28948 32076 29056
rect 32398 29044 32404 29096
rect 32456 29044 32462 29096
rect 34974 29044 34980 29096
rect 35032 29084 35038 29096
rect 35437 29087 35495 29093
rect 35437 29084 35449 29087
rect 35032 29056 35449 29084
rect 35032 29044 35038 29056
rect 35437 29053 35449 29056
rect 35483 29053 35495 29087
rect 40052 29084 40080 29115
rect 40218 29112 40224 29115
rect 40276 29112 40282 29164
rect 40310 29112 40316 29164
rect 40368 29152 40374 29164
rect 40589 29155 40647 29161
rect 40589 29152 40601 29155
rect 40368 29124 40601 29152
rect 40368 29112 40374 29124
rect 40589 29121 40601 29124
rect 40635 29121 40647 29155
rect 40589 29115 40647 29121
rect 40770 29112 40776 29164
rect 40828 29112 40834 29164
rect 41156 29161 41184 29192
rect 42978 29180 42984 29232
rect 43036 29180 43042 29232
rect 43898 29220 43904 29232
rect 43364 29192 43904 29220
rect 40865 29155 40923 29161
rect 40865 29121 40877 29155
rect 40911 29121 40923 29155
rect 40865 29115 40923 29121
rect 41141 29155 41199 29161
rect 41141 29121 41153 29155
rect 41187 29121 41199 29155
rect 41141 29115 41199 29121
rect 40402 29084 40408 29096
rect 40052 29056 40408 29084
rect 35437 29047 35495 29053
rect 40402 29044 40408 29056
rect 40460 29044 40466 29096
rect 40880 29084 40908 29115
rect 41414 29112 41420 29164
rect 41472 29112 41478 29164
rect 41509 29155 41567 29161
rect 41509 29121 41521 29155
rect 41555 29121 41567 29155
rect 41509 29115 41567 29121
rect 41233 29087 41291 29093
rect 41233 29084 41245 29087
rect 40880 29056 41245 29084
rect 41233 29053 41245 29056
rect 41279 29053 41291 29087
rect 41233 29047 41291 29053
rect 41322 29044 41328 29096
rect 41380 29084 41386 29096
rect 41524 29084 41552 29115
rect 41380 29056 41552 29084
rect 41601 29087 41659 29093
rect 41380 29044 41386 29056
rect 41601 29053 41613 29087
rect 41647 29053 41659 29087
rect 41601 29047 41659 29053
rect 41693 29087 41751 29093
rect 41693 29053 41705 29087
rect 41739 29084 41751 29087
rect 43364 29084 43392 29192
rect 43898 29180 43904 29192
rect 43956 29220 43962 29232
rect 43956 29192 44128 29220
rect 43956 29180 43962 29192
rect 43441 29155 43499 29161
rect 43441 29121 43453 29155
rect 43487 29152 43499 29155
rect 43714 29152 43720 29164
rect 43487 29124 43720 29152
rect 43487 29121 43499 29124
rect 43441 29115 43499 29121
rect 43714 29112 43720 29124
rect 43772 29112 43778 29164
rect 44100 29161 44128 29192
rect 43993 29155 44051 29161
rect 43993 29121 44005 29155
rect 44039 29121 44051 29155
rect 43993 29115 44051 29121
rect 44085 29155 44143 29161
rect 44085 29121 44097 29155
rect 44131 29121 44143 29155
rect 44085 29115 44143 29121
rect 41739 29056 43392 29084
rect 41739 29053 41751 29056
rect 41693 29047 41751 29053
rect 40494 28976 40500 29028
rect 40552 29016 40558 29028
rect 41049 29019 41107 29025
rect 41049 29016 41061 29019
rect 40552 28988 41061 29016
rect 40552 28976 40558 28988
rect 41049 28985 41061 28988
rect 41095 28985 41107 29019
rect 41049 28979 41107 28985
rect 41138 28976 41144 29028
rect 41196 29016 41202 29028
rect 41616 29016 41644 29047
rect 43530 29044 43536 29096
rect 43588 29084 43594 29096
rect 44008 29084 44036 29115
rect 44174 29112 44180 29164
rect 44232 29152 44238 29164
rect 44726 29152 44732 29164
rect 44232 29124 44732 29152
rect 44232 29112 44238 29124
rect 44726 29112 44732 29124
rect 44784 29112 44790 29164
rect 46106 29112 46112 29164
rect 46164 29112 46170 29164
rect 44358 29084 44364 29096
rect 43588 29056 44364 29084
rect 43588 29044 43594 29056
rect 44358 29044 44364 29056
rect 44416 29044 44422 29096
rect 45649 29087 45707 29093
rect 45649 29053 45661 29087
rect 45695 29084 45707 29087
rect 45922 29084 45928 29096
rect 45695 29056 45928 29084
rect 45695 29053 45707 29056
rect 45649 29047 45707 29053
rect 45922 29044 45928 29056
rect 45980 29044 45986 29096
rect 41196 28988 41644 29016
rect 42981 29019 43039 29025
rect 41196 28976 41202 28988
rect 42981 28985 42993 29019
rect 43027 29016 43039 29019
rect 43806 29016 43812 29028
rect 43027 28988 43812 29016
rect 43027 28985 43039 28988
rect 42981 28979 43039 28985
rect 43806 28976 43812 28988
rect 43864 28976 43870 29028
rect 32858 28948 32864 28960
rect 32048 28920 32864 28948
rect 32858 28908 32864 28920
rect 32916 28908 32922 28960
rect 33134 28908 33140 28960
rect 33192 28948 33198 28960
rect 33873 28951 33931 28957
rect 33873 28948 33885 28951
rect 33192 28920 33885 28948
rect 33192 28908 33198 28920
rect 33873 28917 33885 28920
rect 33919 28917 33931 28951
rect 33873 28911 33931 28917
rect 39666 28908 39672 28960
rect 39724 28908 39730 28960
rect 43438 28908 43444 28960
rect 43496 28948 43502 28960
rect 43717 28951 43775 28957
rect 43717 28948 43729 28951
rect 43496 28920 43729 28948
rect 43496 28908 43502 28920
rect 43717 28917 43729 28920
rect 43763 28917 43775 28951
rect 43717 28911 43775 28917
rect 1104 28858 58880 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 58880 28858
rect 1104 28784 58880 28806
rect 26510 28704 26516 28756
rect 26568 28744 26574 28756
rect 27341 28747 27399 28753
rect 27341 28744 27353 28747
rect 26568 28716 27353 28744
rect 26568 28704 26574 28716
rect 27341 28713 27353 28716
rect 27387 28713 27399 28747
rect 27341 28707 27399 28713
rect 25593 28611 25651 28617
rect 25593 28577 25605 28611
rect 25639 28608 25651 28611
rect 25866 28608 25872 28620
rect 25639 28580 25872 28608
rect 25639 28577 25651 28580
rect 25593 28571 25651 28577
rect 25866 28568 25872 28580
rect 25924 28568 25930 28620
rect 27356 28540 27384 28707
rect 28810 28704 28816 28756
rect 28868 28704 28874 28756
rect 30650 28704 30656 28756
rect 30708 28704 30714 28756
rect 31846 28704 31852 28756
rect 31904 28744 31910 28756
rect 32309 28747 32367 28753
rect 32309 28744 32321 28747
rect 31904 28716 32321 28744
rect 31904 28704 31910 28716
rect 32309 28713 32321 28716
rect 32355 28713 32367 28747
rect 32309 28707 32367 28713
rect 32398 28704 32404 28756
rect 32456 28744 32462 28756
rect 32493 28747 32551 28753
rect 32493 28744 32505 28747
rect 32456 28716 32505 28744
rect 32456 28704 32462 28716
rect 32493 28713 32505 28716
rect 32539 28713 32551 28747
rect 32493 28707 32551 28713
rect 32677 28747 32735 28753
rect 32677 28713 32689 28747
rect 32723 28744 32735 28747
rect 33778 28744 33784 28756
rect 32723 28716 33784 28744
rect 32723 28713 32735 28716
rect 32677 28707 32735 28713
rect 33778 28704 33784 28716
rect 33836 28704 33842 28756
rect 38010 28704 38016 28756
rect 38068 28704 38074 28756
rect 38194 28704 38200 28756
rect 38252 28744 38258 28756
rect 38565 28747 38623 28753
rect 38565 28744 38577 28747
rect 38252 28716 38577 28744
rect 38252 28704 38258 28716
rect 38565 28713 38577 28716
rect 38611 28713 38623 28747
rect 38565 28707 38623 28713
rect 42426 28704 42432 28756
rect 42484 28744 42490 28756
rect 42981 28747 43039 28753
rect 42981 28744 42993 28747
rect 42484 28716 42993 28744
rect 42484 28704 42490 28716
rect 42981 28713 42993 28716
rect 43027 28713 43039 28747
rect 42981 28707 43039 28713
rect 43070 28704 43076 28756
rect 43128 28744 43134 28756
rect 43717 28747 43775 28753
rect 43717 28744 43729 28747
rect 43128 28716 43729 28744
rect 43128 28704 43134 28716
rect 43717 28713 43729 28716
rect 43763 28713 43775 28747
rect 43717 28707 43775 28713
rect 44177 28747 44235 28753
rect 44177 28713 44189 28747
rect 44223 28744 44235 28747
rect 45186 28744 45192 28756
rect 44223 28716 45192 28744
rect 44223 28713 44235 28716
rect 44177 28707 44235 28713
rect 40586 28636 40592 28688
rect 40644 28676 40650 28688
rect 41322 28676 41328 28688
rect 40644 28648 41328 28676
rect 40644 28636 40650 28648
rect 41322 28636 41328 28648
rect 41380 28636 41386 28688
rect 43162 28636 43168 28688
rect 43220 28676 43226 28688
rect 44192 28676 44220 28707
rect 45186 28704 45192 28716
rect 45244 28704 45250 28756
rect 45741 28747 45799 28753
rect 45741 28713 45753 28747
rect 45787 28744 45799 28747
rect 46106 28744 46112 28756
rect 45787 28716 46112 28744
rect 45787 28713 45799 28716
rect 45741 28707 45799 28713
rect 46106 28704 46112 28716
rect 46164 28704 46170 28756
rect 43220 28648 44220 28676
rect 43220 28636 43226 28648
rect 44358 28636 44364 28688
rect 44416 28676 44422 28688
rect 44453 28679 44511 28685
rect 44453 28676 44465 28679
rect 44416 28648 44465 28676
rect 44416 28636 44422 28648
rect 44453 28645 44465 28648
rect 44499 28676 44511 28679
rect 44818 28676 44824 28688
rect 44499 28648 44824 28676
rect 44499 28645 44511 28648
rect 44453 28639 44511 28645
rect 44818 28636 44824 28648
rect 44876 28636 44882 28688
rect 29288 28580 30236 28608
rect 29288 28552 29316 28580
rect 29181 28543 29239 28549
rect 29181 28540 29193 28543
rect 27356 28512 29193 28540
rect 29181 28509 29193 28512
rect 29227 28540 29239 28543
rect 29270 28540 29276 28552
rect 29227 28512 29276 28540
rect 29227 28509 29239 28512
rect 29181 28503 29239 28509
rect 29270 28500 29276 28512
rect 29328 28500 29334 28552
rect 30208 28549 30236 28580
rect 35986 28568 35992 28620
rect 36044 28568 36050 28620
rect 42705 28611 42763 28617
rect 42705 28577 42717 28611
rect 42751 28608 42763 28611
rect 42751 28580 43300 28608
rect 42751 28577 42763 28580
rect 42705 28571 42763 28577
rect 43272 28552 43300 28580
rect 43625 28553 43683 28559
rect 30009 28543 30067 28549
rect 30009 28509 30021 28543
rect 30055 28509 30067 28543
rect 30009 28503 30067 28509
rect 30193 28543 30251 28549
rect 30193 28509 30205 28543
rect 30239 28509 30251 28543
rect 30193 28503 30251 28509
rect 25869 28475 25927 28481
rect 25869 28441 25881 28475
rect 25915 28472 25927 28475
rect 25958 28472 25964 28484
rect 25915 28444 25964 28472
rect 25915 28441 25927 28444
rect 25869 28435 25927 28441
rect 25958 28432 25964 28444
rect 26016 28432 26022 28484
rect 27430 28472 27436 28484
rect 27094 28444 27436 28472
rect 27430 28432 27436 28444
rect 27488 28432 27494 28484
rect 28997 28475 29055 28481
rect 28997 28441 29009 28475
rect 29043 28441 29055 28475
rect 30024 28472 30052 28503
rect 30466 28500 30472 28552
rect 30524 28500 30530 28552
rect 32490 28500 32496 28552
rect 32548 28540 32554 28552
rect 32677 28543 32735 28549
rect 32677 28540 32689 28543
rect 32548 28512 32689 28540
rect 32548 28500 32554 28512
rect 32677 28509 32689 28512
rect 32723 28509 32735 28543
rect 32677 28503 32735 28509
rect 32858 28500 32864 28552
rect 32916 28540 32922 28552
rect 33045 28543 33103 28549
rect 33045 28540 33057 28543
rect 32916 28512 33057 28540
rect 32916 28500 32922 28512
rect 33045 28509 33057 28512
rect 33091 28509 33103 28543
rect 33045 28503 33103 28509
rect 33134 28500 33140 28552
rect 33192 28500 33198 28552
rect 38749 28543 38807 28549
rect 38749 28509 38761 28543
rect 38795 28540 38807 28543
rect 39666 28540 39672 28552
rect 38795 28512 39672 28540
rect 38795 28509 38807 28512
rect 38749 28503 38807 28509
rect 39666 28500 39672 28512
rect 39724 28500 39730 28552
rect 40218 28500 40224 28552
rect 40276 28500 40282 28552
rect 40375 28543 40433 28549
rect 40375 28509 40387 28543
rect 40421 28540 40433 28543
rect 40494 28540 40500 28552
rect 40421 28512 40500 28540
rect 40421 28509 40433 28512
rect 40375 28503 40433 28509
rect 40494 28500 40500 28512
rect 40552 28500 40558 28552
rect 42794 28500 42800 28552
rect 42852 28500 42858 28552
rect 43162 28500 43168 28552
rect 43220 28500 43226 28552
rect 43254 28500 43260 28552
rect 43312 28500 43318 28552
rect 43438 28500 43444 28552
rect 43496 28500 43502 28552
rect 43533 28543 43591 28549
rect 43533 28509 43545 28543
rect 43579 28509 43591 28543
rect 43625 28519 43637 28553
rect 43671 28550 43683 28553
rect 43714 28550 43720 28552
rect 43671 28522 43720 28550
rect 43671 28519 43683 28522
rect 43625 28513 43683 28519
rect 43533 28503 43591 28509
rect 30558 28472 30564 28484
rect 30024 28444 30564 28472
rect 28997 28435 29055 28441
rect 29012 28404 29040 28435
rect 30558 28432 30564 28444
rect 30616 28432 30622 28484
rect 32122 28432 32128 28484
rect 32180 28432 32186 28484
rect 32325 28475 32383 28481
rect 32325 28441 32337 28475
rect 32371 28472 32383 28475
rect 32766 28472 32772 28484
rect 32371 28444 32772 28472
rect 32371 28441 32383 28444
rect 32325 28435 32383 28441
rect 32766 28432 32772 28444
rect 32824 28432 32830 28484
rect 36262 28432 36268 28484
rect 36320 28432 36326 28484
rect 38010 28472 38016 28484
rect 37490 28444 38016 28472
rect 38010 28432 38016 28444
rect 38068 28432 38074 28484
rect 38378 28432 38384 28484
rect 38436 28472 38442 28484
rect 38473 28475 38531 28481
rect 38473 28472 38485 28475
rect 38436 28444 38485 28472
rect 38436 28432 38442 28444
rect 38473 28441 38485 28444
rect 38519 28472 38531 28475
rect 38930 28472 38936 28484
rect 38519 28444 38936 28472
rect 38519 28441 38531 28444
rect 38473 28435 38531 28441
rect 38930 28432 38936 28444
rect 38988 28432 38994 28484
rect 40236 28472 40264 28500
rect 41230 28472 41236 28484
rect 40236 28444 41236 28472
rect 41230 28432 41236 28444
rect 41288 28432 41294 28484
rect 42242 28432 42248 28484
rect 42300 28472 42306 28484
rect 43548 28472 43576 28503
rect 43714 28500 43720 28522
rect 43772 28500 43778 28552
rect 43806 28500 43812 28552
rect 43864 28540 43870 28552
rect 43901 28543 43959 28549
rect 43901 28540 43913 28543
rect 43864 28512 43913 28540
rect 43864 28500 43870 28512
rect 43901 28509 43913 28512
rect 43947 28509 43959 28543
rect 43901 28503 43959 28509
rect 43990 28500 43996 28552
rect 44048 28540 44054 28552
rect 45005 28543 45063 28549
rect 45005 28540 45017 28543
rect 44048 28512 45017 28540
rect 44048 28500 44054 28512
rect 45005 28509 45017 28512
rect 45051 28509 45063 28543
rect 45005 28503 45063 28509
rect 45186 28500 45192 28552
rect 45244 28500 45250 28552
rect 45278 28500 45284 28552
rect 45336 28500 45342 28552
rect 45646 28500 45652 28552
rect 45704 28500 45710 28552
rect 50614 28500 50620 28552
rect 50672 28540 50678 28552
rect 50893 28543 50951 28549
rect 50893 28540 50905 28543
rect 50672 28512 50905 28540
rect 50672 28500 50678 28512
rect 50893 28509 50905 28512
rect 50939 28509 50951 28543
rect 50893 28503 50951 28509
rect 44174 28472 44180 28484
rect 42300 28444 44180 28472
rect 42300 28432 42306 28444
rect 43916 28416 43944 28444
rect 44174 28432 44180 28444
rect 44232 28432 44238 28484
rect 44726 28432 44732 28484
rect 44784 28432 44790 28484
rect 30006 28404 30012 28416
rect 29012 28376 30012 28404
rect 30006 28364 30012 28376
rect 30064 28404 30070 28416
rect 30285 28407 30343 28413
rect 30285 28404 30297 28407
rect 30064 28376 30297 28404
rect 30064 28364 30070 28376
rect 30285 28373 30297 28376
rect 30331 28373 30343 28407
rect 30285 28367 30343 28373
rect 37734 28364 37740 28416
rect 37792 28364 37798 28416
rect 43898 28364 43904 28416
rect 43956 28364 43962 28416
rect 44266 28364 44272 28416
rect 44324 28364 44330 28416
rect 49878 28364 49884 28416
rect 49936 28404 49942 28416
rect 50341 28407 50399 28413
rect 50341 28404 50353 28407
rect 49936 28376 50353 28404
rect 49936 28364 49942 28376
rect 50341 28373 50353 28376
rect 50387 28373 50399 28407
rect 50341 28367 50399 28373
rect 1104 28314 58880 28336
rect 1104 28262 4874 28314
rect 4926 28262 4938 28314
rect 4990 28262 5002 28314
rect 5054 28262 5066 28314
rect 5118 28262 5130 28314
rect 5182 28262 35594 28314
rect 35646 28262 35658 28314
rect 35710 28262 35722 28314
rect 35774 28262 35786 28314
rect 35838 28262 35850 28314
rect 35902 28262 58880 28314
rect 1104 28240 58880 28262
rect 27430 28160 27436 28212
rect 27488 28200 27494 28212
rect 27488 28172 28764 28200
rect 27488 28160 27494 28172
rect 28537 28135 28595 28141
rect 28537 28101 28549 28135
rect 28583 28132 28595 28135
rect 28626 28132 28632 28144
rect 28583 28104 28632 28132
rect 28583 28101 28595 28104
rect 28537 28095 28595 28101
rect 28626 28092 28632 28104
rect 28684 28092 28690 28144
rect 28736 28132 28764 28172
rect 30006 28160 30012 28212
rect 30064 28160 30070 28212
rect 36262 28160 36268 28212
rect 36320 28200 36326 28212
rect 37277 28203 37335 28209
rect 37277 28200 37289 28203
rect 36320 28172 37289 28200
rect 36320 28160 36326 28172
rect 37277 28169 37289 28172
rect 37323 28169 37335 28203
rect 37277 28163 37335 28169
rect 41230 28160 41236 28212
rect 41288 28200 41294 28212
rect 42702 28200 42708 28212
rect 41288 28172 42708 28200
rect 41288 28160 41294 28172
rect 42702 28160 42708 28172
rect 42760 28200 42766 28212
rect 43714 28200 43720 28212
rect 42760 28172 43720 28200
rect 42760 28160 42766 28172
rect 43714 28160 43720 28172
rect 43772 28160 43778 28212
rect 44174 28160 44180 28212
rect 44232 28200 44238 28212
rect 44232 28172 44588 28200
rect 44232 28160 44238 28172
rect 28736 28104 29026 28132
rect 36538 28092 36544 28144
rect 36596 28132 36602 28144
rect 37001 28135 37059 28141
rect 37001 28132 37013 28135
rect 36596 28104 37013 28132
rect 36596 28092 36602 28104
rect 37001 28101 37013 28104
rect 37047 28132 37059 28135
rect 37826 28132 37832 28144
rect 37047 28104 37832 28132
rect 37047 28101 37059 28104
rect 37001 28095 37059 28101
rect 37826 28092 37832 28104
rect 37884 28092 37890 28144
rect 40034 28092 40040 28144
rect 40092 28132 40098 28144
rect 40129 28135 40187 28141
rect 40129 28132 40141 28135
rect 40092 28104 40141 28132
rect 40092 28092 40098 28104
rect 40129 28101 40141 28104
rect 40175 28101 40187 28135
rect 44560 28132 44588 28172
rect 44910 28160 44916 28212
rect 44968 28200 44974 28212
rect 46845 28203 46903 28209
rect 46845 28200 46857 28203
rect 44968 28172 46857 28200
rect 44968 28160 44974 28172
rect 46845 28169 46857 28172
rect 46891 28200 46903 28203
rect 47765 28203 47823 28209
rect 47765 28200 47777 28203
rect 46891 28172 47777 28200
rect 46891 28169 46903 28172
rect 46845 28163 46903 28169
rect 47765 28169 47777 28172
rect 47811 28169 47823 28203
rect 47765 28163 47823 28169
rect 45189 28135 45247 28141
rect 45189 28132 45201 28135
rect 40129 28095 40187 28101
rect 43088 28104 44496 28132
rect 44560 28104 45201 28132
rect 43088 28076 43116 28104
rect 37645 28067 37703 28073
rect 37645 28033 37657 28067
rect 37691 28064 37703 28067
rect 38930 28064 38936 28076
rect 37691 28036 38936 28064
rect 37691 28033 37703 28036
rect 37645 28027 37703 28033
rect 38930 28024 38936 28036
rect 38988 28024 38994 28076
rect 42242 28024 42248 28076
rect 42300 28024 42306 28076
rect 42702 28024 42708 28076
rect 42760 28024 42766 28076
rect 42794 28024 42800 28076
rect 42852 28024 42858 28076
rect 42886 28024 42892 28076
rect 42944 28064 42950 28076
rect 42981 28067 43039 28073
rect 42981 28064 42993 28067
rect 42944 28036 42993 28064
rect 42944 28024 42950 28036
rect 42981 28033 42993 28036
rect 43027 28033 43039 28067
rect 42981 28027 43039 28033
rect 43070 28024 43076 28076
rect 43128 28024 43134 28076
rect 43717 28067 43775 28073
rect 43717 28033 43729 28067
rect 43763 28064 43775 28067
rect 43990 28064 43996 28076
rect 43763 28036 43996 28064
rect 43763 28033 43775 28036
rect 43717 28027 43775 28033
rect 43990 28024 43996 28036
rect 44048 28024 44054 28076
rect 44085 28067 44143 28073
rect 44085 28033 44097 28067
rect 44131 28064 44143 28067
rect 44468 28064 44496 28104
rect 45189 28101 45201 28104
rect 45235 28132 45247 28135
rect 46937 28135 46995 28141
rect 46937 28132 46949 28135
rect 45235 28104 46949 28132
rect 45235 28101 45247 28104
rect 45189 28095 45247 28101
rect 46937 28101 46949 28104
rect 46983 28132 46995 28135
rect 48130 28132 48136 28144
rect 46983 28104 48136 28132
rect 46983 28101 46995 28104
rect 46937 28095 46995 28101
rect 48130 28092 48136 28104
rect 48188 28092 48194 28144
rect 49694 28092 49700 28144
rect 49752 28132 49758 28144
rect 50985 28135 51043 28141
rect 50985 28132 50997 28135
rect 49752 28104 50997 28132
rect 49752 28092 49758 28104
rect 50985 28101 50997 28104
rect 51031 28101 51043 28135
rect 50985 28095 51043 28101
rect 44545 28067 44603 28073
rect 44545 28064 44557 28067
rect 44131 28036 44404 28064
rect 44468 28036 44557 28064
rect 44131 28033 44143 28036
rect 44085 28027 44143 28033
rect 28258 27956 28264 28008
rect 28316 27956 28322 28008
rect 37734 27956 37740 28008
rect 37792 27956 37798 28008
rect 37826 27956 37832 28008
rect 37884 27956 37890 28008
rect 41782 27956 41788 28008
rect 41840 27996 41846 28008
rect 44376 28005 44404 28036
rect 44545 28033 44557 28036
rect 44591 28064 44603 28067
rect 45005 28067 45063 28073
rect 45005 28064 45017 28067
rect 44591 28036 45017 28064
rect 44591 28033 44603 28036
rect 44545 28027 44603 28033
rect 45005 28033 45017 28036
rect 45051 28033 45063 28067
rect 45005 28027 45063 28033
rect 47578 28024 47584 28076
rect 47636 28024 47642 28076
rect 49602 28024 49608 28076
rect 49660 28024 49666 28076
rect 49878 28024 49884 28076
rect 49936 28024 49942 28076
rect 50062 28024 50068 28076
rect 50120 28064 50126 28076
rect 50249 28067 50307 28073
rect 50249 28064 50261 28067
rect 50120 28036 50261 28064
rect 50120 28024 50126 28036
rect 50249 28033 50261 28036
rect 50295 28033 50307 28067
rect 50249 28027 50307 28033
rect 42153 27999 42211 28005
rect 42153 27996 42165 27999
rect 41840 27968 42165 27996
rect 41840 27956 41846 27968
rect 42153 27965 42165 27968
rect 42199 27996 42211 27999
rect 43257 27999 43315 28005
rect 43257 27996 43269 27999
rect 42199 27968 43269 27996
rect 42199 27965 42211 27968
rect 42153 27959 42211 27965
rect 43257 27965 43269 27968
rect 43303 27965 43315 27999
rect 43257 27959 43315 27965
rect 44361 27999 44419 28005
rect 44361 27965 44373 27999
rect 44407 27965 44419 27999
rect 44361 27959 44419 27965
rect 44634 27956 44640 28008
rect 44692 27956 44698 28008
rect 44726 27956 44732 28008
rect 44784 27956 44790 28008
rect 44818 27956 44824 28008
rect 44876 27956 44882 28008
rect 47121 27999 47179 28005
rect 47121 27965 47133 27999
rect 47167 27996 47179 27999
rect 50890 27996 50896 28008
rect 47167 27968 50896 27996
rect 47167 27965 47179 27968
rect 47121 27959 47179 27965
rect 37752 27928 37780 27956
rect 40494 27928 40500 27940
rect 37752 27900 40500 27928
rect 40494 27888 40500 27900
rect 40552 27928 40558 27940
rect 42978 27928 42984 27940
rect 40552 27900 42984 27928
rect 40552 27888 40558 27900
rect 42978 27888 42984 27900
rect 43036 27888 43042 27940
rect 44085 27931 44143 27937
rect 44085 27928 44097 27931
rect 43088 27900 44097 27928
rect 40589 27863 40647 27869
rect 40589 27829 40601 27863
rect 40635 27860 40647 27863
rect 40954 27860 40960 27872
rect 40635 27832 40960 27860
rect 40635 27829 40647 27832
rect 40589 27823 40647 27829
rect 40954 27820 40960 27832
rect 41012 27820 41018 27872
rect 42521 27863 42579 27869
rect 42521 27829 42533 27863
rect 42567 27860 42579 27863
rect 42610 27860 42616 27872
rect 42567 27832 42616 27860
rect 42567 27829 42579 27832
rect 42521 27823 42579 27829
rect 42610 27820 42616 27832
rect 42668 27820 42674 27872
rect 42702 27820 42708 27872
rect 42760 27860 42766 27872
rect 43088 27860 43116 27900
rect 44085 27897 44097 27900
rect 44131 27928 44143 27931
rect 45646 27928 45652 27940
rect 44131 27900 45652 27928
rect 44131 27897 44143 27900
rect 44085 27891 44143 27897
rect 45646 27888 45652 27900
rect 45704 27888 45710 27940
rect 45922 27888 45928 27940
rect 45980 27928 45986 27940
rect 46385 27931 46443 27937
rect 46385 27928 46397 27931
rect 45980 27900 46397 27928
rect 45980 27888 45986 27900
rect 46385 27897 46397 27900
rect 46431 27928 46443 27931
rect 47136 27928 47164 27959
rect 50890 27956 50896 27968
rect 50948 27956 50954 28008
rect 46431 27900 47164 27928
rect 46431 27897 46443 27900
rect 46385 27891 46443 27897
rect 42760 27832 43116 27860
rect 42760 27820 42766 27832
rect 43622 27820 43628 27872
rect 43680 27860 43686 27872
rect 45373 27863 45431 27869
rect 45373 27860 45385 27863
rect 43680 27832 45385 27860
rect 43680 27820 43686 27832
rect 45373 27829 45385 27832
rect 45419 27829 45431 27863
rect 45373 27823 45431 27829
rect 46474 27820 46480 27872
rect 46532 27820 46538 27872
rect 49418 27820 49424 27872
rect 49476 27820 49482 27872
rect 49786 27820 49792 27872
rect 49844 27820 49850 27872
rect 50062 27820 50068 27872
rect 50120 27820 50126 27872
rect 1104 27770 58880 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 58880 27770
rect 1104 27696 58880 27718
rect 37908 27659 37966 27665
rect 37908 27625 37920 27659
rect 37954 27656 37966 27659
rect 37954 27628 39896 27656
rect 37954 27625 37966 27628
rect 37908 27619 37966 27625
rect 39868 27597 39896 27628
rect 43070 27616 43076 27668
rect 43128 27616 43134 27668
rect 43257 27659 43315 27665
rect 43257 27656 43269 27659
rect 43180 27628 43269 27656
rect 39853 27591 39911 27597
rect 39853 27557 39865 27591
rect 39899 27557 39911 27591
rect 39853 27551 39911 27557
rect 40954 27548 40960 27600
rect 41012 27548 41018 27600
rect 42886 27548 42892 27600
rect 42944 27588 42950 27600
rect 43180 27588 43208 27628
rect 43257 27625 43269 27628
rect 43303 27625 43315 27659
rect 43257 27619 43315 27625
rect 43622 27616 43628 27668
rect 43680 27616 43686 27668
rect 43898 27616 43904 27668
rect 43956 27656 43962 27668
rect 43993 27659 44051 27665
rect 43993 27656 44005 27659
rect 43956 27628 44005 27656
rect 43956 27616 43962 27628
rect 43993 27625 44005 27628
rect 44039 27625 44051 27659
rect 44266 27656 44272 27668
rect 43993 27619 44051 27625
rect 44100 27628 44272 27656
rect 44100 27588 44128 27628
rect 44266 27616 44272 27628
rect 44324 27616 44330 27668
rect 44637 27659 44695 27665
rect 44637 27625 44649 27659
rect 44683 27656 44695 27659
rect 44726 27656 44732 27668
rect 44683 27628 44732 27656
rect 44683 27625 44695 27628
rect 44637 27619 44695 27625
rect 44652 27588 44680 27619
rect 44726 27616 44732 27628
rect 44784 27616 44790 27668
rect 46474 27616 46480 27668
rect 46532 27656 46538 27668
rect 46642 27659 46700 27665
rect 46642 27656 46654 27659
rect 46532 27628 46654 27656
rect 46532 27616 46538 27628
rect 46642 27625 46654 27628
rect 46688 27625 46700 27659
rect 46642 27619 46700 27625
rect 47394 27616 47400 27668
rect 47452 27656 47458 27668
rect 47452 27628 47716 27656
rect 47452 27616 47458 27628
rect 42944 27560 43208 27588
rect 43364 27560 44128 27588
rect 44284 27560 44680 27588
rect 47688 27588 47716 27628
rect 48130 27616 48136 27668
rect 48188 27616 48194 27668
rect 52454 27656 52460 27668
rect 48332 27628 52460 27656
rect 48332 27597 48360 27628
rect 52454 27616 52460 27628
rect 52512 27616 52518 27668
rect 48317 27591 48375 27597
rect 48317 27588 48329 27591
rect 47688 27560 48329 27588
rect 42944 27548 42950 27560
rect 32493 27523 32551 27529
rect 32493 27520 32505 27523
rect 30576 27492 32505 27520
rect 30576 27464 30604 27492
rect 32493 27489 32505 27492
rect 32539 27520 32551 27523
rect 34701 27523 34759 27529
rect 34701 27520 34713 27523
rect 32539 27492 34713 27520
rect 32539 27489 32551 27492
rect 32493 27483 32551 27489
rect 34701 27489 34713 27492
rect 34747 27489 34759 27523
rect 34701 27483 34759 27489
rect 40494 27480 40500 27532
rect 40552 27480 40558 27532
rect 41598 27480 41604 27532
rect 41656 27520 41662 27532
rect 43364 27520 43392 27560
rect 41656 27492 43392 27520
rect 41656 27480 41662 27492
rect 30377 27455 30435 27461
rect 30377 27421 30389 27455
rect 30423 27452 30435 27455
rect 30558 27452 30564 27464
rect 30423 27424 30564 27452
rect 30423 27421 30435 27424
rect 30377 27415 30435 27421
rect 30558 27412 30564 27424
rect 30616 27412 30622 27464
rect 30926 27412 30932 27464
rect 30984 27412 30990 27464
rect 32766 27412 32772 27464
rect 32824 27452 32830 27464
rect 32861 27455 32919 27461
rect 32861 27452 32873 27455
rect 32824 27424 32873 27452
rect 32824 27412 32830 27424
rect 32861 27421 32873 27424
rect 32907 27421 32919 27455
rect 35069 27455 35127 27461
rect 35069 27452 35081 27455
rect 32861 27415 32919 27421
rect 34716 27424 35081 27452
rect 34716 27396 34744 27424
rect 35069 27421 35081 27424
rect 35115 27421 35127 27455
rect 35069 27415 35127 27421
rect 37642 27412 37648 27464
rect 37700 27412 37706 27464
rect 41233 27455 41291 27461
rect 41233 27421 41245 27455
rect 41279 27452 41291 27455
rect 41414 27452 41420 27464
rect 41279 27424 41420 27452
rect 41279 27421 41291 27424
rect 41233 27415 41291 27421
rect 41414 27412 41420 27424
rect 41472 27412 41478 27464
rect 41509 27455 41567 27461
rect 41509 27421 41521 27455
rect 41555 27452 41567 27455
rect 42521 27455 42579 27461
rect 42521 27452 42533 27455
rect 41555 27424 42533 27452
rect 41555 27421 41567 27424
rect 41509 27415 41567 27421
rect 42521 27421 42533 27424
rect 42567 27421 42579 27455
rect 42521 27415 42579 27421
rect 42613 27455 42671 27461
rect 42613 27421 42625 27455
rect 42659 27421 42671 27455
rect 42613 27415 42671 27421
rect 29365 27387 29423 27393
rect 29365 27353 29377 27387
rect 29411 27384 29423 27387
rect 29546 27384 29552 27396
rect 29411 27356 29552 27384
rect 29411 27353 29423 27356
rect 29365 27347 29423 27353
rect 29546 27344 29552 27356
rect 29604 27344 29610 27396
rect 32214 27384 32220 27396
rect 31970 27356 32220 27384
rect 32214 27344 32220 27356
rect 32272 27384 32278 27396
rect 32272 27356 32628 27384
rect 32272 27344 32278 27356
rect 32355 27319 32413 27325
rect 32355 27285 32367 27319
rect 32401 27316 32413 27319
rect 32490 27316 32496 27328
rect 32401 27288 32496 27316
rect 32401 27285 32413 27288
rect 32355 27279 32413 27285
rect 32490 27276 32496 27288
rect 32548 27276 32554 27328
rect 32600 27316 32628 27356
rect 33152 27356 33258 27384
rect 33152 27316 33180 27356
rect 34698 27344 34704 27396
rect 34756 27344 34762 27396
rect 36262 27384 36268 27396
rect 36110 27356 36268 27384
rect 36262 27344 36268 27356
rect 36320 27384 36326 27396
rect 39669 27387 39727 27393
rect 36320 27356 38410 27384
rect 36320 27344 36326 27356
rect 39669 27353 39681 27387
rect 39715 27384 39727 27387
rect 39715 27356 40356 27384
rect 39715 27353 39727 27356
rect 39669 27347 39727 27353
rect 32600 27288 33180 27316
rect 33318 27276 33324 27328
rect 33376 27316 33382 27328
rect 34287 27319 34345 27325
rect 34287 27316 34299 27319
rect 33376 27288 34299 27316
rect 33376 27276 33382 27288
rect 34287 27285 34299 27288
rect 34333 27316 34345 27319
rect 34514 27316 34520 27328
rect 34333 27288 34520 27316
rect 34333 27285 34345 27288
rect 34287 27279 34345 27285
rect 34514 27276 34520 27288
rect 34572 27276 34578 27328
rect 36495 27319 36553 27325
rect 36495 27285 36507 27319
rect 36541 27316 36553 27319
rect 36722 27316 36728 27328
rect 36541 27288 36728 27316
rect 36541 27285 36553 27288
rect 36495 27279 36553 27285
rect 36722 27276 36728 27288
rect 36780 27276 36786 27328
rect 39942 27276 39948 27328
rect 40000 27316 40006 27328
rect 40328 27325 40356 27356
rect 40402 27344 40408 27396
rect 40460 27384 40466 27396
rect 41049 27387 41107 27393
rect 41049 27384 41061 27387
rect 40460 27356 41061 27384
rect 40460 27344 40466 27356
rect 41049 27353 41061 27356
rect 41095 27353 41107 27387
rect 41049 27347 41107 27353
rect 41782 27344 41788 27396
rect 41840 27344 41846 27396
rect 42628 27384 42656 27415
rect 42794 27412 42800 27464
rect 42852 27452 42858 27464
rect 42889 27455 42947 27461
rect 42889 27452 42901 27455
rect 42852 27424 42901 27452
rect 42852 27412 42858 27424
rect 42889 27421 42901 27424
rect 42935 27421 42947 27455
rect 42889 27415 42947 27421
rect 42978 27412 42984 27464
rect 43036 27452 43042 27464
rect 43073 27455 43131 27461
rect 43073 27452 43085 27455
rect 43036 27424 43085 27452
rect 43036 27412 43042 27424
rect 43073 27421 43085 27424
rect 43119 27421 43131 27455
rect 43073 27415 43131 27421
rect 43162 27412 43168 27464
rect 43220 27412 43226 27464
rect 43364 27461 43392 27492
rect 43530 27480 43536 27532
rect 43588 27480 43594 27532
rect 43714 27480 43720 27532
rect 43772 27480 43778 27532
rect 44082 27480 44088 27532
rect 44140 27520 44146 27532
rect 44177 27523 44235 27529
rect 44177 27520 44189 27523
rect 44140 27492 44189 27520
rect 44140 27480 44146 27492
rect 44177 27489 44189 27492
rect 44223 27489 44235 27523
rect 44177 27483 44235 27489
rect 43349 27455 43407 27461
rect 43349 27421 43361 27455
rect 43395 27421 43407 27455
rect 43349 27415 43407 27421
rect 43441 27387 43499 27393
rect 43441 27384 43453 27387
rect 42628 27356 43453 27384
rect 43441 27353 43453 27356
rect 43487 27384 43499 27387
rect 43548 27384 43576 27480
rect 43732 27452 43760 27480
rect 44284 27461 44312 27560
rect 48317 27557 48329 27560
rect 48363 27557 48375 27591
rect 48317 27551 48375 27557
rect 48222 27480 48228 27532
rect 48280 27520 48286 27532
rect 49786 27520 49792 27532
rect 48280 27492 49792 27520
rect 48280 27480 48286 27492
rect 49786 27480 49792 27492
rect 49844 27520 49850 27532
rect 50982 27520 50988 27532
rect 49844 27492 50988 27520
rect 49844 27480 49850 27492
rect 50982 27480 50988 27492
rect 51040 27480 51046 27532
rect 51902 27480 51908 27532
rect 51960 27520 51966 27532
rect 52549 27523 52607 27529
rect 52549 27520 52561 27523
rect 51960 27492 52561 27520
rect 51960 27480 51966 27492
rect 52549 27489 52561 27492
rect 52595 27489 52607 27523
rect 52549 27483 52607 27489
rect 44269 27455 44327 27461
rect 43732 27424 44128 27452
rect 43487 27356 43576 27384
rect 43657 27387 43715 27393
rect 43487 27353 43499 27356
rect 43441 27347 43499 27353
rect 43657 27353 43669 27387
rect 43703 27384 43715 27387
rect 43990 27384 43996 27396
rect 43703 27356 43996 27384
rect 43703 27353 43715 27356
rect 43657 27347 43715 27353
rect 43990 27344 43996 27356
rect 44048 27344 44054 27396
rect 44100 27384 44128 27424
rect 44269 27421 44281 27455
rect 44315 27421 44327 27455
rect 44269 27415 44327 27421
rect 44545 27455 44603 27461
rect 44545 27421 44557 27455
rect 44591 27421 44603 27455
rect 44545 27415 44603 27421
rect 44560 27384 44588 27415
rect 46290 27412 46296 27464
rect 46348 27452 46354 27464
rect 46385 27455 46443 27461
rect 46385 27452 46397 27455
rect 46348 27424 46397 27452
rect 46348 27412 46354 27424
rect 46385 27421 46397 27424
rect 46431 27421 46443 27455
rect 46385 27415 46443 27421
rect 49694 27412 49700 27464
rect 49752 27452 49758 27464
rect 50157 27455 50215 27461
rect 50157 27452 50169 27455
rect 49752 27424 50169 27452
rect 49752 27412 49758 27424
rect 50157 27421 50169 27424
rect 50203 27421 50215 27455
rect 50157 27415 50215 27421
rect 44100 27356 44588 27384
rect 47394 27344 47400 27396
rect 47452 27344 47458 27396
rect 50430 27344 50436 27396
rect 50488 27344 50494 27396
rect 50522 27344 50528 27396
rect 50580 27384 50586 27396
rect 50580 27356 50922 27384
rect 50580 27344 50586 27356
rect 40221 27319 40279 27325
rect 40221 27316 40233 27319
rect 40000 27288 40233 27316
rect 40000 27276 40006 27288
rect 40221 27285 40233 27288
rect 40267 27285 40279 27319
rect 40221 27279 40279 27285
rect 40313 27319 40371 27325
rect 40313 27285 40325 27319
rect 40359 27316 40371 27319
rect 41230 27316 41236 27328
rect 40359 27288 41236 27316
rect 40359 27285 40371 27288
rect 40313 27279 40371 27285
rect 41230 27276 41236 27288
rect 41288 27276 41294 27328
rect 43809 27319 43867 27325
rect 43809 27285 43821 27319
rect 43855 27316 43867 27319
rect 45094 27316 45100 27328
rect 43855 27288 45100 27316
rect 43855 27285 43867 27288
rect 43809 27279 43867 27285
rect 45094 27276 45100 27288
rect 45152 27316 45158 27328
rect 47578 27316 47584 27328
rect 45152 27288 47584 27316
rect 45152 27276 45158 27288
rect 47578 27276 47584 27288
rect 47636 27276 47642 27328
rect 51994 27276 52000 27328
rect 52052 27276 52058 27328
rect 1104 27226 58880 27248
rect 1104 27174 4874 27226
rect 4926 27174 4938 27226
rect 4990 27174 5002 27226
rect 5054 27174 5066 27226
rect 5118 27174 5130 27226
rect 5182 27174 35594 27226
rect 35646 27174 35658 27226
rect 35710 27174 35722 27226
rect 35774 27174 35786 27226
rect 35838 27174 35850 27226
rect 35902 27174 58880 27226
rect 1104 27152 58880 27174
rect 28902 27112 28908 27124
rect 25700 27084 28908 27112
rect 25700 27044 25728 27084
rect 28000 27044 28028 27084
rect 28902 27072 28908 27084
rect 28960 27072 28966 27124
rect 30926 27072 30932 27124
rect 30984 27112 30990 27124
rect 32125 27115 32183 27121
rect 32125 27112 32137 27115
rect 30984 27084 32137 27112
rect 30984 27072 30990 27084
rect 32125 27081 32137 27084
rect 32171 27081 32183 27115
rect 32125 27075 32183 27081
rect 32766 27072 32772 27124
rect 32824 27072 32830 27124
rect 33413 27115 33471 27121
rect 33413 27112 33425 27115
rect 33060 27084 33425 27112
rect 24702 27016 25806 27044
rect 28000 27016 28106 27044
rect 32030 26936 32036 26988
rect 32088 26976 32094 26988
rect 32309 26979 32367 26985
rect 32309 26976 32321 26979
rect 32088 26948 32321 26976
rect 32088 26936 32094 26948
rect 32309 26945 32321 26948
rect 32355 26945 32367 26979
rect 32309 26939 32367 26945
rect 32398 26936 32404 26988
rect 32456 26936 32462 26988
rect 32490 26936 32496 26988
rect 32548 26976 32554 26988
rect 32677 26979 32735 26985
rect 32677 26976 32689 26979
rect 32548 26948 32689 26976
rect 32548 26936 32554 26948
rect 32677 26945 32689 26948
rect 32723 26976 32735 26979
rect 32858 26976 32864 26988
rect 32723 26948 32864 26976
rect 32723 26945 32735 26948
rect 32677 26939 32735 26945
rect 32858 26936 32864 26948
rect 32916 26936 32922 26988
rect 32950 26936 32956 26988
rect 33008 26936 33014 26988
rect 33060 26985 33088 27084
rect 33413 27081 33425 27084
rect 33459 27081 33471 27115
rect 33413 27075 33471 27081
rect 33520 27084 34008 27112
rect 33045 26979 33103 26985
rect 33045 26945 33057 26979
rect 33091 26945 33103 26979
rect 33045 26939 33103 26945
rect 33318 26936 33324 26988
rect 33376 26936 33382 26988
rect 33520 26976 33548 27084
rect 33428 26948 33548 26976
rect 33597 26979 33655 26985
rect 22830 26868 22836 26920
rect 22888 26908 22894 26920
rect 23201 26911 23259 26917
rect 23201 26908 23213 26911
rect 22888 26880 23213 26908
rect 22888 26868 22894 26880
rect 23201 26877 23213 26880
rect 23247 26877 23259 26911
rect 23201 26871 23259 26877
rect 23474 26868 23480 26920
rect 23532 26868 23538 26920
rect 25041 26911 25099 26917
rect 25041 26877 25053 26911
rect 25087 26877 25099 26911
rect 25041 26871 25099 26877
rect 24946 26732 24952 26784
rect 25004 26732 25010 26784
rect 25056 26772 25084 26871
rect 25314 26868 25320 26920
rect 25372 26868 25378 26920
rect 25866 26868 25872 26920
rect 25924 26908 25930 26920
rect 27341 26911 27399 26917
rect 27341 26908 27353 26911
rect 25924 26880 27353 26908
rect 25924 26868 25930 26880
rect 27341 26877 27353 26880
rect 27387 26908 27399 26911
rect 27387 26880 27476 26908
rect 27387 26877 27399 26880
rect 27341 26871 27399 26877
rect 25866 26772 25872 26784
rect 25056 26744 25872 26772
rect 25866 26732 25872 26744
rect 25924 26732 25930 26784
rect 26786 26732 26792 26784
rect 26844 26732 26850 26784
rect 27448 26772 27476 26880
rect 27614 26868 27620 26920
rect 27672 26868 27678 26920
rect 32876 26908 32904 26936
rect 33428 26908 33456 26948
rect 33597 26945 33609 26979
rect 33643 26945 33655 26979
rect 33597 26939 33655 26945
rect 32876 26880 33456 26908
rect 33612 26840 33640 26939
rect 33686 26936 33692 26988
rect 33744 26936 33750 26988
rect 33980 26985 34008 27084
rect 34514 27072 34520 27124
rect 34572 27112 34578 27124
rect 35986 27112 35992 27124
rect 34572 27084 35992 27112
rect 34572 27072 34578 27084
rect 35986 27072 35992 27084
rect 36044 27072 36050 27124
rect 36538 27112 36544 27124
rect 36372 27084 36544 27112
rect 34532 26985 34560 27072
rect 36262 27004 36268 27056
rect 36320 27044 36326 27056
rect 36372 27044 36400 27084
rect 36538 27072 36544 27084
rect 36596 27072 36602 27124
rect 37826 27072 37832 27124
rect 37884 27112 37890 27124
rect 37884 27084 38654 27112
rect 37884 27072 37890 27084
rect 36320 27016 36400 27044
rect 36320 27004 36326 27016
rect 33781 26979 33839 26985
rect 33781 26945 33793 26979
rect 33827 26945 33839 26979
rect 33781 26939 33839 26945
rect 33945 26979 34008 26985
rect 33945 26945 33957 26979
rect 33991 26948 34008 26979
rect 34517 26979 34575 26985
rect 33991 26945 34003 26948
rect 33945 26939 34003 26945
rect 34517 26945 34529 26979
rect 34563 26945 34575 26979
rect 34517 26939 34575 26945
rect 34701 26979 34759 26985
rect 34701 26945 34713 26979
rect 34747 26945 34759 26979
rect 34701 26939 34759 26945
rect 34793 26979 34851 26985
rect 34793 26945 34805 26979
rect 34839 26945 34851 26979
rect 34793 26939 34851 26945
rect 33796 26908 33824 26939
rect 34606 26908 34612 26920
rect 33796 26880 34612 26908
rect 34606 26868 34612 26880
rect 34664 26908 34670 26920
rect 34716 26908 34744 26939
rect 34664 26880 34744 26908
rect 34808 26908 34836 26939
rect 34882 26936 34888 26988
rect 34940 26936 34946 26988
rect 37001 26979 37059 26985
rect 37001 26945 37013 26979
rect 37047 26976 37059 26979
rect 37642 26976 37648 26988
rect 37047 26948 37648 26976
rect 37047 26945 37059 26948
rect 37001 26939 37059 26945
rect 34808 26880 35250 26908
rect 34664 26868 34670 26880
rect 34514 26840 34520 26852
rect 33612 26812 34520 26840
rect 34514 26800 34520 26812
rect 34572 26840 34578 26852
rect 34882 26840 34888 26852
rect 34572 26812 34888 26840
rect 34572 26800 34578 26812
rect 34882 26800 34888 26812
rect 34940 26800 34946 26852
rect 28350 26772 28356 26784
rect 27448 26744 28356 26772
rect 28350 26732 28356 26744
rect 28408 26732 28414 26784
rect 28626 26732 28632 26784
rect 28684 26772 28690 26784
rect 29089 26775 29147 26781
rect 29089 26772 29101 26775
rect 28684 26744 29101 26772
rect 28684 26732 28690 26744
rect 29089 26741 29101 26744
rect 29135 26741 29147 26775
rect 29089 26735 29147 26741
rect 32585 26775 32643 26781
rect 32585 26741 32597 26775
rect 32631 26772 32643 26775
rect 32858 26772 32864 26784
rect 32631 26744 32864 26772
rect 32631 26741 32643 26744
rect 32585 26735 32643 26741
rect 32858 26732 32864 26744
rect 32916 26772 32922 26784
rect 33229 26775 33287 26781
rect 33229 26772 33241 26775
rect 32916 26744 33241 26772
rect 32916 26732 32922 26744
rect 33229 26741 33241 26744
rect 33275 26741 33287 26775
rect 33229 26735 33287 26741
rect 34790 26732 34796 26784
rect 34848 26772 34854 26784
rect 35222 26781 35250 26880
rect 36630 26868 36636 26920
rect 36688 26868 36694 26920
rect 36814 26868 36820 26920
rect 36872 26908 36878 26920
rect 37016 26908 37044 26939
rect 37642 26936 37648 26948
rect 37700 26936 37706 26988
rect 36872 26880 37044 26908
rect 36872 26868 36878 26880
rect 35069 26775 35127 26781
rect 35069 26772 35081 26775
rect 34848 26744 35081 26772
rect 34848 26732 34854 26744
rect 35069 26741 35081 26744
rect 35115 26741 35127 26775
rect 35069 26735 35127 26741
rect 35207 26775 35265 26781
rect 35207 26741 35219 26775
rect 35253 26772 35265 26775
rect 36078 26772 36084 26784
rect 35253 26744 36084 26772
rect 35253 26741 35265 26744
rect 35207 26735 35265 26741
rect 36078 26732 36084 26744
rect 36136 26732 36142 26784
rect 38626 26772 38654 27084
rect 39942 27072 39948 27124
rect 40000 27072 40006 27124
rect 42794 27072 42800 27124
rect 42852 27112 42858 27124
rect 43441 27115 43499 27121
rect 43441 27112 43453 27115
rect 42852 27084 43453 27112
rect 42852 27072 42858 27084
rect 43441 27081 43453 27084
rect 43487 27112 43499 27115
rect 43806 27112 43812 27124
rect 43487 27084 43812 27112
rect 43487 27081 43499 27084
rect 43441 27075 43499 27081
rect 43806 27072 43812 27084
rect 43864 27072 43870 27124
rect 49878 27112 49884 27124
rect 47596 27084 49884 27112
rect 47596 27053 47624 27084
rect 49878 27072 49884 27084
rect 49936 27072 49942 27124
rect 50430 27072 50436 27124
rect 50488 27112 50494 27124
rect 50709 27115 50767 27121
rect 50709 27112 50721 27115
rect 50488 27084 50721 27112
rect 50488 27072 50494 27084
rect 50709 27081 50721 27084
rect 50755 27081 50767 27115
rect 50709 27075 50767 27081
rect 52454 27072 52460 27124
rect 52512 27072 52518 27124
rect 47581 27047 47639 27053
rect 47581 27044 47593 27047
rect 43548 27016 43944 27044
rect 40129 26979 40187 26985
rect 40129 26945 40141 26979
rect 40175 26976 40187 26979
rect 40218 26976 40224 26988
rect 40175 26948 40224 26976
rect 40175 26945 40187 26948
rect 40129 26939 40187 26945
rect 40218 26936 40224 26948
rect 40276 26976 40282 26988
rect 40957 26979 41015 26985
rect 40957 26976 40969 26979
rect 40276 26948 40969 26976
rect 40276 26936 40282 26948
rect 40957 26945 40969 26948
rect 41003 26945 41015 26979
rect 40957 26939 41015 26945
rect 41046 26936 41052 26988
rect 41104 26976 41110 26988
rect 41141 26979 41199 26985
rect 41141 26976 41153 26979
rect 41104 26948 41153 26976
rect 41104 26936 41110 26948
rect 41141 26945 41153 26948
rect 41187 26945 41199 26979
rect 41141 26939 41199 26945
rect 41230 26936 41236 26988
rect 41288 26936 41294 26988
rect 41509 26979 41567 26985
rect 41509 26945 41521 26979
rect 41555 26976 41567 26979
rect 41782 26976 41788 26988
rect 41555 26948 41788 26976
rect 41555 26945 41567 26948
rect 41509 26939 41567 26945
rect 41782 26936 41788 26948
rect 41840 26936 41846 26988
rect 43548 26985 43576 27016
rect 43916 26988 43944 27016
rect 47044 27016 47593 27044
rect 43257 26979 43315 26985
rect 43257 26945 43269 26979
rect 43303 26945 43315 26979
rect 43257 26939 43315 26945
rect 43533 26979 43591 26985
rect 43533 26945 43545 26979
rect 43579 26945 43591 26979
rect 43533 26939 43591 26945
rect 40313 26911 40371 26917
rect 40313 26877 40325 26911
rect 40359 26908 40371 26911
rect 40402 26908 40408 26920
rect 40359 26880 40408 26908
rect 40359 26877 40371 26880
rect 40313 26871 40371 26877
rect 40402 26868 40408 26880
rect 40460 26868 40466 26920
rect 41417 26911 41475 26917
rect 41417 26877 41429 26911
rect 41463 26908 41475 26911
rect 41598 26908 41604 26920
rect 41463 26880 41604 26908
rect 41463 26877 41475 26880
rect 41417 26871 41475 26877
rect 41598 26868 41604 26880
rect 41656 26868 41662 26920
rect 42334 26868 42340 26920
rect 42392 26908 42398 26920
rect 42702 26908 42708 26920
rect 42392 26880 42708 26908
rect 42392 26868 42398 26880
rect 42702 26868 42708 26880
rect 42760 26868 42766 26920
rect 43272 26908 43300 26939
rect 43622 26936 43628 26988
rect 43680 26936 43686 26988
rect 43898 26936 43904 26988
rect 43956 26936 43962 26988
rect 47044 26985 47072 27016
rect 47581 27013 47593 27016
rect 47627 27013 47639 27047
rect 47581 27007 47639 27013
rect 49145 27047 49203 27053
rect 49145 27013 49157 27047
rect 49191 27044 49203 27047
rect 49418 27044 49424 27056
rect 49191 27016 49424 27044
rect 49191 27013 49203 27016
rect 49145 27007 49203 27013
rect 49418 27004 49424 27016
rect 49476 27004 49482 27056
rect 52472 27044 52500 27072
rect 53282 27044 53288 27056
rect 52472 27016 53288 27044
rect 53282 27004 53288 27016
rect 53340 27044 53346 27056
rect 53340 27016 53498 27044
rect 53340 27004 53346 27016
rect 47029 26979 47087 26985
rect 47029 26945 47041 26979
rect 47075 26945 47087 26979
rect 47029 26939 47087 26945
rect 47121 26979 47179 26985
rect 47121 26945 47133 26979
rect 47167 26945 47179 26979
rect 47121 26939 47179 26945
rect 47397 26979 47455 26985
rect 47397 26945 47409 26979
rect 47443 26976 47455 26979
rect 48133 26979 48191 26985
rect 48133 26976 48145 26979
rect 47443 26948 48145 26976
rect 47443 26945 47455 26948
rect 47397 26939 47455 26945
rect 48133 26945 48145 26948
rect 48179 26945 48191 26979
rect 50522 26976 50528 26988
rect 50278 26962 50528 26976
rect 48133 26939 48191 26945
rect 50264 26948 50528 26962
rect 43640 26908 43668 26936
rect 43272 26880 43668 26908
rect 47136 26908 47164 26939
rect 48314 26908 48320 26920
rect 47136 26880 48320 26908
rect 48314 26868 48320 26880
rect 48372 26868 48378 26920
rect 48682 26868 48688 26920
rect 48740 26868 48746 26920
rect 48869 26911 48927 26917
rect 48869 26877 48881 26911
rect 48915 26877 48927 26911
rect 48869 26871 48927 26877
rect 47305 26843 47363 26849
rect 47305 26809 47317 26843
rect 47351 26840 47363 26843
rect 48222 26840 48228 26852
rect 47351 26812 48228 26840
rect 47351 26809 47363 26812
rect 47305 26803 47363 26809
rect 48222 26800 48228 26812
rect 48280 26800 48286 26852
rect 39761 26775 39819 26781
rect 39761 26772 39773 26775
rect 38626 26744 39773 26772
rect 39761 26741 39773 26744
rect 39807 26772 39819 26775
rect 40494 26772 40500 26784
rect 39807 26744 40500 26772
rect 39807 26741 39819 26744
rect 39761 26735 39819 26741
rect 40494 26732 40500 26744
rect 40552 26732 40558 26784
rect 42702 26732 42708 26784
rect 42760 26772 42766 26784
rect 43073 26775 43131 26781
rect 43073 26772 43085 26775
rect 42760 26744 43085 26772
rect 42760 26732 42766 26744
rect 43073 26741 43085 26744
rect 43119 26741 43131 26775
rect 43073 26735 43131 26741
rect 43622 26732 43628 26784
rect 43680 26732 43686 26784
rect 46842 26732 46848 26784
rect 46900 26732 46906 26784
rect 48884 26772 48912 26871
rect 49142 26868 49148 26920
rect 49200 26908 49206 26920
rect 50264 26908 50292 26948
rect 50522 26936 50528 26948
rect 50580 26936 50586 26988
rect 50798 26936 50804 26988
rect 50856 26976 50862 26988
rect 50893 26979 50951 26985
rect 50893 26976 50905 26979
rect 50856 26948 50905 26976
rect 50856 26936 50862 26948
rect 50893 26945 50905 26948
rect 50939 26945 50951 26979
rect 50893 26939 50951 26945
rect 51169 26979 51227 26985
rect 51169 26945 51181 26979
rect 51215 26976 51227 26979
rect 51994 26976 52000 26988
rect 51215 26948 52000 26976
rect 51215 26945 51227 26948
rect 51169 26939 51227 26945
rect 51994 26936 52000 26948
rect 52052 26936 52058 26988
rect 49200 26880 50292 26908
rect 49200 26868 49206 26880
rect 50614 26868 50620 26920
rect 50672 26868 50678 26920
rect 52733 26911 52791 26917
rect 52733 26877 52745 26911
rect 52779 26877 52791 26911
rect 52733 26871 52791 26877
rect 52178 26840 52184 26852
rect 50172 26812 52184 26840
rect 49694 26772 49700 26784
rect 48884 26744 49700 26772
rect 49694 26732 49700 26744
rect 49752 26772 49758 26784
rect 50172 26772 50200 26812
rect 52178 26800 52184 26812
rect 52236 26840 52242 26852
rect 52748 26840 52776 26871
rect 53006 26868 53012 26920
rect 53064 26868 53070 26920
rect 52236 26812 52776 26840
rect 52236 26800 52242 26812
rect 49752 26744 50200 26772
rect 49752 26732 49758 26744
rect 50982 26732 50988 26784
rect 51040 26772 51046 26784
rect 51077 26775 51135 26781
rect 51077 26772 51089 26775
rect 51040 26744 51089 26772
rect 51040 26732 51046 26744
rect 51077 26741 51089 26744
rect 51123 26741 51135 26775
rect 51077 26735 51135 26741
rect 54478 26732 54484 26784
rect 54536 26732 54542 26784
rect 1104 26682 58880 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 58880 26682
rect 1104 26608 58880 26630
rect 23474 26528 23480 26580
rect 23532 26568 23538 26580
rect 24397 26571 24455 26577
rect 24397 26568 24409 26571
rect 23532 26540 24409 26568
rect 23532 26528 23538 26540
rect 24397 26537 24409 26540
rect 24443 26537 24455 26571
rect 24397 26531 24455 26537
rect 25133 26571 25191 26577
rect 25133 26537 25145 26571
rect 25179 26568 25191 26571
rect 25222 26568 25228 26580
rect 25179 26540 25228 26568
rect 25179 26537 25191 26540
rect 25133 26531 25191 26537
rect 25222 26528 25228 26540
rect 25280 26528 25286 26580
rect 29086 26568 29092 26580
rect 28092 26540 29092 26568
rect 25777 26503 25835 26509
rect 25777 26500 25789 26503
rect 25424 26472 25789 26500
rect 25222 26432 25228 26444
rect 24780 26404 25228 26432
rect 24780 26376 24808 26404
rect 25222 26392 25228 26404
rect 25280 26392 25286 26444
rect 24581 26367 24639 26373
rect 24581 26333 24593 26367
rect 24627 26333 24639 26367
rect 24581 26327 24639 26333
rect 24596 26296 24624 26327
rect 24762 26324 24768 26376
rect 24820 26324 24826 26376
rect 24857 26367 24915 26373
rect 24857 26333 24869 26367
rect 24903 26364 24915 26367
rect 24946 26364 24952 26376
rect 24903 26336 24952 26364
rect 24903 26333 24915 26336
rect 24857 26327 24915 26333
rect 24946 26324 24952 26336
rect 25004 26324 25010 26376
rect 25314 26324 25320 26376
rect 25372 26324 25378 26376
rect 25424 26373 25452 26472
rect 25777 26469 25789 26472
rect 25823 26469 25835 26503
rect 25777 26463 25835 26469
rect 27525 26503 27583 26509
rect 27525 26469 27537 26503
rect 27571 26500 27583 26503
rect 27982 26500 27988 26512
rect 27571 26472 27988 26500
rect 27571 26469 27583 26472
rect 27525 26463 27583 26469
rect 27982 26460 27988 26472
rect 28040 26460 28046 26512
rect 25498 26392 25504 26444
rect 25556 26432 25562 26444
rect 25593 26435 25651 26441
rect 25593 26432 25605 26435
rect 25556 26404 25605 26432
rect 25556 26392 25562 26404
rect 25593 26401 25605 26404
rect 25639 26401 25651 26435
rect 26421 26435 26479 26441
rect 26421 26432 26433 26435
rect 25593 26395 25651 26401
rect 25700 26404 26433 26432
rect 25700 26373 25728 26404
rect 26421 26401 26433 26404
rect 26467 26401 26479 26435
rect 27798 26432 27804 26444
rect 26421 26395 26479 26401
rect 26896 26404 27804 26432
rect 25409 26367 25467 26373
rect 25409 26333 25421 26367
rect 25455 26333 25467 26367
rect 25409 26327 25467 26333
rect 25685 26367 25743 26373
rect 25685 26333 25697 26367
rect 25731 26333 25743 26367
rect 25685 26327 25743 26333
rect 25958 26324 25964 26376
rect 26016 26324 26022 26376
rect 26326 26324 26332 26376
rect 26384 26364 26390 26376
rect 26896 26364 26924 26404
rect 27798 26392 27804 26404
rect 27856 26392 27862 26444
rect 26384 26336 26924 26364
rect 26973 26367 27031 26373
rect 26384 26324 26390 26336
rect 26973 26333 26985 26367
rect 27019 26333 27031 26367
rect 26973 26327 27031 26333
rect 24964 26296 24992 26324
rect 26053 26299 26111 26305
rect 26053 26296 26065 26299
rect 24596 26268 24900 26296
rect 24964 26268 26065 26296
rect 24872 26240 24900 26268
rect 26053 26265 26065 26268
rect 26099 26265 26111 26299
rect 26053 26259 26111 26265
rect 26145 26299 26203 26305
rect 26145 26265 26157 26299
rect 26191 26265 26203 26299
rect 26145 26259 26203 26265
rect 22738 26188 22744 26240
rect 22796 26188 22802 26240
rect 24854 26188 24860 26240
rect 24912 26188 24918 26240
rect 25222 26188 25228 26240
rect 25280 26228 25286 26240
rect 26160 26228 26188 26259
rect 26234 26256 26240 26308
rect 26292 26296 26298 26308
rect 26786 26296 26792 26308
rect 26292 26268 26792 26296
rect 26292 26256 26298 26268
rect 26786 26256 26792 26268
rect 26844 26296 26850 26308
rect 26988 26296 27016 26327
rect 27706 26324 27712 26376
rect 27764 26324 27770 26376
rect 28092 26373 28120 26540
rect 29086 26528 29092 26540
rect 29144 26568 29150 26580
rect 30190 26568 30196 26580
rect 29144 26540 30196 26568
rect 29144 26528 29150 26540
rect 30190 26528 30196 26540
rect 30248 26528 30254 26580
rect 32309 26571 32367 26577
rect 32309 26537 32321 26571
rect 32355 26568 32367 26571
rect 32398 26568 32404 26580
rect 32355 26540 32404 26568
rect 32355 26537 32367 26540
rect 32309 26531 32367 26537
rect 32398 26528 32404 26540
rect 32456 26528 32462 26580
rect 34698 26528 34704 26580
rect 34756 26568 34762 26580
rect 34885 26571 34943 26577
rect 34885 26568 34897 26571
rect 34756 26540 34897 26568
rect 34756 26528 34762 26540
rect 34885 26537 34897 26540
rect 34931 26537 34943 26571
rect 34885 26531 34943 26537
rect 35158 26528 35164 26580
rect 35216 26568 35222 26580
rect 35802 26568 35808 26580
rect 35216 26540 35808 26568
rect 35216 26528 35222 26540
rect 35802 26528 35808 26540
rect 35860 26528 35866 26580
rect 36630 26568 36636 26580
rect 36234 26540 36636 26568
rect 28997 26503 29055 26509
rect 28997 26469 29009 26503
rect 29043 26500 29055 26503
rect 32858 26500 32864 26512
rect 29043 26472 32864 26500
rect 29043 26469 29055 26472
rect 28997 26463 29055 26469
rect 32858 26460 32864 26472
rect 32916 26460 32922 26512
rect 33686 26460 33692 26512
rect 33744 26500 33750 26512
rect 33744 26472 35572 26500
rect 33744 26460 33750 26472
rect 29914 26432 29920 26444
rect 28736 26404 29920 26432
rect 28736 26373 28764 26404
rect 29914 26392 29920 26404
rect 29972 26392 29978 26444
rect 30190 26392 30196 26444
rect 30248 26392 30254 26444
rect 33318 26432 33324 26444
rect 32600 26404 33324 26432
rect 28077 26367 28135 26373
rect 28077 26333 28089 26367
rect 28123 26333 28135 26367
rect 28077 26327 28135 26333
rect 28721 26367 28779 26373
rect 28721 26333 28733 26367
rect 28767 26333 28779 26367
rect 28721 26327 28779 26333
rect 28810 26324 28816 26376
rect 28868 26324 28874 26376
rect 29089 26367 29147 26373
rect 29089 26333 29101 26367
rect 29135 26364 29147 26367
rect 29641 26367 29699 26373
rect 29641 26364 29653 26367
rect 29135 26336 29653 26364
rect 29135 26333 29147 26336
rect 29089 26327 29147 26333
rect 29641 26333 29653 26336
rect 29687 26333 29699 26367
rect 29641 26327 29699 26333
rect 32490 26324 32496 26376
rect 32548 26324 32554 26376
rect 32600 26373 32628 26404
rect 33318 26392 33324 26404
rect 33376 26392 33382 26444
rect 34514 26392 34520 26444
rect 34572 26432 34578 26444
rect 34698 26432 34704 26444
rect 34572 26404 34704 26432
rect 34572 26392 34578 26404
rect 34698 26392 34704 26404
rect 34756 26392 34762 26444
rect 34790 26392 34796 26444
rect 34848 26432 34854 26444
rect 35345 26435 35403 26441
rect 34848 26404 35204 26432
rect 34848 26392 34854 26404
rect 32585 26367 32643 26373
rect 32585 26333 32597 26367
rect 32631 26333 32643 26367
rect 32585 26327 32643 26333
rect 32861 26367 32919 26373
rect 32861 26333 32873 26367
rect 32907 26364 32919 26367
rect 33042 26364 33048 26376
rect 32907 26336 33048 26364
rect 32907 26333 32919 26336
rect 32861 26327 32919 26333
rect 33042 26324 33048 26336
rect 33100 26324 33106 26376
rect 33134 26324 33140 26376
rect 33192 26364 33198 26376
rect 34422 26364 34428 26376
rect 33192 26336 34428 26364
rect 33192 26324 33198 26336
rect 34422 26324 34428 26336
rect 34480 26364 34486 26376
rect 35066 26364 35072 26376
rect 34480 26336 35072 26364
rect 34480 26324 34486 26336
rect 35066 26324 35072 26336
rect 35124 26324 35130 26376
rect 35176 26373 35204 26404
rect 35345 26401 35357 26435
rect 35391 26401 35403 26435
rect 35345 26395 35403 26401
rect 35544 26432 35572 26472
rect 35894 26460 35900 26512
rect 35952 26500 35958 26512
rect 36081 26503 36139 26509
rect 36081 26500 36093 26503
rect 35952 26472 36093 26500
rect 35952 26460 35958 26472
rect 36081 26469 36093 26472
rect 36127 26469 36139 26503
rect 36234 26500 36262 26540
rect 36630 26528 36636 26540
rect 36688 26528 36694 26580
rect 38930 26528 38936 26580
rect 38988 26528 38994 26580
rect 40218 26528 40224 26580
rect 40276 26528 40282 26580
rect 40494 26528 40500 26580
rect 40552 26568 40558 26580
rect 44174 26568 44180 26580
rect 40552 26540 44180 26568
rect 40552 26528 40558 26540
rect 44174 26528 44180 26540
rect 44232 26528 44238 26580
rect 48317 26571 48375 26577
rect 48317 26537 48329 26571
rect 48363 26568 48375 26571
rect 48682 26568 48688 26580
rect 48363 26540 48688 26568
rect 48363 26537 48375 26540
rect 48317 26531 48375 26537
rect 48682 26528 48688 26540
rect 48740 26528 48746 26580
rect 49329 26571 49387 26577
rect 49329 26537 49341 26571
rect 49375 26568 49387 26571
rect 49602 26568 49608 26580
rect 49375 26540 49608 26568
rect 49375 26537 49387 26540
rect 49329 26531 49387 26537
rect 49602 26528 49608 26540
rect 49660 26528 49666 26580
rect 49712 26540 49888 26568
rect 36722 26500 36728 26512
rect 36081 26463 36139 26469
rect 36188 26472 36262 26500
rect 36372 26472 36728 26500
rect 36188 26441 36216 26472
rect 36173 26435 36231 26441
rect 35544 26404 36032 26432
rect 35161 26367 35219 26373
rect 35161 26333 35173 26367
rect 35207 26333 35219 26367
rect 35161 26327 35219 26333
rect 27801 26299 27859 26305
rect 27801 26296 27813 26299
rect 26844 26268 27813 26296
rect 26844 26256 26850 26268
rect 27801 26265 27813 26268
rect 27847 26265 27859 26299
rect 27801 26259 27859 26265
rect 27893 26299 27951 26305
rect 27893 26265 27905 26299
rect 27939 26265 27951 26299
rect 27893 26259 27951 26265
rect 27706 26228 27712 26240
rect 25280 26200 27712 26228
rect 25280 26188 25286 26200
rect 27706 26188 27712 26200
rect 27764 26228 27770 26240
rect 27908 26228 27936 26259
rect 28350 26256 28356 26308
rect 28408 26296 28414 26308
rect 30558 26296 30564 26308
rect 28408 26268 30564 26296
rect 28408 26256 28414 26268
rect 30558 26256 30564 26268
rect 30616 26256 30622 26308
rect 32398 26256 32404 26308
rect 32456 26296 32462 26308
rect 32677 26299 32735 26305
rect 32677 26296 32689 26299
rect 32456 26268 32689 26296
rect 32456 26256 32462 26268
rect 32677 26265 32689 26268
rect 32723 26296 32735 26299
rect 35360 26296 35388 26395
rect 35544 26373 35572 26404
rect 35437 26367 35495 26373
rect 35437 26333 35449 26367
rect 35483 26364 35495 26367
rect 35529 26367 35587 26373
rect 35529 26364 35541 26367
rect 35483 26336 35541 26364
rect 35483 26333 35495 26336
rect 35437 26327 35495 26333
rect 35529 26333 35541 26336
rect 35575 26333 35587 26367
rect 35529 26327 35587 26333
rect 35618 26324 35624 26376
rect 35676 26364 35682 26376
rect 35713 26367 35771 26373
rect 35713 26364 35725 26367
rect 35676 26336 35725 26364
rect 35676 26324 35682 26336
rect 35713 26333 35725 26336
rect 35759 26333 35771 26367
rect 35713 26327 35771 26333
rect 35894 26324 35900 26376
rect 35952 26324 35958 26376
rect 36004 26364 36032 26404
rect 36173 26401 36185 26435
rect 36219 26401 36231 26435
rect 36372 26432 36400 26472
rect 36722 26460 36728 26472
rect 36780 26500 36786 26512
rect 39022 26500 39028 26512
rect 36780 26472 39028 26500
rect 36780 26460 36786 26472
rect 39022 26460 39028 26472
rect 39080 26460 39086 26512
rect 39117 26503 39175 26509
rect 39117 26469 39129 26503
rect 39163 26500 39175 26503
rect 40126 26500 40132 26512
rect 39163 26472 40132 26500
rect 39163 26469 39175 26472
rect 39117 26463 39175 26469
rect 40126 26460 40132 26472
rect 40184 26460 40190 26512
rect 36633 26435 36691 26441
rect 36633 26432 36645 26435
rect 36173 26395 36231 26401
rect 36280 26404 36400 26432
rect 36556 26404 36645 26432
rect 36280 26364 36308 26404
rect 36004 26336 36308 26364
rect 36354 26324 36360 26376
rect 36412 26324 36418 26376
rect 36446 26324 36452 26376
rect 36504 26324 36510 26376
rect 35805 26299 35863 26305
rect 32723 26268 35296 26296
rect 35360 26268 35664 26296
rect 32723 26265 32735 26268
rect 32677 26259 32735 26265
rect 35268 26240 35296 26268
rect 27764 26200 27936 26228
rect 27764 26188 27770 26200
rect 28534 26188 28540 26240
rect 28592 26188 28598 26240
rect 30926 26188 30932 26240
rect 30984 26228 30990 26240
rect 33226 26228 33232 26240
rect 30984 26200 33232 26228
rect 30984 26188 30990 26200
rect 33226 26188 33232 26200
rect 33284 26188 33290 26240
rect 35250 26188 35256 26240
rect 35308 26228 35314 26240
rect 35526 26228 35532 26240
rect 35308 26200 35532 26228
rect 35308 26188 35314 26200
rect 35526 26188 35532 26200
rect 35584 26188 35590 26240
rect 35636 26228 35664 26268
rect 35805 26265 35817 26299
rect 35851 26296 35863 26299
rect 36262 26296 36268 26308
rect 35851 26268 36268 26296
rect 35851 26265 35863 26268
rect 35805 26259 35863 26265
rect 36262 26256 36268 26268
rect 36320 26256 36326 26308
rect 36170 26228 36176 26240
rect 35636 26200 36176 26228
rect 36170 26188 36176 26200
rect 36228 26228 36234 26240
rect 36556 26228 36584 26404
rect 36633 26401 36645 26404
rect 36679 26401 36691 26435
rect 36633 26395 36691 26401
rect 38654 26392 38660 26444
rect 38712 26432 38718 26444
rect 39669 26435 39727 26441
rect 39669 26432 39681 26435
rect 38712 26404 39681 26432
rect 38712 26392 38718 26404
rect 39669 26401 39681 26404
rect 39715 26401 39727 26435
rect 40236 26432 40264 26528
rect 42886 26460 42892 26512
rect 42944 26500 42950 26512
rect 43438 26500 43444 26512
rect 42944 26472 43444 26500
rect 42944 26460 42950 26472
rect 43438 26460 43444 26472
rect 43496 26460 43502 26512
rect 45830 26460 45836 26512
rect 45888 26500 45894 26512
rect 45925 26503 45983 26509
rect 45925 26500 45937 26503
rect 45888 26472 45937 26500
rect 45888 26460 45894 26472
rect 45925 26469 45937 26472
rect 45971 26500 45983 26503
rect 46385 26503 46443 26509
rect 46385 26500 46397 26503
rect 45971 26472 46397 26500
rect 45971 26469 45983 26472
rect 45925 26463 45983 26469
rect 46385 26469 46397 26472
rect 46431 26469 46443 26503
rect 49510 26500 49516 26512
rect 46385 26463 46443 26469
rect 48286 26472 49516 26500
rect 40589 26435 40647 26441
rect 40589 26432 40601 26435
rect 40236 26404 40601 26432
rect 39669 26395 39727 26401
rect 40589 26401 40601 26404
rect 40635 26401 40647 26435
rect 41233 26435 41291 26441
rect 41233 26432 41245 26435
rect 40589 26395 40647 26401
rect 40788 26404 41245 26432
rect 36725 26367 36783 26373
rect 36725 26333 36737 26367
rect 36771 26364 36783 26367
rect 37182 26364 37188 26376
rect 36771 26336 37188 26364
rect 36771 26333 36783 26336
rect 36725 26327 36783 26333
rect 37182 26324 37188 26336
rect 37240 26324 37246 26376
rect 38841 26367 38899 26373
rect 38841 26333 38853 26367
rect 38887 26333 38899 26367
rect 38841 26327 38899 26333
rect 39025 26367 39083 26373
rect 39025 26333 39037 26367
rect 39071 26364 39083 26367
rect 39485 26367 39543 26373
rect 39071 26336 39436 26364
rect 39071 26333 39083 26336
rect 39025 26327 39083 26333
rect 36228 26200 36584 26228
rect 38856 26228 38884 26327
rect 39298 26228 39304 26240
rect 38856 26200 39304 26228
rect 36228 26188 36234 26200
rect 39298 26188 39304 26200
rect 39356 26188 39362 26240
rect 39408 26237 39436 26336
rect 39485 26333 39497 26367
rect 39531 26364 39543 26367
rect 39942 26364 39948 26376
rect 39531 26336 39948 26364
rect 39531 26333 39543 26336
rect 39485 26327 39543 26333
rect 39942 26324 39948 26336
rect 40000 26324 40006 26376
rect 40175 26333 40233 26339
rect 40175 26299 40187 26333
rect 40221 26330 40233 26333
rect 40221 26299 40234 26330
rect 40494 26324 40500 26376
rect 40552 26364 40558 26376
rect 40681 26367 40739 26373
rect 40681 26364 40693 26367
rect 40552 26336 40693 26364
rect 40552 26324 40558 26336
rect 40681 26333 40693 26336
rect 40727 26333 40739 26367
rect 40681 26327 40739 26333
rect 40175 26296 40234 26299
rect 40405 26299 40463 26305
rect 40175 26293 40248 26296
rect 40206 26268 40248 26293
rect 40220 26240 40248 26268
rect 40405 26265 40417 26299
rect 40451 26296 40463 26299
rect 40512 26296 40540 26324
rect 40451 26268 40540 26296
rect 40451 26265 40463 26268
rect 40405 26259 40463 26265
rect 39393 26231 39451 26237
rect 39393 26197 39405 26231
rect 39439 26228 39451 26231
rect 39482 26228 39488 26240
rect 39439 26200 39488 26228
rect 39439 26197 39451 26200
rect 39393 26191 39451 26197
rect 39482 26188 39488 26200
rect 39540 26188 39546 26240
rect 40034 26188 40040 26240
rect 40092 26188 40098 26240
rect 40218 26188 40224 26240
rect 40276 26228 40282 26240
rect 40788 26228 40816 26404
rect 41233 26401 41245 26404
rect 41279 26432 41291 26435
rect 42058 26432 42064 26444
rect 41279 26404 42064 26432
rect 41279 26401 41291 26404
rect 41233 26395 41291 26401
rect 42058 26392 42064 26404
rect 42116 26432 42122 26444
rect 42426 26432 42432 26444
rect 42116 26404 42432 26432
rect 42116 26392 42122 26404
rect 42426 26392 42432 26404
rect 42484 26392 42490 26444
rect 45554 26392 45560 26444
rect 45612 26432 45618 26444
rect 46290 26432 46296 26444
rect 45612 26404 46296 26432
rect 45612 26392 45618 26404
rect 46290 26392 46296 26404
rect 46348 26432 46354 26444
rect 46569 26435 46627 26441
rect 46569 26432 46581 26435
rect 46348 26404 46581 26432
rect 46348 26392 46354 26404
rect 46569 26401 46581 26404
rect 46615 26401 46627 26435
rect 46569 26395 46627 26401
rect 46842 26392 46848 26444
rect 46900 26392 46906 26444
rect 48038 26392 48044 26444
rect 48096 26432 48102 26444
rect 48286 26432 48314 26472
rect 49510 26460 49516 26472
rect 49568 26460 49574 26512
rect 48096 26404 48314 26432
rect 48096 26392 48102 26404
rect 40957 26367 41015 26373
rect 40957 26333 40969 26367
rect 41003 26364 41015 26367
rect 42886 26364 42892 26376
rect 41003 26336 42892 26364
rect 41003 26333 41015 26336
rect 40957 26327 41015 26333
rect 42886 26324 42892 26336
rect 42944 26324 42950 26376
rect 46201 26367 46259 26373
rect 46201 26333 46213 26367
rect 46247 26333 46259 26367
rect 46201 26327 46259 26333
rect 46477 26367 46535 26373
rect 46477 26333 46489 26367
rect 46523 26333 46535 26367
rect 46477 26327 46535 26333
rect 43346 26256 43352 26308
rect 43404 26296 43410 26308
rect 44910 26296 44916 26308
rect 43404 26268 44916 26296
rect 43404 26256 43410 26268
rect 44910 26256 44916 26268
rect 44968 26256 44974 26308
rect 46216 26296 46244 26327
rect 46492 26296 46520 26327
rect 48682 26324 48688 26376
rect 48740 26364 48746 26376
rect 49510 26373 49516 26376
rect 48740 26336 49280 26364
rect 48740 26324 48746 26336
rect 47118 26296 47124 26308
rect 46216 26268 46428 26296
rect 46492 26268 47124 26296
rect 40276 26200 40816 26228
rect 40276 26188 40282 26200
rect 42150 26188 42156 26240
rect 42208 26228 42214 26240
rect 43622 26228 43628 26240
rect 42208 26200 43628 26228
rect 42208 26188 42214 26200
rect 43622 26188 43628 26200
rect 43680 26188 43686 26240
rect 45922 26188 45928 26240
rect 45980 26228 45986 26240
rect 46017 26231 46075 26237
rect 46017 26228 46029 26231
rect 45980 26200 46029 26228
rect 45980 26188 45986 26200
rect 46017 26197 46029 26200
rect 46063 26197 46075 26231
rect 46400 26228 46428 26268
rect 47118 26256 47124 26268
rect 47176 26256 47182 26308
rect 48130 26296 48136 26308
rect 48070 26268 48136 26296
rect 48130 26256 48136 26268
rect 48188 26296 48194 26308
rect 48774 26296 48780 26308
rect 48188 26268 48780 26296
rect 48188 26256 48194 26268
rect 48774 26256 48780 26268
rect 48832 26296 48838 26308
rect 49142 26296 49148 26308
rect 48832 26268 49148 26296
rect 48832 26256 48838 26268
rect 49142 26256 49148 26268
rect 49200 26256 49206 26308
rect 49252 26296 49280 26336
rect 49508 26327 49516 26373
rect 49568 26364 49574 26376
rect 49712 26364 49740 26540
rect 49860 26500 49888 26540
rect 50798 26528 50804 26580
rect 50856 26528 50862 26580
rect 52457 26571 52515 26577
rect 52457 26537 52469 26571
rect 52503 26568 52515 26571
rect 53006 26568 53012 26580
rect 52503 26540 53012 26568
rect 52503 26537 52515 26540
rect 52457 26531 52515 26537
rect 53006 26528 53012 26540
rect 53064 26528 53070 26580
rect 50614 26500 50620 26512
rect 49860 26472 50620 26500
rect 50614 26460 50620 26472
rect 50672 26500 50678 26512
rect 51902 26500 51908 26512
rect 50672 26472 51908 26500
rect 50672 26460 50678 26472
rect 51902 26460 51908 26472
rect 51960 26460 51966 26512
rect 57882 26460 57888 26512
rect 57940 26500 57946 26512
rect 58437 26503 58495 26509
rect 58437 26500 58449 26503
rect 57940 26472 58449 26500
rect 57940 26460 57946 26472
rect 58437 26469 58449 26472
rect 58483 26469 58495 26503
rect 58437 26463 58495 26469
rect 50430 26392 50436 26444
rect 50488 26432 50494 26444
rect 50488 26404 50665 26432
rect 50488 26392 50494 26404
rect 49880 26367 49938 26373
rect 49880 26364 49892 26367
rect 49568 26336 49608 26364
rect 49712 26336 49892 26364
rect 49510 26324 49516 26327
rect 49568 26324 49574 26336
rect 49880 26333 49892 26336
rect 49926 26333 49938 26367
rect 49880 26327 49938 26333
rect 49970 26324 49976 26376
rect 50028 26364 50034 26376
rect 50157 26367 50215 26373
rect 50157 26364 50169 26367
rect 50028 26336 50169 26364
rect 50028 26324 50034 26336
rect 50157 26333 50169 26336
rect 50203 26333 50215 26367
rect 50157 26327 50215 26333
rect 50250 26367 50308 26373
rect 50250 26333 50262 26367
rect 50296 26333 50308 26367
rect 50250 26327 50308 26333
rect 49326 26296 49332 26308
rect 49252 26268 49332 26296
rect 49326 26256 49332 26268
rect 49384 26296 49390 26308
rect 49605 26299 49663 26305
rect 49605 26296 49617 26299
rect 49384 26268 49617 26296
rect 49384 26256 49390 26268
rect 49605 26265 49617 26268
rect 49651 26265 49663 26299
rect 49605 26259 49663 26265
rect 49694 26256 49700 26308
rect 49752 26256 49758 26308
rect 49786 26256 49792 26308
rect 49844 26296 49850 26308
rect 50265 26296 50293 26327
rect 50522 26324 50528 26376
rect 50580 26324 50586 26376
rect 50637 26373 50665 26404
rect 50982 26392 50988 26444
rect 51040 26432 51046 26444
rect 52825 26435 52883 26441
rect 52825 26432 52837 26435
rect 51040 26404 52837 26432
rect 51040 26392 51046 26404
rect 52825 26401 52837 26404
rect 52871 26401 52883 26435
rect 52825 26395 52883 26401
rect 50622 26367 50680 26373
rect 50622 26333 50634 26367
rect 50668 26333 50680 26367
rect 50622 26327 50680 26333
rect 52638 26324 52644 26376
rect 52696 26324 52702 26376
rect 52917 26367 52975 26373
rect 52917 26333 52929 26367
rect 52963 26364 52975 26367
rect 53561 26367 53619 26373
rect 53561 26364 53573 26367
rect 52963 26336 53573 26364
rect 52963 26333 52975 26336
rect 52917 26327 52975 26333
rect 53561 26333 53573 26336
rect 53607 26333 53619 26367
rect 53561 26327 53619 26333
rect 54113 26367 54171 26373
rect 54113 26333 54125 26367
rect 54159 26364 54171 26367
rect 54478 26364 54484 26376
rect 54159 26336 54484 26364
rect 54159 26333 54171 26336
rect 54113 26327 54171 26333
rect 49844 26268 50293 26296
rect 49844 26256 49850 26268
rect 48222 26228 48228 26240
rect 46400 26200 48228 26228
rect 46017 26191 46075 26197
rect 48222 26188 48228 26200
rect 48280 26188 48286 26240
rect 49050 26188 49056 26240
rect 49108 26228 49114 26240
rect 49970 26228 49976 26240
rect 49108 26200 49976 26228
rect 49108 26188 49114 26200
rect 49970 26188 49976 26200
rect 50028 26188 50034 26240
rect 50265 26228 50293 26268
rect 50430 26256 50436 26308
rect 50488 26256 50494 26308
rect 54128 26296 54156 26327
rect 54478 26324 54484 26336
rect 54536 26324 54542 26376
rect 58250 26324 58256 26376
rect 58308 26324 58314 26376
rect 53024 26268 54156 26296
rect 53024 26240 53052 26268
rect 53006 26228 53012 26240
rect 50265 26200 53012 26228
rect 53006 26188 53012 26200
rect 53064 26188 53070 26240
rect 1104 26138 58880 26160
rect 1104 26086 4874 26138
rect 4926 26086 4938 26138
rect 4990 26086 5002 26138
rect 5054 26086 5066 26138
rect 5118 26086 5130 26138
rect 5182 26086 35594 26138
rect 35646 26086 35658 26138
rect 35710 26086 35722 26138
rect 35774 26086 35786 26138
rect 35838 26086 35850 26138
rect 35902 26086 58880 26138
rect 1104 26064 58880 26086
rect 22278 25984 22284 26036
rect 22336 25984 22342 26036
rect 22738 25984 22744 26036
rect 22796 26024 22802 26036
rect 24673 26027 24731 26033
rect 24673 26024 24685 26027
rect 22796 25996 24685 26024
rect 22796 25984 22802 25996
rect 24673 25993 24685 25996
rect 24719 26024 24731 26027
rect 30101 26027 30159 26033
rect 24719 25996 25636 26024
rect 24719 25993 24731 25996
rect 24673 25987 24731 25993
rect 20162 25956 20168 25968
rect 19076 25928 20168 25956
rect 19076 25897 19104 25928
rect 20162 25916 20168 25928
rect 20220 25916 20226 25968
rect 22296 25956 22324 25984
rect 25133 25959 25191 25965
rect 22112 25928 22324 25956
rect 22480 25928 23428 25956
rect 19061 25891 19119 25897
rect 19061 25857 19073 25891
rect 19107 25857 19119 25891
rect 19061 25851 19119 25857
rect 19153 25891 19211 25897
rect 19153 25857 19165 25891
rect 19199 25857 19211 25891
rect 19153 25851 19211 25857
rect 19429 25891 19487 25897
rect 19429 25857 19441 25891
rect 19475 25888 19487 25891
rect 19610 25888 19616 25900
rect 19475 25860 19616 25888
rect 19475 25857 19487 25860
rect 19429 25851 19487 25857
rect 19168 25820 19196 25851
rect 19610 25848 19616 25860
rect 19668 25848 19674 25900
rect 22112 25897 22140 25928
rect 22092 25891 22150 25897
rect 22092 25857 22104 25891
rect 22138 25857 22150 25891
rect 22092 25851 22150 25857
rect 22189 25891 22247 25897
rect 22189 25857 22201 25891
rect 22235 25857 22247 25891
rect 22189 25851 22247 25857
rect 22281 25891 22339 25897
rect 22281 25857 22293 25891
rect 22327 25888 22339 25891
rect 22370 25888 22376 25900
rect 22327 25860 22376 25888
rect 22327 25857 22339 25860
rect 22281 25851 22339 25857
rect 19794 25820 19800 25832
rect 19168 25792 19800 25820
rect 19794 25780 19800 25792
rect 19852 25780 19858 25832
rect 20530 25780 20536 25832
rect 20588 25820 20594 25832
rect 22204 25820 22232 25851
rect 22370 25848 22376 25860
rect 22428 25848 22434 25900
rect 22480 25897 22508 25928
rect 22464 25891 22522 25897
rect 22464 25857 22476 25891
rect 22510 25857 22522 25891
rect 22464 25851 22522 25857
rect 22557 25891 22615 25897
rect 22557 25857 22569 25891
rect 22603 25888 22615 25891
rect 22738 25888 22744 25900
rect 22603 25860 22744 25888
rect 22603 25857 22615 25860
rect 22557 25851 22615 25857
rect 22738 25848 22744 25860
rect 22796 25848 22802 25900
rect 22833 25891 22891 25897
rect 22833 25857 22845 25891
rect 22879 25888 22891 25891
rect 23290 25888 23296 25900
rect 22879 25860 23296 25888
rect 22879 25857 22891 25860
rect 22833 25851 22891 25857
rect 23290 25848 23296 25860
rect 23348 25848 23354 25900
rect 23400 25832 23428 25928
rect 25133 25925 25145 25959
rect 25179 25925 25191 25959
rect 25133 25919 25191 25925
rect 23474 25848 23480 25900
rect 23532 25888 23538 25900
rect 24118 25888 24124 25900
rect 23532 25860 24124 25888
rect 23532 25848 23538 25860
rect 24118 25848 24124 25860
rect 24176 25888 24182 25900
rect 25038 25897 25044 25900
rect 24995 25891 25044 25897
rect 24995 25888 25007 25891
rect 24176 25860 25007 25888
rect 24176 25848 24182 25860
rect 24995 25857 25007 25860
rect 25041 25857 25044 25891
rect 24995 25851 25044 25857
rect 25038 25848 25044 25851
rect 25096 25848 25102 25900
rect 23014 25820 23020 25832
rect 20588 25792 23020 25820
rect 20588 25780 20594 25792
rect 23014 25780 23020 25792
rect 23072 25780 23078 25832
rect 23109 25823 23167 25829
rect 23109 25789 23121 25823
rect 23155 25820 23167 25823
rect 23201 25823 23259 25829
rect 23201 25820 23213 25823
rect 23155 25792 23213 25820
rect 23155 25789 23167 25792
rect 23109 25783 23167 25789
rect 23201 25789 23213 25792
rect 23247 25789 23259 25823
rect 23201 25783 23259 25789
rect 23382 25780 23388 25832
rect 23440 25820 23446 25832
rect 23753 25823 23811 25829
rect 23753 25820 23765 25823
rect 23440 25792 23765 25820
rect 23440 25780 23446 25792
rect 23753 25789 23765 25792
rect 23799 25820 23811 25823
rect 25148 25820 25176 25919
rect 25222 25848 25228 25900
rect 25280 25848 25286 25900
rect 25408 25891 25466 25897
rect 25408 25857 25420 25891
rect 25454 25857 25466 25891
rect 25408 25851 25466 25857
rect 25501 25891 25559 25897
rect 25501 25857 25513 25891
rect 25547 25888 25559 25891
rect 25608 25888 25636 25996
rect 27724 25996 29960 26024
rect 26510 25916 26516 25968
rect 26568 25956 26574 25968
rect 27724 25956 27752 25996
rect 26568 25928 27752 25956
rect 26568 25916 26574 25928
rect 27798 25916 27804 25968
rect 27856 25956 27862 25968
rect 27856 25928 28304 25956
rect 27856 25916 27862 25928
rect 25547 25860 25636 25888
rect 25547 25857 25559 25860
rect 25501 25851 25559 25857
rect 25424 25820 25452 25851
rect 27614 25848 27620 25900
rect 27672 25888 27678 25900
rect 27709 25891 27767 25897
rect 27709 25888 27721 25891
rect 27672 25860 27721 25888
rect 27672 25848 27678 25860
rect 27709 25857 27721 25860
rect 27755 25857 27767 25891
rect 27709 25851 27767 25857
rect 27893 25891 27951 25897
rect 27893 25857 27905 25891
rect 27939 25857 27951 25891
rect 27893 25851 27951 25857
rect 26234 25820 26240 25832
rect 23799 25792 25268 25820
rect 25424 25792 26240 25820
rect 23799 25789 23811 25792
rect 23753 25783 23811 25789
rect 19337 25755 19395 25761
rect 19337 25721 19349 25755
rect 19383 25752 19395 25755
rect 24762 25752 24768 25764
rect 19383 25724 24768 25752
rect 19383 25721 19395 25724
rect 19337 25715 19395 25721
rect 18230 25644 18236 25696
rect 18288 25684 18294 25696
rect 18877 25687 18935 25693
rect 18877 25684 18889 25687
rect 18288 25656 18889 25684
rect 18288 25644 18294 25656
rect 18877 25653 18889 25656
rect 18923 25653 18935 25687
rect 18877 25647 18935 25653
rect 21174 25644 21180 25696
rect 21232 25684 21238 25696
rect 21913 25687 21971 25693
rect 21913 25684 21925 25687
rect 21232 25656 21925 25684
rect 21232 25644 21238 25656
rect 21913 25653 21925 25656
rect 21959 25653 21971 25687
rect 21913 25647 21971 25653
rect 22002 25644 22008 25696
rect 22060 25684 22066 25696
rect 23032 25693 23060 25724
rect 24762 25712 24768 25724
rect 24820 25712 24826 25764
rect 24854 25712 24860 25764
rect 24912 25712 24918 25764
rect 22649 25687 22707 25693
rect 22649 25684 22661 25687
rect 22060 25656 22661 25684
rect 22060 25644 22066 25656
rect 22649 25653 22661 25656
rect 22695 25653 22707 25687
rect 22649 25647 22707 25653
rect 23017 25687 23075 25693
rect 23017 25653 23029 25687
rect 23063 25653 23075 25687
rect 25240 25684 25268 25792
rect 26234 25780 26240 25792
rect 26292 25780 26298 25832
rect 26970 25780 26976 25832
rect 27028 25820 27034 25832
rect 27908 25820 27936 25851
rect 27982 25848 27988 25900
rect 28040 25848 28046 25900
rect 28276 25897 28304 25928
rect 28534 25916 28540 25968
rect 28592 25956 28598 25968
rect 28629 25959 28687 25965
rect 28629 25956 28641 25959
rect 28592 25928 28641 25956
rect 28592 25916 28598 25928
rect 28629 25925 28641 25928
rect 28675 25925 28687 25959
rect 28629 25919 28687 25925
rect 28902 25916 28908 25968
rect 28960 25956 28966 25968
rect 29932 25956 29960 25996
rect 30101 25993 30113 26027
rect 30147 26024 30159 26027
rect 30190 26024 30196 26036
rect 30147 25996 30196 26024
rect 30147 25993 30159 25996
rect 30101 25987 30159 25993
rect 30190 25984 30196 25996
rect 30248 25984 30254 26036
rect 31726 25996 35480 26024
rect 31726 25956 31754 25996
rect 28960 25928 29118 25956
rect 29932 25928 31754 25956
rect 32401 25959 32459 25965
rect 28960 25916 28966 25928
rect 32401 25925 32413 25959
rect 32447 25956 32459 25959
rect 32950 25956 32956 25968
rect 32447 25928 32956 25956
rect 32447 25925 32459 25928
rect 32401 25919 32459 25925
rect 32950 25916 32956 25928
rect 33008 25916 33014 25968
rect 35452 25956 35480 25996
rect 35526 25984 35532 26036
rect 35584 26024 35590 26036
rect 35584 25996 35940 26024
rect 35584 25984 35590 25996
rect 35618 25956 35624 25968
rect 35452 25928 35624 25956
rect 35618 25916 35624 25928
rect 35676 25916 35682 25968
rect 35912 25965 35940 25996
rect 37642 25984 37648 26036
rect 37700 26024 37706 26036
rect 39235 26027 39293 26033
rect 37700 25996 39160 26024
rect 37700 25984 37706 25996
rect 35897 25959 35955 25965
rect 35897 25925 35909 25959
rect 35943 25956 35955 25959
rect 36906 25956 36912 25968
rect 35943 25928 36912 25956
rect 35943 25925 35955 25928
rect 35897 25919 35955 25925
rect 36906 25916 36912 25928
rect 36964 25916 36970 25968
rect 38930 25916 38936 25968
rect 38988 25956 38994 25968
rect 39025 25959 39083 25965
rect 39025 25956 39037 25959
rect 38988 25928 39037 25956
rect 38988 25916 38994 25928
rect 39025 25925 39037 25928
rect 39071 25925 39083 25959
rect 39132 25956 39160 25996
rect 39235 25993 39247 26027
rect 39281 26024 39293 26027
rect 40034 26024 40040 26036
rect 39281 25996 40040 26024
rect 39281 25993 39293 25996
rect 39235 25987 39293 25993
rect 40034 25984 40040 25996
rect 40092 25984 40098 26036
rect 42518 25984 42524 26036
rect 42576 26024 42582 26036
rect 42613 26027 42671 26033
rect 42613 26024 42625 26027
rect 42576 25996 42625 26024
rect 42576 25984 42582 25996
rect 42613 25993 42625 25996
rect 42659 26024 42671 26027
rect 42659 25996 42840 26024
rect 42659 25993 42671 25996
rect 42613 25987 42671 25993
rect 40862 25956 40868 25968
rect 39132 25928 40868 25956
rect 39025 25919 39083 25925
rect 40862 25916 40868 25928
rect 40920 25916 40926 25968
rect 42702 25916 42708 25968
rect 42760 25916 42766 25968
rect 42812 25956 42840 25996
rect 42886 25984 42892 26036
rect 42944 26033 42950 26036
rect 42944 26027 42963 26033
rect 42951 25993 42963 26027
rect 42944 25987 42963 25993
rect 44545 26027 44603 26033
rect 44545 25993 44557 26027
rect 44591 26024 44603 26027
rect 45738 26024 45744 26036
rect 44591 25996 45744 26024
rect 44591 25993 44603 25996
rect 44545 25987 44603 25993
rect 42944 25984 42950 25987
rect 43806 25956 43812 25968
rect 42812 25928 43812 25956
rect 43806 25916 43812 25928
rect 43864 25916 43870 25968
rect 28261 25891 28319 25897
rect 28261 25857 28273 25891
rect 28307 25857 28319 25891
rect 28261 25851 28319 25857
rect 27028 25792 27936 25820
rect 28276 25820 28304 25851
rect 28350 25848 28356 25900
rect 28408 25848 28414 25900
rect 32122 25848 32128 25900
rect 32180 25848 32186 25900
rect 32309 25891 32367 25897
rect 32309 25857 32321 25891
rect 32355 25888 32367 25891
rect 32493 25891 32551 25897
rect 32355 25860 32444 25888
rect 32355 25857 32367 25860
rect 32309 25851 32367 25857
rect 32416 25832 32444 25860
rect 32493 25857 32505 25891
rect 32539 25888 32551 25891
rect 32582 25888 32588 25900
rect 32539 25860 32588 25888
rect 32539 25857 32551 25860
rect 32493 25851 32551 25857
rect 32582 25848 32588 25860
rect 32640 25888 32646 25900
rect 35158 25888 35164 25900
rect 32640 25860 35164 25888
rect 32640 25848 32646 25860
rect 35158 25848 35164 25860
rect 35216 25888 35222 25900
rect 35713 25891 35771 25897
rect 35713 25888 35725 25891
rect 35216 25860 35725 25888
rect 35216 25848 35222 25860
rect 35713 25857 35725 25860
rect 35759 25857 35771 25891
rect 35713 25851 35771 25857
rect 28626 25820 28632 25832
rect 28276 25792 28632 25820
rect 27028 25780 27034 25792
rect 28626 25780 28632 25792
rect 28684 25780 28690 25832
rect 32398 25780 32404 25832
rect 32456 25780 32462 25832
rect 35250 25780 35256 25832
rect 35308 25820 35314 25832
rect 35526 25820 35532 25832
rect 35308 25792 35532 25820
rect 35308 25780 35314 25792
rect 35526 25780 35532 25792
rect 35584 25780 35590 25832
rect 35728 25820 35756 25851
rect 35802 25848 35808 25900
rect 35860 25848 35866 25900
rect 36078 25848 36084 25900
rect 36136 25888 36142 25900
rect 37182 25888 37188 25900
rect 36136 25860 37188 25888
rect 36136 25848 36142 25860
rect 37182 25848 37188 25860
rect 37240 25848 37246 25900
rect 39298 25848 39304 25900
rect 39356 25888 39362 25900
rect 39666 25888 39672 25900
rect 39356 25860 39672 25888
rect 39356 25848 39362 25860
rect 39666 25848 39672 25860
rect 39724 25848 39730 25900
rect 42334 25888 42340 25900
rect 39776 25860 42340 25888
rect 36722 25820 36728 25832
rect 35728 25792 36728 25820
rect 36722 25780 36728 25792
rect 36780 25780 36786 25832
rect 39390 25820 39396 25832
rect 38626 25792 39396 25820
rect 25314 25712 25320 25764
rect 25372 25752 25378 25764
rect 25869 25755 25927 25761
rect 25869 25752 25881 25755
rect 25372 25724 25881 25752
rect 25372 25712 25378 25724
rect 25869 25721 25881 25724
rect 25915 25752 25927 25755
rect 38626 25752 38654 25792
rect 39390 25780 39396 25792
rect 39448 25780 39454 25832
rect 39482 25780 39488 25832
rect 39540 25780 39546 25832
rect 39776 25752 39804 25860
rect 42334 25848 42340 25860
rect 42392 25848 42398 25900
rect 43901 25891 43959 25897
rect 43901 25888 43913 25891
rect 43364 25860 43913 25888
rect 39942 25780 39948 25832
rect 40000 25780 40006 25832
rect 40037 25823 40095 25829
rect 40037 25789 40049 25823
rect 40083 25820 40095 25823
rect 40310 25820 40316 25832
rect 40083 25792 40316 25820
rect 40083 25789 40095 25792
rect 40037 25783 40095 25789
rect 40310 25780 40316 25792
rect 40368 25780 40374 25832
rect 41966 25780 41972 25832
rect 42024 25820 42030 25832
rect 43364 25829 43392 25860
rect 43901 25857 43913 25860
rect 43947 25857 43959 25891
rect 43901 25851 43959 25857
rect 43993 25891 44051 25897
rect 43993 25857 44005 25891
rect 44039 25857 44051 25891
rect 43993 25851 44051 25857
rect 43165 25823 43223 25829
rect 43165 25820 43177 25823
rect 42024 25792 43177 25820
rect 42024 25780 42030 25792
rect 43165 25789 43177 25792
rect 43211 25789 43223 25823
rect 43165 25783 43223 25789
rect 43349 25823 43407 25829
rect 43349 25789 43361 25823
rect 43395 25789 43407 25823
rect 43349 25783 43407 25789
rect 25915 25724 28304 25752
rect 25915 25721 25927 25724
rect 25869 25715 25927 25721
rect 25406 25684 25412 25696
rect 25240 25656 25412 25684
rect 23017 25647 23075 25653
rect 25406 25644 25412 25656
rect 25464 25644 25470 25696
rect 25498 25644 25504 25696
rect 25556 25684 25562 25696
rect 26142 25684 26148 25696
rect 25556 25656 26148 25684
rect 25556 25644 25562 25656
rect 26142 25644 26148 25656
rect 26200 25684 26206 25696
rect 28169 25687 28227 25693
rect 28169 25684 28181 25687
rect 26200 25656 28181 25684
rect 26200 25644 26206 25656
rect 28169 25653 28181 25656
rect 28215 25653 28227 25687
rect 28276 25684 28304 25724
rect 32600 25724 38654 25752
rect 39224 25724 39804 25752
rect 28718 25684 28724 25696
rect 28276 25656 28724 25684
rect 28169 25647 28227 25653
rect 28718 25644 28724 25656
rect 28776 25644 28782 25696
rect 31754 25644 31760 25696
rect 31812 25684 31818 25696
rect 32600 25684 32628 25724
rect 31812 25656 32628 25684
rect 32677 25687 32735 25693
rect 31812 25644 31818 25656
rect 32677 25653 32689 25687
rect 32723 25684 32735 25687
rect 33318 25684 33324 25696
rect 32723 25656 33324 25684
rect 32723 25653 32735 25656
rect 32677 25647 32735 25653
rect 33318 25644 33324 25656
rect 33376 25644 33382 25696
rect 35526 25644 35532 25696
rect 35584 25644 35590 25696
rect 35618 25644 35624 25696
rect 35676 25684 35682 25696
rect 37734 25684 37740 25696
rect 35676 25656 37740 25684
rect 35676 25644 35682 25656
rect 37734 25644 37740 25656
rect 37792 25644 37798 25696
rect 38746 25644 38752 25696
rect 38804 25684 38810 25696
rect 39224 25693 39252 25724
rect 39850 25712 39856 25764
rect 39908 25752 39914 25764
rect 43073 25755 43131 25761
rect 39908 25724 43024 25752
rect 39908 25712 39914 25724
rect 39209 25687 39267 25693
rect 39209 25684 39221 25687
rect 38804 25656 39221 25684
rect 38804 25644 38810 25656
rect 39209 25653 39221 25656
rect 39255 25653 39267 25687
rect 39209 25647 39267 25653
rect 39390 25644 39396 25696
rect 39448 25684 39454 25696
rect 40221 25687 40279 25693
rect 40221 25684 40233 25687
rect 39448 25656 40233 25684
rect 39448 25644 39454 25656
rect 40221 25653 40233 25656
rect 40267 25684 40279 25687
rect 40586 25684 40592 25696
rect 40267 25656 40592 25684
rect 40267 25653 40279 25656
rect 40221 25647 40279 25653
rect 40586 25644 40592 25656
rect 40644 25644 40650 25696
rect 42610 25644 42616 25696
rect 42668 25684 42674 25696
rect 42889 25687 42947 25693
rect 42889 25684 42901 25687
rect 42668 25656 42901 25684
rect 42668 25644 42674 25656
rect 42889 25653 42901 25656
rect 42935 25653 42947 25687
rect 42996 25684 43024 25724
rect 43073 25721 43085 25755
rect 43119 25752 43131 25755
rect 43364 25752 43392 25783
rect 43438 25780 43444 25832
rect 43496 25820 43502 25832
rect 44008 25820 44036 25851
rect 44174 25848 44180 25900
rect 44232 25888 44238 25900
rect 44560 25888 44588 25987
rect 45738 25984 45744 25996
rect 45796 25984 45802 26036
rect 47118 25984 47124 26036
rect 47176 26024 47182 26036
rect 47581 26027 47639 26033
rect 47581 26024 47593 26027
rect 47176 25996 47593 26024
rect 47176 25984 47182 25996
rect 47581 25993 47593 25996
rect 47627 25993 47639 26027
rect 47581 25987 47639 25993
rect 48314 25984 48320 26036
rect 48372 25984 48378 26036
rect 49694 26024 49700 26036
rect 48700 25996 49700 26024
rect 45833 25959 45891 25965
rect 45833 25925 45845 25959
rect 45879 25956 45891 25959
rect 45922 25956 45928 25968
rect 45879 25928 45928 25956
rect 45879 25925 45891 25928
rect 45833 25919 45891 25925
rect 45922 25916 45928 25928
rect 45980 25916 45986 25968
rect 47210 25956 47216 25968
rect 47058 25928 47216 25956
rect 47210 25916 47216 25928
rect 47268 25956 47274 25968
rect 48130 25956 48136 25968
rect 47268 25928 48136 25956
rect 47268 25916 47274 25928
rect 48130 25916 48136 25928
rect 48188 25916 48194 25968
rect 48700 25900 48728 25996
rect 49694 25984 49700 25996
rect 49752 26024 49758 26036
rect 50430 26024 50436 26036
rect 49752 25996 50436 26024
rect 49752 25984 49758 25996
rect 50430 25984 50436 25996
rect 50488 26024 50494 26036
rect 52181 26027 52239 26033
rect 50488 25996 51856 26024
rect 50488 25984 50494 25996
rect 50522 25956 50528 25968
rect 48884 25928 50528 25956
rect 44232 25860 44588 25888
rect 44232 25848 44238 25860
rect 47946 25848 47952 25900
rect 48004 25888 48010 25900
rect 48501 25891 48559 25897
rect 48501 25888 48513 25891
rect 48004 25860 48513 25888
rect 48004 25848 48010 25860
rect 48501 25857 48513 25860
rect 48547 25857 48559 25891
rect 48501 25851 48559 25857
rect 48593 25891 48651 25897
rect 48593 25857 48605 25891
rect 48639 25857 48651 25891
rect 48593 25851 48651 25857
rect 43496 25792 44036 25820
rect 43496 25780 43502 25792
rect 45554 25780 45560 25832
rect 45612 25780 45618 25832
rect 47302 25780 47308 25832
rect 47360 25820 47366 25832
rect 48133 25823 48191 25829
rect 48133 25820 48145 25823
rect 47360 25792 48145 25820
rect 47360 25780 47366 25792
rect 48133 25789 48145 25792
rect 48179 25820 48191 25823
rect 48608 25820 48636 25851
rect 48682 25848 48688 25900
rect 48740 25848 48746 25900
rect 48884 25897 48912 25928
rect 50522 25916 50528 25928
rect 50580 25916 50586 25968
rect 51828 25965 51856 25996
rect 52181 25993 52193 26027
rect 52227 26024 52239 26027
rect 52638 26024 52644 26036
rect 52227 25996 52644 26024
rect 52227 25993 52239 25996
rect 52181 25987 52239 25993
rect 52638 25984 52644 25996
rect 52696 25984 52702 26036
rect 51813 25959 51871 25965
rect 51813 25925 51825 25959
rect 51859 25925 51871 25959
rect 51813 25919 51871 25925
rect 51902 25916 51908 25968
rect 51960 25916 51966 25968
rect 53006 25916 53012 25968
rect 53064 25916 53070 25968
rect 53101 25959 53159 25965
rect 53101 25925 53113 25959
rect 53147 25956 53159 25959
rect 54202 25956 54208 25968
rect 53147 25928 54208 25956
rect 53147 25925 53159 25928
rect 53101 25919 53159 25925
rect 54202 25916 54208 25928
rect 54260 25916 54266 25968
rect 56704 25928 57192 25956
rect 56704 25900 56732 25928
rect 48869 25891 48927 25897
rect 48869 25857 48881 25891
rect 48915 25857 48927 25891
rect 48869 25851 48927 25857
rect 49510 25848 49516 25900
rect 49568 25888 49574 25900
rect 49973 25891 50031 25897
rect 49973 25888 49985 25891
rect 49568 25860 49985 25888
rect 49568 25848 49574 25860
rect 49973 25857 49985 25860
rect 50019 25857 50031 25891
rect 49973 25851 50031 25857
rect 50249 25891 50307 25897
rect 50249 25857 50261 25891
rect 50295 25888 50307 25891
rect 50338 25888 50344 25900
rect 50295 25860 50344 25888
rect 50295 25857 50307 25860
rect 50249 25851 50307 25857
rect 50338 25848 50344 25860
rect 50396 25848 50402 25900
rect 51350 25848 51356 25900
rect 51408 25888 51414 25900
rect 51537 25891 51595 25897
rect 51537 25888 51549 25891
rect 51408 25860 51549 25888
rect 51408 25848 51414 25860
rect 51537 25857 51549 25860
rect 51583 25857 51595 25891
rect 51537 25851 51595 25857
rect 51626 25848 51632 25900
rect 51684 25888 51690 25900
rect 52043 25891 52101 25897
rect 51684 25860 51729 25888
rect 51684 25848 51690 25860
rect 52043 25857 52055 25891
rect 52089 25888 52101 25891
rect 52638 25888 52644 25900
rect 52089 25860 52644 25888
rect 52089 25857 52101 25860
rect 52043 25851 52101 25857
rect 52638 25848 52644 25860
rect 52696 25888 52702 25900
rect 52871 25891 52929 25897
rect 52871 25888 52883 25891
rect 52696 25860 52883 25888
rect 52696 25848 52702 25860
rect 52871 25857 52883 25860
rect 52917 25857 52929 25891
rect 53229 25891 53287 25897
rect 53229 25888 53241 25891
rect 52871 25851 52929 25857
rect 53208 25857 53241 25888
rect 53275 25857 53287 25891
rect 53208 25851 53287 25857
rect 53377 25891 53435 25897
rect 53377 25857 53389 25891
rect 53423 25888 53435 25891
rect 53466 25888 53472 25900
rect 53423 25860 53472 25888
rect 53423 25857 53435 25860
rect 53377 25851 53435 25857
rect 48179 25792 48636 25820
rect 48179 25789 48191 25792
rect 48133 25783 48191 25789
rect 49142 25780 49148 25832
rect 49200 25820 49206 25832
rect 49786 25820 49792 25832
rect 49200 25792 49792 25820
rect 49200 25780 49206 25792
rect 49786 25780 49792 25792
rect 49844 25780 49850 25832
rect 50154 25780 50160 25832
rect 50212 25780 50218 25832
rect 50706 25780 50712 25832
rect 50764 25820 50770 25832
rect 53208 25820 53236 25851
rect 53466 25848 53472 25860
rect 53524 25848 53530 25900
rect 53742 25848 53748 25900
rect 53800 25888 53806 25900
rect 53800 25860 54878 25888
rect 53800 25848 53806 25860
rect 56686 25848 56692 25900
rect 56744 25848 56750 25900
rect 56870 25848 56876 25900
rect 56928 25848 56934 25900
rect 57164 25897 57192 25928
rect 57057 25891 57115 25897
rect 57057 25857 57069 25891
rect 57103 25857 57115 25891
rect 57057 25851 57115 25857
rect 57149 25891 57207 25897
rect 57149 25857 57161 25891
rect 57195 25857 57207 25891
rect 57149 25851 57207 25857
rect 57241 25891 57299 25897
rect 57241 25857 57253 25891
rect 57287 25888 57299 25891
rect 57885 25891 57943 25897
rect 57885 25888 57897 25891
rect 57287 25860 57897 25888
rect 57287 25857 57299 25860
rect 57241 25851 57299 25857
rect 57885 25857 57897 25860
rect 57931 25857 57943 25891
rect 57885 25851 57943 25857
rect 54481 25823 54539 25829
rect 54481 25820 54493 25823
rect 50764 25792 54493 25820
rect 50764 25780 50770 25792
rect 54481 25789 54493 25792
rect 54527 25820 54539 25823
rect 55306 25820 55312 25832
rect 54527 25792 55312 25820
rect 54527 25789 54539 25792
rect 54481 25783 54539 25789
rect 55306 25780 55312 25792
rect 55364 25780 55370 25832
rect 55950 25780 55956 25832
rect 56008 25780 56014 25832
rect 56226 25780 56232 25832
rect 56284 25780 56290 25832
rect 57072 25820 57100 25851
rect 56520 25792 57100 25820
rect 49602 25752 49608 25764
rect 43119 25724 43392 25752
rect 46860 25724 49608 25752
rect 43119 25721 43131 25724
rect 43073 25715 43131 25721
rect 43806 25684 43812 25696
rect 42996 25656 43812 25684
rect 42889 25647 42947 25653
rect 43806 25644 43812 25656
rect 43864 25644 43870 25696
rect 44266 25644 44272 25696
rect 44324 25684 44330 25696
rect 44361 25687 44419 25693
rect 44361 25684 44373 25687
rect 44324 25656 44373 25684
rect 44324 25644 44330 25656
rect 44361 25653 44373 25656
rect 44407 25653 44419 25687
rect 44361 25647 44419 25653
rect 44450 25644 44456 25696
rect 44508 25684 44514 25696
rect 46860 25684 46888 25724
rect 49602 25712 49608 25724
rect 49660 25712 49666 25764
rect 50430 25712 50436 25764
rect 50488 25712 50494 25764
rect 56520 25696 56548 25792
rect 58250 25780 58256 25832
rect 58308 25820 58314 25832
rect 58437 25823 58495 25829
rect 58437 25820 58449 25823
rect 58308 25792 58449 25820
rect 58308 25780 58314 25792
rect 58437 25789 58449 25792
rect 58483 25789 58495 25823
rect 58437 25783 58495 25789
rect 44508 25656 46888 25684
rect 44508 25644 44514 25656
rect 49970 25644 49976 25696
rect 50028 25644 50034 25696
rect 51350 25644 51356 25696
rect 51408 25644 51414 25696
rect 51810 25644 51816 25696
rect 51868 25684 51874 25696
rect 52733 25687 52791 25693
rect 52733 25684 52745 25687
rect 51868 25656 52745 25684
rect 51868 25644 51874 25656
rect 52733 25653 52745 25656
rect 52779 25653 52791 25687
rect 52733 25647 52791 25653
rect 56502 25644 56508 25696
rect 56560 25644 56566 25696
rect 57514 25644 57520 25696
rect 57572 25644 57578 25696
rect 1104 25594 58880 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 58880 25594
rect 1104 25520 58880 25542
rect 17576 25483 17634 25489
rect 17576 25449 17588 25483
rect 17622 25480 17634 25483
rect 19981 25483 20039 25489
rect 19981 25480 19993 25483
rect 17622 25452 19993 25480
rect 17622 25449 17634 25452
rect 17576 25443 17634 25449
rect 19981 25449 19993 25452
rect 20027 25449 20039 25483
rect 19981 25443 20039 25449
rect 20441 25483 20499 25489
rect 20441 25449 20453 25483
rect 20487 25480 20499 25483
rect 20993 25483 21051 25489
rect 20993 25480 21005 25483
rect 20487 25452 21005 25480
rect 20487 25449 20499 25452
rect 20441 25443 20499 25449
rect 20993 25449 21005 25452
rect 21039 25480 21051 25483
rect 21542 25480 21548 25492
rect 21039 25452 21548 25480
rect 21039 25449 21051 25452
rect 20993 25443 21051 25449
rect 21542 25440 21548 25452
rect 21600 25440 21606 25492
rect 22186 25440 22192 25492
rect 22244 25480 22250 25492
rect 22370 25480 22376 25492
rect 22244 25452 22376 25480
rect 22244 25440 22250 25452
rect 22370 25440 22376 25452
rect 22428 25440 22434 25492
rect 23290 25440 23296 25492
rect 23348 25440 23354 25492
rect 25792 25452 26648 25480
rect 25038 25412 25044 25424
rect 19904 25384 20944 25412
rect 17313 25347 17371 25353
rect 17313 25313 17325 25347
rect 17359 25344 17371 25347
rect 17954 25344 17960 25356
rect 17359 25316 17960 25344
rect 17359 25313 17371 25316
rect 17313 25307 17371 25313
rect 17954 25304 17960 25316
rect 18012 25304 18018 25356
rect 19061 25347 19119 25353
rect 19061 25313 19073 25347
rect 19107 25344 19119 25347
rect 19107 25316 19840 25344
rect 19107 25313 19119 25316
rect 19061 25307 19119 25313
rect 19518 25236 19524 25288
rect 19576 25236 19582 25288
rect 19426 25208 19432 25220
rect 18814 25180 19432 25208
rect 19426 25168 19432 25180
rect 19484 25168 19490 25220
rect 19610 25168 19616 25220
rect 19668 25168 19674 25220
rect 19702 25168 19708 25220
rect 19760 25168 19766 25220
rect 19812 25208 19840 25316
rect 19904 25285 19932 25384
rect 19995 25316 20392 25344
rect 19889 25279 19947 25285
rect 19889 25245 19901 25279
rect 19935 25245 19947 25279
rect 19889 25239 19947 25245
rect 19995 25208 20023 25316
rect 20162 25236 20168 25288
rect 20220 25236 20226 25288
rect 20257 25279 20315 25285
rect 20257 25245 20269 25279
rect 20303 25245 20315 25279
rect 20364 25276 20392 25316
rect 20916 25288 20944 25384
rect 23676 25384 25044 25412
rect 21453 25347 21511 25353
rect 21453 25313 21465 25347
rect 21499 25344 21511 25347
rect 21818 25344 21824 25356
rect 21499 25316 21824 25344
rect 21499 25313 21511 25316
rect 21453 25307 21511 25313
rect 21818 25304 21824 25316
rect 21876 25304 21882 25356
rect 23201 25347 23259 25353
rect 23201 25313 23213 25347
rect 23247 25344 23259 25347
rect 23382 25344 23388 25356
rect 23247 25316 23388 25344
rect 23247 25313 23259 25316
rect 23201 25307 23259 25313
rect 23382 25304 23388 25316
rect 23440 25304 23446 25356
rect 20530 25276 20536 25288
rect 20364 25248 20536 25276
rect 20257 25239 20315 25245
rect 19812 25180 20023 25208
rect 19337 25143 19395 25149
rect 19337 25109 19349 25143
rect 19383 25140 19395 25143
rect 20272 25140 20300 25239
rect 20530 25236 20536 25248
rect 20588 25236 20594 25288
rect 20898 25236 20904 25288
rect 20956 25236 20962 25288
rect 21174 25236 21180 25288
rect 21232 25236 21238 25288
rect 23290 25236 23296 25288
rect 23348 25276 23354 25288
rect 23474 25285 23480 25288
rect 23472 25276 23480 25285
rect 23348 25248 23480 25276
rect 23348 25236 23354 25248
rect 23472 25239 23480 25248
rect 23474 25236 23480 25239
rect 23532 25236 23538 25288
rect 21729 25211 21787 25217
rect 21729 25177 21741 25211
rect 21775 25208 21787 25211
rect 22002 25208 22008 25220
rect 21775 25180 22008 25208
rect 21775 25177 21787 25180
rect 21729 25171 21787 25177
rect 22002 25168 22008 25180
rect 22060 25168 22066 25220
rect 23014 25208 23020 25220
rect 22954 25180 23020 25208
rect 23014 25168 23020 25180
rect 23072 25168 23078 25220
rect 23566 25168 23572 25220
rect 23624 25168 23630 25220
rect 23676 25217 23704 25384
rect 25038 25372 25044 25384
rect 25096 25412 25102 25424
rect 25222 25412 25228 25424
rect 25096 25384 25228 25412
rect 25096 25372 25102 25384
rect 25222 25372 25228 25384
rect 25280 25372 25286 25424
rect 24946 25344 24952 25356
rect 23860 25316 24952 25344
rect 23860 25285 23888 25316
rect 24946 25304 24952 25316
rect 25004 25344 25010 25356
rect 25682 25344 25688 25356
rect 25004 25316 25688 25344
rect 25004 25304 25010 25316
rect 25682 25304 25688 25316
rect 25740 25304 25746 25356
rect 23844 25279 23902 25285
rect 23844 25245 23856 25279
rect 23890 25245 23902 25279
rect 23844 25239 23902 25245
rect 23937 25279 23995 25285
rect 23937 25245 23949 25279
rect 23983 25276 23995 25279
rect 23983 25248 24164 25276
rect 23983 25245 23995 25248
rect 23937 25239 23995 25245
rect 23661 25211 23719 25217
rect 23661 25177 23673 25211
rect 23707 25177 23719 25211
rect 23661 25171 23719 25177
rect 19383 25112 20300 25140
rect 21361 25143 21419 25149
rect 19383 25109 19395 25112
rect 19337 25103 19395 25109
rect 21361 25109 21373 25143
rect 21407 25140 21419 25143
rect 22370 25140 22376 25152
rect 21407 25112 22376 25140
rect 21407 25109 21419 25112
rect 21361 25103 21419 25109
rect 22370 25100 22376 25112
rect 22428 25100 22434 25152
rect 23290 25100 23296 25152
rect 23348 25140 23354 25152
rect 23676 25140 23704 25171
rect 24136 25149 24164 25248
rect 25222 25236 25228 25288
rect 25280 25276 25286 25288
rect 25792 25285 25820 25452
rect 26234 25372 26240 25424
rect 26292 25372 26298 25424
rect 26620 25421 26648 25452
rect 28810 25440 28816 25492
rect 28868 25480 28874 25492
rect 28905 25483 28963 25489
rect 28905 25480 28917 25483
rect 28868 25452 28917 25480
rect 28868 25440 28874 25452
rect 28905 25449 28917 25452
rect 28951 25449 28963 25483
rect 28905 25443 28963 25449
rect 31846 25440 31852 25492
rect 31904 25480 31910 25492
rect 34330 25480 34336 25492
rect 31904 25452 34336 25480
rect 31904 25440 31910 25452
rect 34330 25440 34336 25452
rect 34388 25440 34394 25492
rect 36262 25440 36268 25492
rect 36320 25480 36326 25492
rect 36495 25483 36553 25489
rect 36495 25480 36507 25483
rect 36320 25452 36507 25480
rect 36320 25440 36326 25452
rect 36495 25449 36507 25452
rect 36541 25480 36553 25483
rect 38930 25480 38936 25492
rect 36541 25452 36952 25480
rect 36541 25449 36553 25452
rect 36495 25443 36553 25449
rect 26605 25415 26663 25421
rect 26605 25381 26617 25415
rect 26651 25412 26663 25415
rect 30190 25412 30196 25424
rect 26651 25384 30196 25412
rect 26651 25381 26663 25384
rect 26605 25375 26663 25381
rect 30190 25372 30196 25384
rect 30248 25372 30254 25424
rect 32858 25372 32864 25424
rect 32916 25412 32922 25424
rect 33505 25415 33563 25421
rect 33505 25412 33517 25415
rect 32916 25384 33517 25412
rect 32916 25372 32922 25384
rect 33505 25381 33517 25384
rect 33551 25381 33563 25415
rect 33505 25375 33563 25381
rect 26252 25344 26280 25372
rect 26160 25316 26280 25344
rect 26421 25347 26479 25353
rect 26160 25285 26188 25316
rect 26421 25313 26433 25347
rect 26467 25344 26479 25347
rect 26467 25316 29684 25344
rect 26467 25313 26479 25316
rect 26421 25307 26479 25313
rect 25772 25279 25830 25285
rect 25772 25276 25784 25279
rect 25280 25248 25784 25276
rect 25280 25236 25286 25248
rect 25772 25245 25784 25248
rect 25818 25245 25830 25279
rect 25772 25239 25830 25245
rect 25869 25279 25927 25285
rect 25869 25245 25881 25279
rect 25915 25245 25927 25279
rect 25869 25239 25927 25245
rect 26144 25279 26202 25285
rect 26144 25245 26156 25279
rect 26190 25245 26202 25279
rect 26144 25239 26202 25245
rect 26237 25279 26295 25285
rect 26237 25245 26249 25279
rect 26283 25276 26295 25279
rect 26436 25276 26464 25307
rect 26283 25248 26464 25276
rect 26283 25245 26295 25248
rect 26237 25239 26295 25245
rect 25406 25168 25412 25220
rect 25464 25208 25470 25220
rect 25884 25208 25912 25239
rect 28350 25236 28356 25288
rect 28408 25236 28414 25288
rect 28442 25236 28448 25288
rect 28500 25276 28506 25288
rect 28721 25279 28779 25285
rect 28721 25276 28733 25279
rect 28500 25248 28733 25276
rect 28500 25236 28506 25248
rect 28721 25245 28733 25248
rect 28767 25245 28779 25279
rect 28721 25239 28779 25245
rect 28810 25236 28816 25288
rect 28868 25276 28874 25288
rect 29273 25279 29331 25285
rect 29273 25276 29285 25279
rect 28868 25248 29285 25276
rect 28868 25236 28874 25248
rect 29273 25245 29285 25248
rect 29319 25276 29331 25279
rect 29549 25279 29607 25285
rect 29549 25276 29561 25279
rect 29319 25248 29561 25276
rect 29319 25245 29331 25248
rect 29273 25239 29331 25245
rect 29549 25245 29561 25248
rect 29595 25245 29607 25279
rect 29549 25239 29607 25245
rect 25464 25180 25912 25208
rect 25961 25211 26019 25217
rect 25464 25168 25470 25180
rect 25961 25177 25973 25211
rect 26007 25208 26019 25211
rect 26007 25180 26832 25208
rect 26007 25177 26019 25180
rect 25961 25171 26019 25177
rect 23348 25112 23704 25140
rect 24121 25143 24179 25149
rect 23348 25100 23354 25112
rect 24121 25109 24133 25143
rect 24167 25140 24179 25143
rect 24210 25140 24216 25152
rect 24167 25112 24216 25140
rect 24167 25109 24179 25112
rect 24121 25103 24179 25109
rect 24210 25100 24216 25112
rect 24268 25100 24274 25152
rect 25593 25143 25651 25149
rect 25593 25109 25605 25143
rect 25639 25140 25651 25143
rect 26050 25140 26056 25152
rect 25639 25112 26056 25140
rect 25639 25109 25651 25112
rect 25593 25103 25651 25109
rect 26050 25100 26056 25112
rect 26108 25100 26114 25152
rect 26804 25149 26832 25180
rect 27706 25168 27712 25220
rect 27764 25208 27770 25220
rect 28537 25211 28595 25217
rect 28537 25208 28549 25211
rect 27764 25180 28549 25208
rect 27764 25168 27770 25180
rect 28537 25177 28549 25180
rect 28583 25177 28595 25211
rect 28537 25171 28595 25177
rect 28626 25168 28632 25220
rect 28684 25168 28690 25220
rect 26789 25143 26847 25149
rect 26789 25109 26801 25143
rect 26835 25140 26847 25143
rect 27338 25140 27344 25152
rect 26835 25112 27344 25140
rect 26835 25109 26847 25112
rect 26789 25103 26847 25109
rect 27338 25100 27344 25112
rect 27396 25100 27402 25152
rect 28166 25100 28172 25152
rect 28224 25140 28230 25152
rect 29089 25143 29147 25149
rect 29089 25140 29101 25143
rect 28224 25112 29101 25140
rect 28224 25100 28230 25112
rect 29089 25109 29101 25112
rect 29135 25109 29147 25143
rect 29656 25140 29684 25316
rect 30558 25304 30564 25356
rect 30616 25344 30622 25356
rect 31113 25347 31171 25353
rect 31113 25344 31125 25347
rect 30616 25316 31125 25344
rect 30616 25304 30622 25316
rect 31113 25313 31125 25316
rect 31159 25313 31171 25347
rect 31113 25307 31171 25313
rect 31481 25347 31539 25353
rect 31481 25313 31493 25347
rect 31527 25344 31539 25347
rect 33045 25347 33103 25353
rect 33045 25344 33057 25347
rect 31527 25316 33057 25344
rect 31527 25313 31539 25316
rect 31481 25307 31539 25313
rect 33045 25313 33057 25316
rect 33091 25313 33103 25347
rect 33045 25307 33103 25313
rect 34701 25347 34759 25353
rect 34701 25313 34713 25347
rect 34747 25344 34759 25347
rect 34974 25344 34980 25356
rect 34747 25316 34980 25344
rect 34747 25313 34759 25316
rect 34701 25307 34759 25313
rect 34974 25304 34980 25316
rect 35032 25344 35038 25356
rect 36814 25344 36820 25356
rect 35032 25316 36820 25344
rect 35032 25304 35038 25316
rect 36814 25304 36820 25316
rect 36872 25304 36878 25356
rect 36924 25344 36952 25452
rect 38626 25452 38936 25480
rect 37185 25415 37243 25421
rect 37185 25381 37197 25415
rect 37231 25412 37243 25415
rect 37458 25412 37464 25424
rect 37231 25384 37464 25412
rect 37231 25381 37243 25384
rect 37185 25375 37243 25381
rect 37458 25372 37464 25384
rect 37516 25372 37522 25424
rect 37090 25344 37096 25356
rect 36924 25316 37096 25344
rect 33226 25236 33232 25288
rect 33284 25236 33290 25288
rect 33318 25236 33324 25288
rect 33376 25236 33382 25288
rect 33597 25279 33655 25285
rect 33597 25245 33609 25279
rect 33643 25245 33655 25279
rect 33597 25239 33655 25245
rect 32214 25168 32220 25220
rect 32272 25168 32278 25220
rect 32907 25211 32965 25217
rect 32907 25177 32919 25211
rect 32953 25208 32965 25211
rect 33042 25208 33048 25220
rect 32953 25180 33048 25208
rect 32953 25177 32965 25180
rect 32907 25171 32965 25177
rect 33042 25168 33048 25180
rect 33100 25208 33106 25220
rect 33612 25208 33640 25239
rect 35066 25236 35072 25288
rect 35124 25236 35130 25288
rect 35986 25236 35992 25288
rect 36044 25276 36050 25288
rect 36924 25285 36952 25316
rect 37090 25304 37096 25316
rect 37148 25304 37154 25356
rect 37734 25304 37740 25356
rect 37792 25344 37798 25356
rect 38197 25347 38255 25353
rect 37792 25316 37964 25344
rect 37792 25304 37798 25316
rect 36633 25279 36691 25285
rect 36633 25276 36645 25279
rect 36044 25248 36645 25276
rect 36044 25236 36050 25248
rect 36633 25245 36645 25248
rect 36679 25245 36691 25279
rect 36633 25239 36691 25245
rect 36909 25279 36967 25285
rect 36909 25245 36921 25279
rect 36955 25245 36967 25279
rect 36909 25239 36967 25245
rect 36998 25236 37004 25288
rect 37056 25236 37062 25288
rect 37182 25236 37188 25288
rect 37240 25276 37246 25288
rect 37829 25279 37887 25285
rect 37829 25276 37841 25279
rect 37240 25248 37841 25276
rect 37240 25236 37246 25248
rect 37829 25245 37841 25248
rect 37875 25245 37887 25279
rect 37829 25239 37887 25245
rect 33100 25180 33640 25208
rect 33100 25168 33106 25180
rect 36078 25168 36084 25220
rect 36136 25208 36142 25220
rect 36538 25208 36544 25220
rect 36136 25180 36544 25208
rect 36136 25168 36142 25180
rect 36538 25168 36544 25180
rect 36596 25168 36602 25220
rect 36814 25168 36820 25220
rect 36872 25208 36878 25220
rect 37461 25211 37519 25217
rect 37461 25208 37473 25211
rect 36872 25180 37473 25208
rect 36872 25168 36878 25180
rect 37461 25177 37473 25180
rect 37507 25208 37519 25211
rect 37642 25208 37648 25220
rect 37507 25180 37648 25208
rect 37507 25177 37519 25180
rect 37461 25171 37519 25177
rect 37642 25168 37648 25180
rect 37700 25168 37706 25220
rect 37936 25208 37964 25316
rect 38197 25313 38209 25347
rect 38243 25344 38255 25347
rect 38626 25344 38654 25452
rect 38930 25440 38936 25452
rect 38988 25480 38994 25492
rect 40218 25480 40224 25492
rect 38988 25452 40224 25480
rect 38988 25440 38994 25452
rect 40218 25440 40224 25452
rect 40276 25440 40282 25492
rect 41506 25440 41512 25492
rect 41564 25480 41570 25492
rect 41601 25483 41659 25489
rect 41601 25480 41613 25483
rect 41564 25452 41613 25480
rect 41564 25440 41570 25452
rect 41601 25449 41613 25452
rect 41647 25480 41659 25483
rect 42702 25480 42708 25492
rect 41647 25452 42708 25480
rect 41647 25449 41659 25452
rect 41601 25443 41659 25449
rect 42702 25440 42708 25452
rect 42760 25440 42766 25492
rect 42981 25483 43039 25489
rect 42981 25449 42993 25483
rect 43027 25449 43039 25483
rect 42981 25443 43039 25449
rect 38838 25372 38844 25424
rect 38896 25412 38902 25424
rect 39393 25415 39451 25421
rect 39393 25412 39405 25415
rect 38896 25384 39405 25412
rect 38896 25372 38902 25384
rect 39393 25381 39405 25384
rect 39439 25381 39451 25415
rect 39393 25375 39451 25381
rect 41785 25415 41843 25421
rect 41785 25381 41797 25415
rect 41831 25412 41843 25415
rect 42521 25415 42579 25421
rect 42521 25412 42533 25415
rect 41831 25384 42533 25412
rect 41831 25381 41843 25384
rect 41785 25375 41843 25381
rect 42521 25381 42533 25384
rect 42567 25381 42579 25415
rect 42521 25375 42579 25381
rect 38243 25316 38654 25344
rect 38243 25313 38255 25316
rect 38197 25307 38255 25313
rect 39482 25304 39488 25356
rect 39540 25344 39546 25356
rect 39540 25316 40172 25344
rect 39540 25304 39546 25316
rect 38654 25285 38660 25288
rect 38105 25279 38163 25285
rect 38105 25245 38117 25279
rect 38151 25276 38163 25279
rect 38652 25276 38660 25285
rect 38151 25248 38660 25276
rect 38151 25245 38163 25248
rect 38105 25239 38163 25245
rect 38652 25239 38660 25248
rect 38654 25236 38660 25239
rect 38712 25236 38718 25288
rect 38746 25236 38752 25288
rect 38804 25236 38810 25288
rect 39022 25236 39028 25288
rect 39080 25236 39086 25288
rect 39114 25236 39120 25288
rect 39172 25236 39178 25288
rect 39390 25276 39396 25288
rect 39224 25248 39396 25276
rect 37936 25180 38608 25208
rect 31754 25140 31760 25152
rect 29656 25112 31760 25140
rect 29089 25103 29147 25109
rect 31754 25100 31760 25112
rect 31812 25100 31818 25152
rect 32030 25100 32036 25152
rect 32088 25140 32094 25152
rect 33226 25140 33232 25152
rect 32088 25112 33232 25140
rect 32088 25100 32094 25112
rect 33226 25100 33232 25112
rect 33284 25100 33290 25152
rect 36998 25100 37004 25152
rect 37056 25140 37062 25152
rect 37277 25143 37335 25149
rect 37277 25140 37289 25143
rect 37056 25112 37289 25140
rect 37056 25100 37062 25112
rect 37277 25109 37289 25112
rect 37323 25109 37335 25143
rect 37277 25103 37335 25109
rect 37550 25100 37556 25152
rect 37608 25140 37614 25152
rect 38381 25143 38439 25149
rect 38381 25140 38393 25143
rect 37608 25112 38393 25140
rect 37608 25100 37614 25112
rect 38381 25109 38393 25112
rect 38427 25109 38439 25143
rect 38381 25103 38439 25109
rect 38470 25100 38476 25152
rect 38528 25100 38534 25152
rect 38580 25140 38608 25180
rect 38838 25168 38844 25220
rect 38896 25168 38902 25220
rect 39224 25149 39252 25248
rect 39390 25236 39396 25248
rect 39448 25276 39454 25288
rect 39850 25276 39856 25288
rect 39448 25248 39856 25276
rect 39448 25236 39454 25248
rect 39850 25236 39856 25248
rect 39908 25236 39914 25288
rect 40034 25285 40040 25288
rect 40012 25279 40040 25285
rect 40012 25245 40024 25279
rect 40012 25239 40040 25245
rect 40034 25236 40040 25239
rect 40092 25236 40098 25288
rect 40144 25285 40172 25316
rect 40310 25304 40316 25356
rect 40368 25344 40374 25356
rect 40497 25347 40555 25353
rect 40497 25344 40509 25347
rect 40368 25316 40509 25344
rect 40368 25304 40374 25316
rect 40497 25313 40509 25316
rect 40543 25344 40555 25347
rect 41230 25344 41236 25356
rect 40543 25316 41236 25344
rect 40543 25313 40555 25316
rect 40497 25307 40555 25313
rect 41230 25304 41236 25316
rect 41288 25304 41294 25356
rect 41966 25304 41972 25356
rect 42024 25304 42030 25356
rect 42058 25304 42064 25356
rect 42116 25304 42122 25356
rect 42153 25347 42211 25353
rect 42153 25313 42165 25347
rect 42199 25344 42211 25347
rect 42334 25344 42340 25356
rect 42199 25316 42340 25344
rect 42199 25313 42211 25316
rect 42153 25307 42211 25313
rect 42334 25304 42340 25316
rect 42392 25304 42398 25356
rect 42536 25344 42564 25375
rect 42794 25372 42800 25424
rect 42852 25412 42858 25424
rect 42996 25412 43024 25443
rect 43346 25440 43352 25492
rect 43404 25440 43410 25492
rect 43806 25440 43812 25492
rect 43864 25440 43870 25492
rect 43990 25440 43996 25492
rect 44048 25480 44054 25492
rect 44048 25452 48176 25480
rect 44048 25440 44054 25452
rect 44269 25415 44327 25421
rect 44269 25412 44281 25415
rect 42852 25384 44281 25412
rect 42852 25372 42858 25384
rect 44269 25381 44281 25384
rect 44315 25412 44327 25415
rect 44450 25412 44456 25424
rect 44315 25384 44456 25412
rect 44315 25381 44327 25384
rect 44269 25375 44327 25381
rect 44450 25372 44456 25384
rect 44508 25372 44514 25424
rect 48148 25412 48176 25452
rect 48222 25440 48228 25492
rect 48280 25440 48286 25492
rect 50154 25440 50160 25492
rect 50212 25440 50218 25492
rect 52638 25440 52644 25492
rect 52696 25480 52702 25492
rect 52696 25452 54248 25480
rect 52696 25440 52702 25452
rect 49605 25415 49663 25421
rect 48148 25384 49556 25412
rect 42536 25316 43576 25344
rect 41325 25289 41383 25295
rect 40129 25279 40187 25285
rect 40129 25245 40141 25279
rect 40175 25276 40187 25279
rect 41325 25276 41337 25289
rect 40175 25255 41337 25276
rect 41371 25276 41383 25289
rect 42245 25279 42303 25285
rect 41371 25255 41676 25276
rect 40175 25248 41676 25255
rect 40175 25245 40187 25248
rect 40129 25239 40187 25245
rect 39666 25168 39672 25220
rect 39724 25208 39730 25220
rect 40221 25211 40279 25217
rect 40221 25208 40233 25211
rect 39724 25180 40233 25208
rect 39724 25168 39730 25180
rect 40221 25177 40233 25180
rect 40267 25208 40279 25211
rect 40267 25180 41368 25208
rect 40267 25177 40279 25180
rect 40221 25171 40279 25177
rect 39209 25143 39267 25149
rect 39209 25140 39221 25143
rect 38580 25112 39221 25140
rect 39209 25109 39221 25112
rect 39255 25109 39267 25143
rect 39209 25103 39267 25109
rect 39298 25100 39304 25152
rect 39356 25140 39362 25152
rect 39853 25143 39911 25149
rect 39853 25140 39865 25143
rect 39356 25112 39865 25140
rect 39356 25100 39362 25112
rect 39853 25109 39865 25112
rect 39899 25109 39911 25143
rect 39853 25103 39911 25109
rect 40954 25100 40960 25152
rect 41012 25140 41018 25152
rect 41233 25143 41291 25149
rect 41233 25140 41245 25143
rect 41012 25112 41245 25140
rect 41012 25100 41018 25112
rect 41233 25109 41245 25112
rect 41279 25109 41291 25143
rect 41340 25140 41368 25180
rect 41414 25168 41420 25220
rect 41472 25168 41478 25220
rect 41648 25217 41676 25248
rect 42245 25245 42257 25279
rect 42291 25276 42303 25279
rect 42518 25276 42524 25288
rect 42291 25248 42524 25276
rect 42291 25245 42303 25248
rect 42245 25239 42303 25245
rect 42518 25236 42524 25248
rect 42576 25236 42582 25288
rect 42797 25279 42855 25285
rect 42797 25245 42809 25279
rect 42843 25276 42855 25279
rect 42886 25276 42892 25288
rect 42843 25248 42892 25276
rect 42843 25245 42855 25248
rect 42797 25239 42855 25245
rect 42886 25236 42892 25248
rect 42944 25236 42950 25288
rect 43548 25285 43576 25316
rect 43806 25304 43812 25356
rect 43864 25344 43870 25356
rect 44361 25347 44419 25353
rect 44361 25344 44373 25347
rect 43864 25316 44373 25344
rect 43864 25304 43870 25316
rect 44361 25313 44373 25316
rect 44407 25313 44419 25347
rect 44361 25307 44419 25313
rect 43533 25279 43591 25285
rect 43533 25245 43545 25279
rect 43579 25245 43591 25279
rect 43533 25239 43591 25245
rect 43622 25236 43628 25288
rect 43680 25236 43686 25288
rect 41633 25211 41691 25217
rect 41633 25177 41645 25211
rect 41679 25208 41691 25211
rect 42610 25208 42616 25220
rect 41679 25180 42616 25208
rect 41679 25177 41691 25180
rect 41633 25171 41691 25177
rect 42610 25168 42616 25180
rect 42668 25168 42674 25220
rect 42702 25168 42708 25220
rect 42760 25168 42766 25220
rect 41506 25140 41512 25152
rect 41340 25112 41512 25140
rect 41233 25103 41291 25109
rect 41506 25100 41512 25112
rect 41564 25100 41570 25152
rect 42429 25143 42487 25149
rect 42429 25109 42441 25143
rect 42475 25140 42487 25143
rect 43990 25140 43996 25152
rect 42475 25112 43996 25140
rect 42475 25109 42487 25112
rect 42429 25103 42487 25109
rect 43990 25100 43996 25112
rect 44048 25100 44054 25152
rect 44376 25140 44404 25307
rect 46474 25304 46480 25356
rect 46532 25344 46538 25356
rect 47489 25347 47547 25353
rect 47489 25344 47501 25347
rect 46532 25316 47501 25344
rect 46532 25304 46538 25316
rect 47489 25313 47501 25316
rect 47535 25313 47547 25347
rect 47489 25307 47547 25313
rect 47946 25304 47952 25356
rect 48004 25344 48010 25356
rect 49528 25344 49556 25384
rect 49605 25381 49617 25415
rect 49651 25412 49663 25415
rect 50246 25412 50252 25424
rect 49651 25384 50252 25412
rect 49651 25381 49663 25384
rect 49605 25375 49663 25381
rect 50246 25372 50252 25384
rect 50304 25372 50310 25424
rect 50351 25384 50844 25412
rect 50351 25344 50379 25384
rect 48004 25316 48314 25344
rect 48004 25304 48010 25316
rect 45646 25236 45652 25288
rect 45704 25236 45710 25288
rect 48041 25279 48099 25285
rect 48041 25276 48053 25279
rect 47780 25248 48053 25276
rect 45922 25168 45928 25220
rect 45980 25168 45986 25220
rect 47210 25208 47216 25220
rect 47150 25180 47216 25208
rect 47210 25168 47216 25180
rect 47268 25208 47274 25220
rect 47486 25208 47492 25220
rect 47268 25180 47492 25208
rect 47268 25168 47274 25180
rect 47486 25168 47492 25180
rect 47544 25168 47550 25220
rect 47780 25152 47808 25248
rect 48041 25245 48053 25248
rect 48087 25245 48099 25279
rect 48286 25276 48314 25316
rect 48791 25316 49372 25344
rect 49528 25316 50379 25344
rect 48791 25285 48819 25316
rect 49344 25288 49372 25316
rect 48363 25279 48421 25285
rect 48363 25276 48375 25279
rect 48286 25248 48375 25276
rect 48041 25239 48099 25245
rect 48363 25245 48375 25248
rect 48409 25245 48421 25279
rect 48363 25239 48421 25245
rect 48776 25279 48834 25285
rect 48776 25245 48788 25279
rect 48822 25245 48834 25279
rect 48776 25239 48834 25245
rect 48869 25279 48927 25285
rect 48869 25245 48881 25279
rect 48915 25276 48927 25279
rect 48958 25276 48964 25288
rect 48915 25248 48964 25276
rect 48915 25245 48927 25248
rect 48869 25239 48927 25245
rect 48056 25208 48084 25239
rect 48958 25236 48964 25248
rect 49016 25236 49022 25288
rect 49053 25279 49111 25285
rect 49053 25245 49065 25279
rect 49099 25276 49111 25279
rect 49142 25276 49148 25288
rect 49099 25248 49148 25276
rect 49099 25245 49111 25248
rect 49053 25239 49111 25245
rect 49142 25236 49148 25248
rect 49200 25236 49206 25288
rect 49326 25236 49332 25288
rect 49384 25236 49390 25288
rect 49418 25236 49424 25288
rect 49476 25276 49482 25288
rect 49697 25279 49755 25285
rect 49697 25276 49709 25279
rect 49476 25248 49709 25276
rect 49476 25236 49482 25248
rect 49697 25245 49709 25248
rect 49743 25245 49755 25279
rect 49697 25239 49755 25245
rect 50154 25236 50160 25288
rect 50212 25276 50218 25288
rect 50295 25279 50353 25285
rect 50295 25276 50307 25279
rect 50212 25248 50307 25276
rect 50212 25236 50218 25248
rect 50295 25245 50307 25248
rect 50341 25245 50353 25279
rect 50295 25239 50353 25245
rect 50433 25279 50491 25285
rect 50433 25245 50445 25279
rect 50479 25276 50491 25279
rect 50614 25276 50620 25288
rect 50479 25248 50620 25276
rect 50479 25245 50491 25248
rect 50433 25239 50491 25245
rect 50614 25236 50620 25248
rect 50672 25236 50678 25288
rect 50706 25236 50712 25288
rect 50764 25236 50770 25288
rect 50816 25285 50844 25384
rect 52104 25384 52316 25412
rect 52104 25353 52132 25384
rect 52089 25347 52147 25353
rect 52089 25313 52101 25347
rect 52135 25313 52147 25347
rect 52089 25307 52147 25313
rect 52178 25304 52184 25356
rect 52236 25304 52242 25356
rect 52288 25344 52316 25384
rect 52822 25344 52828 25356
rect 52288 25316 52828 25344
rect 52822 25304 52828 25316
rect 52880 25304 52886 25356
rect 53466 25304 53472 25356
rect 53524 25344 53530 25356
rect 53524 25316 54064 25344
rect 53524 25304 53530 25316
rect 50801 25279 50859 25285
rect 50801 25245 50813 25279
rect 50847 25245 50859 25279
rect 50801 25239 50859 25245
rect 51810 25236 51816 25288
rect 51868 25236 51874 25288
rect 51994 25236 52000 25288
rect 52052 25236 52058 25288
rect 54036 25285 54064 25316
rect 54021 25279 54079 25285
rect 54021 25245 54033 25279
rect 54067 25245 54079 25279
rect 54021 25239 54079 25245
rect 54114 25279 54172 25285
rect 54114 25245 54126 25279
rect 54160 25245 54172 25279
rect 54220 25276 54248 25452
rect 55950 25440 55956 25492
rect 56008 25480 56014 25492
rect 56045 25483 56103 25489
rect 56045 25480 56057 25483
rect 56008 25452 56057 25480
rect 56008 25440 56014 25452
rect 56045 25449 56057 25452
rect 56091 25449 56103 25483
rect 56045 25443 56103 25449
rect 58250 25440 58256 25492
rect 58308 25440 58314 25492
rect 54665 25415 54723 25421
rect 54665 25381 54677 25415
rect 54711 25381 54723 25415
rect 54665 25375 54723 25381
rect 54680 25344 54708 25375
rect 56226 25372 56232 25424
rect 56284 25372 56290 25424
rect 56244 25344 56272 25372
rect 56873 25347 56931 25353
rect 56873 25344 56885 25347
rect 54680 25316 55536 25344
rect 56244 25316 56885 25344
rect 54486 25279 54544 25285
rect 54486 25276 54498 25279
rect 54220 25248 54498 25276
rect 54114 25239 54172 25245
rect 54486 25245 54498 25248
rect 54532 25276 54544 25279
rect 54532 25248 54708 25276
rect 54532 25245 54544 25248
rect 54486 25239 54544 25245
rect 48501 25211 48559 25217
rect 48501 25208 48513 25211
rect 48056 25180 48513 25208
rect 48501 25177 48513 25180
rect 48547 25177 48559 25211
rect 48501 25171 48559 25177
rect 48590 25168 48596 25220
rect 48648 25168 48654 25220
rect 49237 25211 49295 25217
rect 49237 25177 49249 25211
rect 49283 25177 49295 25211
rect 49237 25171 49295 25177
rect 50525 25211 50583 25217
rect 50525 25177 50537 25211
rect 50571 25177 50583 25211
rect 50525 25171 50583 25177
rect 51629 25211 51687 25217
rect 51629 25177 51641 25211
rect 51675 25208 51687 25211
rect 52457 25211 52515 25217
rect 52457 25208 52469 25211
rect 51675 25180 52469 25208
rect 51675 25177 51687 25180
rect 51629 25171 51687 25177
rect 52457 25177 52469 25180
rect 52503 25177 52515 25211
rect 53742 25208 53748 25220
rect 53682 25180 53748 25208
rect 52457 25171 52515 25177
rect 46934 25140 46940 25152
rect 44376 25112 46940 25140
rect 46934 25100 46940 25112
rect 46992 25100 46998 25152
rect 47397 25143 47455 25149
rect 47397 25109 47409 25143
rect 47443 25140 47455 25143
rect 47762 25140 47768 25152
rect 47443 25112 47768 25140
rect 47443 25109 47455 25112
rect 47397 25103 47455 25109
rect 47762 25100 47768 25112
rect 47820 25100 47826 25152
rect 48774 25100 48780 25152
rect 48832 25140 48838 25152
rect 49252 25140 49280 25171
rect 48832 25112 49280 25140
rect 48832 25100 48838 25112
rect 49786 25100 49792 25152
rect 49844 25140 49850 25152
rect 49881 25143 49939 25149
rect 49881 25140 49893 25143
rect 49844 25112 49893 25140
rect 49844 25100 49850 25112
rect 49881 25109 49893 25112
rect 49927 25140 49939 25143
rect 50540 25140 50568 25171
rect 53742 25168 53748 25180
rect 53800 25168 53806 25220
rect 53834 25168 53840 25220
rect 53892 25208 53898 25220
rect 54129 25208 54157 25239
rect 53892 25180 54157 25208
rect 53892 25168 53898 25180
rect 54202 25168 54208 25220
rect 54260 25208 54266 25220
rect 54297 25211 54355 25217
rect 54297 25208 54309 25211
rect 54260 25180 54309 25208
rect 54260 25168 54266 25180
rect 54297 25177 54309 25180
rect 54343 25177 54355 25211
rect 54297 25171 54355 25177
rect 54389 25211 54447 25217
rect 54389 25177 54401 25211
rect 54435 25177 54447 25211
rect 54680 25208 54708 25248
rect 55306 25236 55312 25288
rect 55364 25236 55370 25288
rect 55508 25276 55536 25316
rect 56873 25313 56885 25316
rect 56919 25313 56931 25347
rect 56873 25307 56931 25313
rect 56229 25279 56287 25285
rect 56229 25276 56241 25279
rect 55508 25248 56241 25276
rect 56229 25245 56241 25248
rect 56275 25245 56287 25279
rect 56229 25239 56287 25245
rect 56410 25236 56416 25288
rect 56468 25236 56474 25288
rect 56505 25279 56563 25285
rect 56505 25245 56517 25279
rect 56551 25245 56563 25279
rect 56505 25239 56563 25245
rect 57140 25279 57198 25285
rect 57140 25245 57152 25279
rect 57186 25276 57198 25279
rect 57514 25276 57520 25288
rect 57186 25248 57520 25276
rect 57186 25245 57198 25248
rect 57140 25239 57198 25245
rect 55674 25208 55680 25220
rect 54680 25180 55680 25208
rect 54389 25171 54447 25177
rect 49927 25112 50568 25140
rect 49927 25109 49939 25112
rect 49881 25103 49939 25109
rect 50798 25100 50804 25152
rect 50856 25140 50862 25152
rect 50893 25143 50951 25149
rect 50893 25140 50905 25143
rect 50856 25112 50905 25140
rect 50856 25100 50862 25112
rect 50893 25109 50905 25112
rect 50939 25109 50951 25143
rect 50893 25103 50951 25109
rect 53374 25100 53380 25152
rect 53432 25140 53438 25152
rect 53929 25143 53987 25149
rect 53929 25140 53941 25143
rect 53432 25112 53941 25140
rect 53432 25100 53438 25112
rect 53929 25109 53941 25112
rect 53975 25140 53987 25143
rect 54404 25140 54432 25171
rect 55674 25168 55680 25180
rect 55732 25168 55738 25220
rect 55953 25211 56011 25217
rect 55953 25177 55965 25211
rect 55999 25208 56011 25211
rect 56520 25208 56548 25239
rect 57514 25236 57520 25248
rect 57572 25236 57578 25288
rect 55999 25180 56548 25208
rect 55999 25177 56011 25180
rect 55953 25171 56011 25177
rect 53975 25112 54432 25140
rect 53975 25109 53987 25112
rect 53929 25103 53987 25109
rect 1104 25050 58880 25072
rect 1104 24998 4874 25050
rect 4926 24998 4938 25050
rect 4990 24998 5002 25050
rect 5054 24998 5066 25050
rect 5118 24998 5130 25050
rect 5182 24998 35594 25050
rect 35646 24998 35658 25050
rect 35710 24998 35722 25050
rect 35774 24998 35786 25050
rect 35838 24998 35850 25050
rect 35902 24998 58880 25050
rect 1104 24976 58880 24998
rect 19794 24896 19800 24948
rect 19852 24896 19858 24948
rect 20898 24896 20904 24948
rect 20956 24936 20962 24948
rect 23566 24936 23572 24948
rect 20956 24908 23572 24936
rect 20956 24896 20962 24908
rect 23566 24896 23572 24908
rect 23624 24896 23630 24948
rect 26326 24936 26332 24948
rect 25056 24908 26332 24936
rect 18230 24828 18236 24880
rect 18288 24828 18294 24880
rect 19702 24828 19708 24880
rect 19760 24868 19766 24880
rect 19886 24868 19892 24880
rect 19760 24840 19892 24868
rect 19760 24828 19766 24840
rect 19886 24828 19892 24840
rect 19944 24868 19950 24880
rect 20165 24871 20223 24877
rect 20165 24868 20177 24871
rect 19944 24840 20177 24868
rect 19944 24828 19950 24840
rect 20165 24837 20177 24840
rect 20211 24837 20223 24871
rect 20165 24831 20223 24837
rect 22097 24871 22155 24877
rect 22097 24837 22109 24871
rect 22143 24868 22155 24871
rect 22370 24868 22376 24880
rect 22143 24840 22376 24868
rect 22143 24837 22155 24840
rect 22097 24831 22155 24837
rect 22370 24828 22376 24840
rect 22428 24828 22434 24880
rect 22554 24828 22560 24880
rect 22612 24828 22618 24880
rect 17954 24760 17960 24812
rect 18012 24760 18018 24812
rect 19981 24803 20039 24809
rect 19352 24596 19380 24786
rect 19981 24769 19993 24803
rect 20027 24769 20039 24803
rect 19981 24763 20039 24769
rect 19996 24732 20024 24763
rect 20070 24760 20076 24812
rect 20128 24760 20134 24812
rect 20349 24803 20407 24809
rect 20349 24769 20361 24803
rect 20395 24800 20407 24803
rect 20530 24800 20536 24812
rect 20395 24772 20536 24800
rect 20395 24769 20407 24772
rect 20349 24763 20407 24769
rect 20530 24760 20536 24772
rect 20588 24760 20594 24812
rect 24949 24803 25007 24809
rect 24949 24769 24961 24803
rect 24995 24800 25007 24803
rect 25056 24800 25084 24908
rect 26326 24896 26332 24908
rect 26384 24896 26390 24948
rect 26513 24939 26571 24945
rect 26513 24905 26525 24939
rect 26559 24936 26571 24939
rect 26559 24908 30144 24936
rect 26559 24905 26571 24908
rect 26513 24899 26571 24905
rect 25133 24871 25191 24877
rect 25133 24837 25145 24871
rect 25179 24868 25191 24871
rect 25590 24868 25596 24880
rect 25179 24840 25596 24868
rect 25179 24837 25191 24840
rect 25133 24831 25191 24837
rect 25590 24828 25596 24840
rect 25648 24828 25654 24880
rect 25682 24828 25688 24880
rect 25740 24868 25746 24880
rect 26528 24868 26556 24899
rect 25740 24840 25912 24868
rect 25740 24828 25746 24840
rect 25225 24803 25283 24809
rect 25225 24800 25237 24803
rect 24995 24772 25084 24800
rect 25148 24772 25237 24800
rect 24995 24769 25007 24772
rect 24949 24763 25007 24769
rect 21726 24732 21732 24744
rect 19996 24704 21732 24732
rect 21726 24692 21732 24704
rect 21784 24692 21790 24744
rect 21818 24692 21824 24744
rect 21876 24732 21882 24744
rect 22830 24732 22836 24744
rect 21876 24704 22836 24732
rect 21876 24692 21882 24704
rect 22830 24692 22836 24704
rect 22888 24692 22894 24744
rect 19610 24624 19616 24676
rect 19668 24664 19674 24676
rect 19705 24667 19763 24673
rect 19705 24664 19717 24667
rect 19668 24636 19717 24664
rect 19668 24624 19674 24636
rect 19705 24633 19717 24636
rect 19751 24664 19763 24667
rect 20622 24664 20628 24676
rect 19751 24636 20628 24664
rect 19751 24633 19763 24636
rect 19705 24627 19763 24633
rect 20622 24624 20628 24636
rect 20680 24624 20686 24676
rect 20806 24624 20812 24676
rect 20864 24664 20870 24676
rect 20864 24636 21680 24664
rect 20864 24624 20870 24636
rect 20438 24596 20444 24608
rect 19352 24568 20444 24596
rect 20438 24556 20444 24568
rect 20496 24596 20502 24608
rect 21545 24599 21603 24605
rect 21545 24596 21557 24599
rect 20496 24568 21557 24596
rect 20496 24556 20502 24568
rect 21545 24565 21557 24568
rect 21591 24565 21603 24599
rect 21652 24596 21680 24636
rect 23106 24624 23112 24676
rect 23164 24664 23170 24676
rect 25148 24664 25176 24772
rect 25225 24769 25237 24772
rect 25271 24769 25283 24803
rect 25225 24763 25283 24769
rect 25314 24760 25320 24812
rect 25372 24760 25378 24812
rect 25884 24809 25912 24840
rect 25976 24840 26556 24868
rect 30116 24868 30144 24908
rect 30190 24896 30196 24948
rect 30248 24936 30254 24948
rect 31846 24936 31852 24948
rect 30248 24908 31852 24936
rect 30248 24896 30254 24908
rect 31846 24896 31852 24908
rect 31904 24896 31910 24948
rect 32125 24939 32183 24945
rect 32125 24905 32137 24939
rect 32171 24905 32183 24939
rect 32125 24899 32183 24905
rect 35360 24908 38240 24936
rect 31478 24868 31484 24880
rect 30116 24840 31484 24868
rect 25976 24812 26004 24840
rect 31478 24828 31484 24840
rect 31536 24828 31542 24880
rect 32030 24868 32036 24880
rect 31588 24840 32036 24868
rect 25777 24803 25835 24809
rect 25777 24769 25789 24803
rect 25823 24769 25835 24803
rect 25777 24763 25835 24769
rect 25869 24803 25927 24809
rect 25869 24769 25881 24803
rect 25915 24769 25927 24803
rect 25869 24763 25927 24769
rect 23164 24636 25176 24664
rect 23164 24624 23170 24636
rect 25406 24624 25412 24676
rect 25464 24664 25470 24676
rect 25593 24667 25651 24673
rect 25593 24664 25605 24667
rect 25464 24636 25605 24664
rect 25464 24624 25470 24636
rect 25593 24633 25605 24636
rect 25639 24633 25651 24667
rect 25593 24627 25651 24633
rect 23290 24596 23296 24608
rect 21652 24568 23296 24596
rect 21545 24559 21603 24565
rect 23290 24556 23296 24568
rect 23348 24556 23354 24608
rect 23566 24556 23572 24608
rect 23624 24556 23630 24608
rect 24857 24599 24915 24605
rect 24857 24565 24869 24599
rect 24903 24596 24915 24599
rect 25314 24596 25320 24608
rect 24903 24568 25320 24596
rect 24903 24565 24915 24568
rect 24857 24559 24915 24565
rect 25314 24556 25320 24568
rect 25372 24556 25378 24608
rect 25498 24556 25504 24608
rect 25556 24556 25562 24608
rect 25792 24596 25820 24763
rect 25958 24760 25964 24812
rect 26016 24760 26022 24812
rect 26050 24760 26056 24812
rect 26108 24760 26114 24812
rect 26145 24803 26203 24809
rect 26145 24769 26157 24803
rect 26191 24800 26203 24803
rect 27430 24800 27436 24812
rect 26191 24772 27436 24800
rect 26191 24769 26203 24772
rect 26145 24763 26203 24769
rect 27430 24760 27436 24772
rect 27488 24760 27494 24812
rect 28902 24760 28908 24812
rect 28960 24760 28966 24812
rect 31588 24809 31616 24840
rect 32030 24828 32036 24840
rect 32088 24828 32094 24880
rect 31573 24803 31631 24809
rect 31573 24769 31585 24803
rect 31619 24769 31631 24803
rect 31573 24763 31631 24769
rect 31665 24803 31723 24809
rect 31665 24769 31677 24803
rect 31711 24769 31723 24803
rect 31665 24763 31723 24769
rect 27522 24692 27528 24744
rect 27580 24692 27586 24744
rect 27798 24692 27804 24744
rect 27856 24692 27862 24744
rect 28350 24692 28356 24744
rect 28408 24732 28414 24744
rect 29273 24735 29331 24741
rect 29273 24732 29285 24735
rect 28408 24704 29285 24732
rect 28408 24692 28414 24704
rect 29273 24701 29285 24704
rect 29319 24732 29331 24735
rect 29917 24735 29975 24741
rect 29917 24732 29929 24735
rect 29319 24704 29929 24732
rect 29319 24701 29331 24704
rect 29273 24695 29331 24701
rect 29917 24701 29929 24704
rect 29963 24701 29975 24735
rect 31680 24732 31708 24763
rect 31846 24760 31852 24812
rect 31904 24800 31910 24812
rect 31941 24803 31999 24809
rect 31941 24800 31953 24803
rect 31904 24772 31953 24800
rect 31904 24760 31910 24772
rect 31941 24769 31953 24772
rect 31987 24769 31999 24803
rect 31941 24763 31999 24769
rect 32140 24732 32168 24899
rect 32401 24871 32459 24877
rect 32401 24837 32413 24871
rect 32447 24868 32459 24871
rect 33042 24868 33048 24880
rect 32447 24840 33048 24868
rect 32447 24837 32459 24840
rect 32401 24831 32459 24837
rect 33042 24828 33048 24840
rect 33100 24828 33106 24880
rect 33134 24828 33140 24880
rect 33192 24868 33198 24880
rect 35360 24868 35388 24908
rect 33192 24840 35388 24868
rect 33192 24828 33198 24840
rect 35434 24828 35440 24880
rect 35492 24868 35498 24880
rect 38010 24877 38016 24880
rect 35989 24871 36047 24877
rect 35989 24868 36001 24871
rect 35492 24840 35664 24868
rect 35492 24828 35498 24840
rect 32309 24803 32367 24809
rect 32309 24769 32321 24803
rect 32355 24769 32367 24803
rect 32309 24763 32367 24769
rect 31680 24704 32168 24732
rect 32324 24732 32352 24763
rect 32490 24760 32496 24812
rect 32548 24760 32554 24812
rect 32674 24760 32680 24812
rect 32732 24760 32738 24812
rect 33410 24800 33416 24812
rect 32784 24772 33416 24800
rect 32582 24732 32588 24744
rect 32324 24704 32588 24732
rect 29917 24695 29975 24701
rect 32582 24692 32588 24704
rect 32640 24732 32646 24744
rect 32784 24732 32812 24772
rect 33410 24760 33416 24772
rect 33468 24760 33474 24812
rect 34974 24760 34980 24812
rect 35032 24760 35038 24812
rect 35066 24760 35072 24812
rect 35124 24800 35130 24812
rect 35636 24809 35664 24840
rect 35820 24840 36001 24868
rect 35345 24803 35403 24809
rect 35345 24800 35357 24803
rect 35124 24772 35357 24800
rect 35124 24760 35130 24772
rect 35345 24769 35357 24772
rect 35391 24769 35403 24803
rect 35345 24763 35403 24769
rect 35529 24803 35587 24809
rect 35529 24769 35541 24803
rect 35575 24769 35587 24803
rect 35529 24763 35587 24769
rect 35621 24803 35679 24809
rect 35621 24769 35633 24803
rect 35667 24769 35679 24803
rect 35621 24763 35679 24769
rect 32640 24704 32812 24732
rect 32640 24692 32646 24704
rect 33226 24692 33232 24744
rect 33284 24732 33290 24744
rect 34422 24732 34428 24744
rect 33284 24704 34428 24732
rect 33284 24692 33290 24704
rect 34422 24692 34428 24704
rect 34480 24732 34486 24744
rect 35544 24732 35572 24763
rect 35710 24760 35716 24812
rect 35768 24800 35774 24812
rect 35820 24800 35848 24840
rect 35989 24837 36001 24840
rect 36035 24837 36047 24871
rect 35989 24831 36047 24837
rect 37997 24871 38016 24877
rect 37997 24837 38009 24871
rect 37997 24831 38016 24837
rect 38010 24828 38016 24831
rect 38068 24828 38074 24880
rect 38212 24877 38240 24908
rect 42426 24896 42432 24948
rect 42484 24936 42490 24948
rect 42702 24936 42708 24948
rect 42484 24908 42708 24936
rect 42484 24896 42490 24908
rect 42702 24896 42708 24908
rect 42760 24896 42766 24948
rect 45830 24896 45836 24948
rect 45888 24896 45894 24948
rect 45922 24896 45928 24948
rect 45980 24896 45986 24948
rect 47394 24896 47400 24948
rect 47452 24936 47458 24948
rect 49418 24936 49424 24948
rect 47452 24908 49424 24936
rect 47452 24896 47458 24908
rect 49418 24896 49424 24908
rect 49476 24896 49482 24948
rect 49970 24896 49976 24948
rect 50028 24936 50034 24948
rect 50065 24939 50123 24945
rect 50065 24936 50077 24939
rect 50028 24908 50077 24936
rect 50028 24896 50034 24908
rect 50065 24905 50077 24908
rect 50111 24905 50123 24939
rect 50065 24899 50123 24905
rect 50433 24939 50491 24945
rect 50433 24905 50445 24939
rect 50479 24936 50491 24939
rect 50522 24936 50528 24948
rect 50479 24908 50528 24936
rect 50479 24905 50491 24908
rect 50433 24899 50491 24905
rect 50522 24896 50528 24908
rect 50580 24896 50586 24948
rect 51994 24896 52000 24948
rect 52052 24936 52058 24948
rect 54110 24936 54116 24948
rect 52052 24908 54116 24936
rect 52052 24896 52058 24908
rect 54110 24896 54116 24908
rect 54168 24896 54174 24948
rect 55306 24896 55312 24948
rect 55364 24896 55370 24948
rect 38197 24871 38255 24877
rect 38197 24837 38209 24871
rect 38243 24837 38255 24871
rect 38197 24831 38255 24837
rect 39761 24871 39819 24877
rect 39761 24837 39773 24871
rect 39807 24868 39819 24871
rect 40034 24868 40040 24880
rect 39807 24840 40040 24868
rect 39807 24837 39819 24840
rect 39761 24831 39819 24837
rect 40034 24828 40040 24840
rect 40092 24868 40098 24880
rect 43257 24871 43315 24877
rect 43257 24868 43269 24871
rect 40092 24840 41092 24868
rect 40092 24828 40098 24840
rect 35768 24772 35848 24800
rect 35897 24803 35955 24809
rect 35768 24760 35774 24772
rect 35897 24769 35909 24803
rect 35943 24800 35955 24803
rect 36262 24800 36268 24812
rect 35943 24772 36268 24800
rect 35943 24769 35955 24772
rect 35897 24763 35955 24769
rect 36262 24760 36268 24772
rect 36320 24760 36326 24812
rect 37461 24803 37519 24809
rect 37461 24769 37473 24803
rect 37507 24800 37519 24803
rect 37550 24800 37556 24812
rect 37507 24772 37556 24800
rect 37507 24769 37519 24772
rect 37461 24763 37519 24769
rect 37550 24760 37556 24772
rect 37608 24760 37614 24812
rect 37737 24803 37795 24809
rect 37737 24769 37749 24803
rect 37783 24800 37795 24803
rect 38470 24800 38476 24812
rect 37783 24772 38476 24800
rect 37783 24769 37795 24772
rect 37737 24763 37795 24769
rect 38470 24760 38476 24772
rect 38528 24760 38534 24812
rect 39853 24803 39911 24809
rect 39853 24769 39865 24803
rect 39899 24800 39911 24803
rect 39942 24800 39948 24812
rect 39899 24772 39948 24800
rect 39899 24769 39911 24772
rect 39853 24763 39911 24769
rect 39942 24760 39948 24772
rect 40000 24760 40006 24812
rect 40865 24803 40923 24809
rect 40865 24769 40877 24803
rect 40911 24769 40923 24803
rect 40865 24763 40923 24769
rect 34480 24704 35572 24732
rect 35805 24735 35863 24741
rect 34480 24692 34486 24704
rect 35805 24701 35817 24735
rect 35851 24732 35863 24735
rect 36078 24732 36084 24744
rect 35851 24704 36084 24732
rect 35851 24701 35863 24704
rect 35805 24695 35863 24701
rect 36078 24692 36084 24704
rect 36136 24692 36142 24744
rect 37645 24735 37703 24741
rect 37645 24701 37657 24735
rect 37691 24701 37703 24735
rect 37645 24695 37703 24701
rect 25958 24624 25964 24676
rect 26016 24664 26022 24676
rect 26016 24636 26464 24664
rect 26016 24624 26022 24636
rect 26326 24596 26332 24608
rect 25792 24568 26332 24596
rect 26326 24556 26332 24568
rect 26384 24556 26390 24608
rect 26436 24596 26464 24636
rect 32306 24624 32312 24676
rect 32364 24664 32370 24676
rect 37660 24664 37688 24695
rect 37829 24667 37887 24673
rect 37829 24664 37841 24667
rect 32364 24636 37596 24664
rect 37660 24636 37841 24664
rect 32364 24624 32370 24636
rect 28994 24596 29000 24608
rect 26436 24568 29000 24596
rect 28994 24556 29000 24568
rect 29052 24556 29058 24608
rect 29362 24556 29368 24608
rect 29420 24556 29426 24608
rect 31386 24556 31392 24608
rect 31444 24556 31450 24608
rect 31754 24556 31760 24608
rect 31812 24596 31818 24608
rect 31849 24599 31907 24605
rect 31849 24596 31861 24599
rect 31812 24568 31861 24596
rect 31812 24556 31818 24568
rect 31849 24565 31861 24568
rect 31895 24596 31907 24599
rect 32766 24596 32772 24608
rect 31895 24568 32772 24596
rect 31895 24565 31907 24568
rect 31849 24559 31907 24565
rect 32766 24556 32772 24568
rect 32824 24556 32830 24608
rect 34514 24556 34520 24608
rect 34572 24596 34578 24608
rect 37277 24599 37335 24605
rect 37277 24596 37289 24599
rect 34572 24568 37289 24596
rect 34572 24556 34578 24568
rect 37277 24565 37289 24568
rect 37323 24565 37335 24599
rect 37277 24559 37335 24565
rect 37458 24556 37464 24608
rect 37516 24556 37522 24608
rect 37568 24596 37596 24636
rect 37829 24633 37841 24636
rect 37875 24633 37887 24667
rect 38746 24664 38752 24676
rect 37829 24627 37887 24633
rect 37936 24636 38752 24664
rect 37936 24596 37964 24636
rect 38746 24624 38752 24636
rect 38804 24624 38810 24676
rect 39850 24624 39856 24676
rect 39908 24664 39914 24676
rect 40589 24667 40647 24673
rect 40589 24664 40601 24667
rect 39908 24636 40601 24664
rect 39908 24624 39914 24636
rect 40589 24633 40601 24636
rect 40635 24633 40647 24667
rect 40880 24664 40908 24763
rect 40954 24760 40960 24812
rect 41012 24760 41018 24812
rect 41064 24809 41092 24840
rect 41616 24840 43269 24868
rect 41049 24803 41107 24809
rect 41049 24769 41061 24803
rect 41095 24769 41107 24803
rect 41049 24763 41107 24769
rect 41233 24803 41291 24809
rect 41233 24769 41245 24803
rect 41279 24800 41291 24803
rect 41414 24800 41420 24812
rect 41279 24772 41420 24800
rect 41279 24769 41291 24772
rect 41233 24763 41291 24769
rect 41414 24760 41420 24772
rect 41472 24800 41478 24812
rect 41616 24809 41644 24840
rect 43257 24837 43269 24840
rect 43303 24837 43315 24871
rect 45848 24868 45876 24896
rect 45848 24840 46336 24868
rect 43257 24831 43315 24837
rect 41601 24803 41659 24809
rect 41601 24800 41613 24803
rect 41472 24772 41613 24800
rect 41472 24760 41478 24772
rect 41601 24769 41613 24772
rect 41647 24769 41659 24803
rect 41601 24763 41659 24769
rect 41782 24760 41788 24812
rect 41840 24760 41846 24812
rect 41877 24803 41935 24809
rect 41877 24769 41889 24803
rect 41923 24769 41935 24803
rect 41877 24763 41935 24769
rect 41969 24803 42027 24809
rect 41969 24769 41981 24803
rect 42015 24800 42027 24803
rect 42150 24800 42156 24812
rect 42015 24772 42156 24800
rect 42015 24769 42027 24772
rect 41969 24763 42027 24769
rect 40972 24732 41000 24760
rect 41322 24732 41328 24744
rect 40972 24704 41328 24732
rect 41322 24692 41328 24704
rect 41380 24732 41386 24744
rect 41892 24732 41920 24763
rect 41380 24704 41920 24732
rect 41380 24692 41386 24704
rect 41984 24664 42012 24763
rect 42150 24760 42156 24772
rect 42208 24760 42214 24812
rect 42613 24803 42671 24809
rect 42613 24769 42625 24803
rect 42659 24769 42671 24803
rect 42613 24763 42671 24769
rect 42628 24732 42656 24763
rect 42702 24760 42708 24812
rect 42760 24760 42766 24812
rect 46106 24760 46112 24812
rect 46164 24760 46170 24812
rect 46308 24809 46336 24840
rect 48774 24828 48780 24880
rect 48832 24828 48838 24880
rect 48958 24828 48964 24880
rect 49016 24868 49022 24880
rect 49789 24871 49847 24877
rect 49789 24868 49801 24871
rect 49016 24840 49801 24868
rect 49016 24828 49022 24840
rect 49789 24837 49801 24840
rect 49835 24868 49847 24871
rect 50154 24868 50160 24880
rect 49835 24840 50160 24868
rect 49835 24837 49847 24840
rect 49789 24831 49847 24837
rect 50154 24828 50160 24840
rect 50212 24828 50218 24880
rect 50706 24868 50712 24880
rect 50540 24840 50712 24868
rect 46293 24803 46351 24809
rect 46293 24769 46305 24803
rect 46339 24769 46351 24803
rect 46293 24763 46351 24769
rect 46385 24803 46443 24809
rect 46385 24769 46397 24803
rect 46431 24800 46443 24803
rect 46474 24800 46480 24812
rect 46431 24772 46480 24800
rect 46431 24769 46443 24772
rect 46385 24763 46443 24769
rect 46474 24760 46480 24772
rect 46532 24760 46538 24812
rect 46569 24803 46627 24809
rect 46569 24769 46581 24803
rect 46615 24800 46627 24803
rect 49605 24803 49663 24809
rect 49605 24800 49617 24803
rect 46615 24772 47808 24800
rect 46615 24769 46627 24772
rect 46569 24763 46627 24769
rect 42886 24732 42892 24744
rect 40880 24636 42012 24664
rect 42076 24704 42892 24732
rect 40589 24627 40647 24633
rect 37568 24568 37964 24596
rect 38013 24599 38071 24605
rect 38013 24565 38025 24599
rect 38059 24596 38071 24599
rect 38286 24596 38292 24608
rect 38059 24568 38292 24596
rect 38059 24565 38071 24568
rect 38013 24559 38071 24565
rect 38286 24556 38292 24568
rect 38344 24556 38350 24608
rect 39574 24556 39580 24608
rect 39632 24556 39638 24608
rect 39666 24556 39672 24608
rect 39724 24596 39730 24608
rect 40037 24599 40095 24605
rect 40037 24596 40049 24599
rect 39724 24568 40049 24596
rect 39724 24556 39730 24568
rect 40037 24565 40049 24568
rect 40083 24596 40095 24599
rect 40126 24596 40132 24608
rect 40083 24568 40132 24596
rect 40083 24565 40095 24568
rect 40037 24559 40095 24565
rect 40126 24556 40132 24568
rect 40184 24596 40190 24608
rect 40494 24596 40500 24608
rect 40184 24568 40500 24596
rect 40184 24556 40190 24568
rect 40494 24556 40500 24568
rect 40552 24556 40558 24608
rect 41782 24556 41788 24608
rect 41840 24596 41846 24608
rect 42076 24596 42104 24704
rect 42886 24692 42892 24704
rect 42944 24692 42950 24744
rect 42978 24692 42984 24744
rect 43036 24732 43042 24744
rect 43806 24732 43812 24744
rect 43036 24704 43812 24732
rect 43036 24692 43042 24704
rect 43806 24692 43812 24704
rect 43864 24692 43870 24744
rect 42245 24667 42303 24673
rect 42245 24633 42257 24667
rect 42291 24664 42303 24667
rect 42794 24664 42800 24676
rect 42291 24636 42800 24664
rect 42291 24633 42303 24636
rect 42245 24627 42303 24633
rect 42794 24624 42800 24636
rect 42852 24624 42858 24676
rect 42904 24664 42932 24692
rect 43533 24667 43591 24673
rect 43533 24664 43545 24667
rect 42904 24636 43545 24664
rect 43533 24633 43545 24636
rect 43579 24664 43591 24667
rect 43622 24664 43628 24676
rect 43579 24636 43628 24664
rect 43579 24633 43591 24636
rect 43533 24627 43591 24633
rect 43622 24624 43628 24636
rect 43680 24624 43686 24676
rect 47581 24667 47639 24673
rect 47581 24664 47593 24667
rect 46400 24636 47593 24664
rect 46400 24608 46428 24636
rect 47581 24633 47593 24636
rect 47627 24633 47639 24667
rect 47581 24627 47639 24633
rect 41840 24568 42104 24596
rect 41840 24556 41846 24568
rect 42426 24556 42432 24608
rect 42484 24556 42490 24608
rect 42889 24599 42947 24605
rect 42889 24565 42901 24599
rect 42935 24596 42947 24599
rect 42978 24596 42984 24608
rect 42935 24568 42984 24596
rect 42935 24565 42947 24568
rect 42889 24559 42947 24565
rect 42978 24556 42984 24568
rect 43036 24556 43042 24608
rect 43714 24556 43720 24608
rect 43772 24556 43778 24608
rect 46382 24556 46388 24608
rect 46440 24556 46446 24608
rect 46845 24599 46903 24605
rect 46845 24565 46857 24599
rect 46891 24596 46903 24599
rect 47026 24596 47032 24608
rect 46891 24568 47032 24596
rect 46891 24565 46903 24568
rect 46845 24559 46903 24565
rect 47026 24556 47032 24568
rect 47084 24556 47090 24608
rect 47121 24599 47179 24605
rect 47121 24565 47133 24599
rect 47167 24596 47179 24599
rect 47210 24596 47216 24608
rect 47167 24568 47216 24596
rect 47167 24565 47179 24568
rect 47121 24559 47179 24565
rect 47210 24556 47216 24568
rect 47268 24556 47274 24608
rect 47305 24599 47363 24605
rect 47305 24565 47317 24599
rect 47351 24596 47363 24599
rect 47780 24596 47808 24772
rect 49252 24772 49617 24800
rect 49252 24744 49280 24772
rect 49605 24769 49617 24772
rect 49651 24769 49663 24803
rect 49605 24763 49663 24769
rect 49697 24803 49755 24809
rect 49697 24769 49709 24803
rect 49743 24769 49755 24803
rect 49697 24763 49755 24769
rect 49234 24692 49240 24744
rect 49292 24692 49298 24744
rect 49712 24732 49740 24763
rect 49970 24760 49976 24812
rect 50028 24760 50034 24812
rect 50246 24760 50252 24812
rect 50304 24760 50310 24812
rect 50540 24809 50568 24840
rect 50706 24828 50712 24840
rect 50764 24828 50770 24880
rect 55324 24868 55352 24896
rect 55585 24871 55643 24877
rect 55585 24868 55597 24871
rect 55324 24840 55597 24868
rect 55585 24837 55597 24840
rect 55631 24837 55643 24871
rect 56226 24868 56232 24880
rect 55585 24831 55643 24837
rect 55968 24840 56232 24868
rect 50525 24803 50583 24809
rect 50525 24769 50537 24803
rect 50571 24769 50583 24803
rect 50525 24763 50583 24769
rect 50614 24760 50620 24812
rect 50672 24800 50678 24812
rect 51350 24800 51356 24812
rect 50672 24772 51356 24800
rect 50672 24760 50678 24772
rect 51350 24760 51356 24772
rect 51408 24760 51414 24812
rect 52822 24760 52828 24812
rect 52880 24760 52886 24812
rect 53466 24760 53472 24812
rect 53524 24800 53530 24812
rect 55398 24809 55404 24812
rect 55217 24803 55275 24809
rect 55217 24800 55229 24803
rect 53524 24772 55229 24800
rect 53524 24760 53530 24772
rect 55217 24769 55229 24772
rect 55263 24769 55275 24803
rect 55217 24763 55275 24769
rect 55365 24803 55404 24809
rect 55365 24769 55377 24803
rect 55365 24763 55404 24769
rect 55398 24760 55404 24763
rect 55456 24760 55462 24812
rect 55493 24803 55551 24809
rect 55493 24769 55505 24803
rect 55539 24769 55551 24803
rect 55493 24763 55551 24769
rect 51626 24732 51632 24744
rect 49712 24704 51632 24732
rect 51626 24692 51632 24704
rect 51684 24732 51690 24744
rect 53374 24732 53380 24744
rect 51684 24704 53380 24732
rect 51684 24692 51690 24704
rect 53374 24692 53380 24704
rect 53432 24692 53438 24744
rect 49602 24664 49608 24676
rect 48700 24636 49608 24664
rect 48700 24596 48728 24636
rect 49602 24624 49608 24636
rect 49660 24624 49666 24676
rect 50890 24624 50896 24676
rect 50948 24664 50954 24676
rect 55306 24664 55312 24676
rect 50948 24636 55312 24664
rect 50948 24624 50954 24636
rect 55306 24624 55312 24636
rect 55364 24624 55370 24676
rect 47351 24568 48728 24596
rect 47351 24565 47363 24568
rect 47305 24559 47363 24565
rect 48958 24556 48964 24608
rect 49016 24596 49022 24608
rect 49053 24599 49111 24605
rect 49053 24596 49065 24599
rect 49016 24568 49065 24596
rect 49016 24556 49022 24568
rect 49053 24565 49065 24568
rect 49099 24565 49111 24599
rect 49053 24559 49111 24565
rect 49418 24556 49424 24608
rect 49476 24556 49482 24608
rect 54202 24556 54208 24608
rect 54260 24596 54266 24608
rect 55508 24596 55536 24763
rect 55674 24760 55680 24812
rect 55732 24809 55738 24812
rect 55732 24800 55740 24809
rect 55732 24772 55777 24800
rect 55732 24763 55740 24772
rect 55732 24760 55738 24763
rect 55968 24741 55996 24840
rect 56226 24828 56232 24840
rect 56284 24828 56290 24880
rect 56502 24828 56508 24880
rect 56560 24868 56566 24880
rect 56560 24840 56718 24868
rect 56560 24828 56566 24840
rect 55953 24735 56011 24741
rect 55953 24732 55965 24735
rect 55600 24704 55965 24732
rect 55600 24676 55628 24704
rect 55953 24701 55965 24704
rect 55999 24701 56011 24735
rect 55953 24695 56011 24701
rect 56226 24692 56232 24744
rect 56284 24692 56290 24744
rect 55582 24624 55588 24676
rect 55640 24624 55646 24676
rect 54260 24568 55536 24596
rect 55861 24599 55919 24605
rect 54260 24556 54266 24568
rect 55861 24565 55873 24599
rect 55907 24596 55919 24599
rect 56318 24596 56324 24608
rect 55907 24568 56324 24596
rect 55907 24565 55919 24568
rect 55861 24559 55919 24565
rect 56318 24556 56324 24568
rect 56376 24556 56382 24608
rect 57698 24556 57704 24608
rect 57756 24556 57762 24608
rect 1104 24506 58880 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 58880 24506
rect 1104 24432 58880 24454
rect 20438 24352 20444 24404
rect 20496 24392 20502 24404
rect 22554 24392 22560 24404
rect 20496 24364 22560 24392
rect 20496 24352 20502 24364
rect 22554 24352 22560 24364
rect 22612 24352 22618 24404
rect 22833 24395 22891 24401
rect 22833 24361 22845 24395
rect 22879 24392 22891 24395
rect 22922 24392 22928 24404
rect 22879 24364 22928 24392
rect 22879 24361 22891 24364
rect 22833 24355 22891 24361
rect 22922 24352 22928 24364
rect 22980 24352 22986 24404
rect 23106 24352 23112 24404
rect 23164 24352 23170 24404
rect 24949 24395 25007 24401
rect 24949 24361 24961 24395
rect 24995 24392 25007 24395
rect 25130 24392 25136 24404
rect 24995 24364 25136 24392
rect 24995 24361 25007 24364
rect 24949 24355 25007 24361
rect 25130 24352 25136 24364
rect 25188 24352 25194 24404
rect 25409 24395 25467 24401
rect 25409 24361 25421 24395
rect 25455 24392 25467 24395
rect 26145 24395 26203 24401
rect 26145 24392 26157 24395
rect 25455 24364 26157 24392
rect 25455 24361 25467 24364
rect 25409 24355 25467 24361
rect 26145 24361 26157 24364
rect 26191 24361 26203 24395
rect 26145 24355 26203 24361
rect 26510 24352 26516 24404
rect 26568 24352 26574 24404
rect 27798 24352 27804 24404
rect 27856 24392 27862 24404
rect 27985 24395 28043 24401
rect 27985 24392 27997 24395
rect 27856 24364 27997 24392
rect 27856 24352 27862 24364
rect 27985 24361 27997 24364
rect 28031 24361 28043 24395
rect 27985 24355 28043 24361
rect 28445 24395 28503 24401
rect 28445 24361 28457 24395
rect 28491 24392 28503 24395
rect 31754 24392 31760 24404
rect 28491 24364 31760 24392
rect 28491 24361 28503 24364
rect 28445 24355 28503 24361
rect 31754 24352 31760 24364
rect 31812 24352 31818 24404
rect 31846 24352 31852 24404
rect 31904 24392 31910 24404
rect 32122 24392 32128 24404
rect 31904 24364 32128 24392
rect 31904 24352 31910 24364
rect 32122 24352 32128 24364
rect 32180 24392 32186 24404
rect 32582 24392 32588 24404
rect 32180 24364 32588 24392
rect 32180 24352 32186 24364
rect 32582 24352 32588 24364
rect 32640 24392 32646 24404
rect 32815 24395 32873 24401
rect 32815 24392 32827 24395
rect 32640 24364 32827 24392
rect 32640 24352 32646 24364
rect 32815 24361 32827 24364
rect 32861 24392 32873 24395
rect 33134 24392 33140 24404
rect 32861 24364 33140 24392
rect 32861 24361 32873 24364
rect 32815 24355 32873 24361
rect 33134 24352 33140 24364
rect 33192 24352 33198 24404
rect 34054 24352 34060 24404
rect 34112 24352 34118 24404
rect 34514 24352 34520 24404
rect 34572 24352 34578 24404
rect 35986 24352 35992 24404
rect 36044 24352 36050 24404
rect 36078 24352 36084 24404
rect 36136 24392 36142 24404
rect 36136 24364 36400 24392
rect 36136 24352 36142 24364
rect 21818 24284 21824 24336
rect 21876 24324 21882 24336
rect 21876 24296 23060 24324
rect 21876 24284 21882 24296
rect 19705 24259 19763 24265
rect 19705 24225 19717 24259
rect 19751 24256 19763 24259
rect 21542 24256 21548 24268
rect 19751 24228 21548 24256
rect 19751 24225 19763 24228
rect 19705 24219 19763 24225
rect 21542 24216 21548 24228
rect 21600 24216 21606 24268
rect 22554 24216 22560 24268
rect 22612 24256 22618 24268
rect 22612 24228 22784 24256
rect 22612 24216 22618 24228
rect 19429 24191 19487 24197
rect 19429 24157 19441 24191
rect 19475 24157 19487 24191
rect 19429 24151 19487 24157
rect 18506 24012 18512 24064
rect 18564 24052 18570 24064
rect 19245 24055 19303 24061
rect 19245 24052 19257 24055
rect 18564 24024 19257 24052
rect 18564 24012 18570 24024
rect 19245 24021 19257 24024
rect 19291 24021 19303 24055
rect 19444 24052 19472 24151
rect 19518 24148 19524 24200
rect 19576 24148 19582 24200
rect 19797 24191 19855 24197
rect 19797 24157 19809 24191
rect 19843 24188 19855 24191
rect 19978 24188 19984 24200
rect 19843 24160 19984 24188
rect 19843 24157 19855 24160
rect 19797 24151 19855 24157
rect 19978 24148 19984 24160
rect 20036 24148 20042 24200
rect 22278 24148 22284 24200
rect 22336 24188 22342 24200
rect 22373 24191 22431 24197
rect 22373 24188 22385 24191
rect 22336 24160 22385 24188
rect 22336 24148 22342 24160
rect 22373 24157 22385 24160
rect 22419 24157 22431 24191
rect 22373 24151 22431 24157
rect 22462 24148 22468 24200
rect 22520 24148 22526 24200
rect 22756 24197 22784 24228
rect 23032 24197 23060 24296
rect 23124 24197 23152 24352
rect 23290 24284 23296 24336
rect 23348 24284 23354 24336
rect 25314 24284 25320 24336
rect 25372 24324 25378 24336
rect 26050 24324 26056 24336
rect 25372 24296 26056 24324
rect 25372 24284 25378 24296
rect 26050 24284 26056 24296
rect 26108 24324 26114 24336
rect 26108 24296 26832 24324
rect 26108 24284 26114 24296
rect 23566 24216 23572 24268
rect 23624 24256 23630 24268
rect 26418 24256 26424 24268
rect 23624 24228 26424 24256
rect 23624 24216 23630 24228
rect 26418 24216 26424 24228
rect 26476 24216 26482 24268
rect 22741 24191 22799 24197
rect 22741 24157 22753 24191
rect 22787 24157 22799 24191
rect 22741 24151 22799 24157
rect 23017 24191 23075 24197
rect 23017 24157 23029 24191
rect 23063 24157 23075 24191
rect 23017 24151 23075 24157
rect 23109 24191 23167 24197
rect 23109 24157 23121 24191
rect 23155 24157 23167 24191
rect 23109 24151 23167 24157
rect 23367 24191 23425 24197
rect 23367 24157 23379 24191
rect 23413 24188 23425 24191
rect 23658 24188 23664 24200
rect 23413 24182 23428 24188
rect 23487 24182 23664 24188
rect 23413 24160 23664 24182
rect 23413 24157 23515 24160
rect 23367 24154 23515 24157
rect 23367 24151 23425 24154
rect 23658 24148 23664 24160
rect 23716 24148 23722 24200
rect 25038 24148 25044 24200
rect 25096 24188 25102 24200
rect 25133 24191 25191 24197
rect 25133 24188 25145 24191
rect 25096 24160 25145 24188
rect 25096 24148 25102 24160
rect 25133 24157 25145 24160
rect 25179 24157 25191 24191
rect 25133 24151 25191 24157
rect 25222 24148 25228 24200
rect 25280 24148 25286 24200
rect 25406 24148 25412 24200
rect 25464 24148 25470 24200
rect 25498 24148 25504 24200
rect 25556 24148 25562 24200
rect 25594 24191 25652 24197
rect 25594 24157 25606 24191
rect 25640 24157 25652 24191
rect 25594 24151 25652 24157
rect 22094 24080 22100 24132
rect 22152 24120 22158 24132
rect 22557 24123 22615 24129
rect 22557 24120 22569 24123
rect 22152 24092 22569 24120
rect 22152 24080 22158 24092
rect 22557 24089 22569 24092
rect 22603 24089 22615 24123
rect 22557 24083 22615 24089
rect 22922 24080 22928 24132
rect 22980 24120 22986 24132
rect 25608 24120 25636 24151
rect 25774 24148 25780 24200
rect 25832 24148 25838 24200
rect 26007 24191 26065 24197
rect 26007 24157 26019 24191
rect 26053 24188 26065 24191
rect 26053 24160 26740 24188
rect 26053 24157 26065 24160
rect 26007 24151 26065 24157
rect 22980 24092 25636 24120
rect 22980 24080 22986 24092
rect 25866 24080 25872 24132
rect 25924 24080 25930 24132
rect 26326 24080 26332 24132
rect 26384 24080 26390 24132
rect 20254 24052 20260 24064
rect 19444 24024 20260 24052
rect 19245 24015 19303 24021
rect 20254 24012 20260 24024
rect 20312 24052 20318 24064
rect 21818 24052 21824 24064
rect 20312 24024 21824 24052
rect 20312 24012 20318 24024
rect 21818 24012 21824 24024
rect 21876 24012 21882 24064
rect 22186 24012 22192 24064
rect 22244 24012 22250 24064
rect 24946 24012 24952 24064
rect 25004 24052 25010 24064
rect 25590 24052 25596 24064
rect 25004 24024 25596 24052
rect 25004 24012 25010 24024
rect 25590 24012 25596 24024
rect 25648 24012 25654 24064
rect 25682 24012 25688 24064
rect 25740 24052 25746 24064
rect 26344 24052 26372 24080
rect 26712 24061 26740 24160
rect 26804 24120 26832 24296
rect 27430 24284 27436 24336
rect 27488 24324 27494 24336
rect 29917 24327 29975 24333
rect 29917 24324 29929 24327
rect 27488 24296 29929 24324
rect 27488 24284 27494 24296
rect 29917 24293 29929 24296
rect 29963 24293 29975 24327
rect 29917 24287 29975 24293
rect 33781 24327 33839 24333
rect 33781 24293 33793 24327
rect 33827 24324 33839 24327
rect 34974 24324 34980 24336
rect 33827 24296 34376 24324
rect 33827 24293 33839 24296
rect 33781 24287 33839 24293
rect 28074 24216 28080 24268
rect 28132 24256 28138 24268
rect 28350 24256 28356 24268
rect 28132 24228 28356 24256
rect 28132 24216 28138 24228
rect 28350 24216 28356 24228
rect 28408 24216 28414 24268
rect 29362 24256 29368 24268
rect 28644 24228 29368 24256
rect 26970 24148 26976 24200
rect 27028 24188 27034 24200
rect 28166 24188 28172 24200
rect 27028 24160 28172 24188
rect 27028 24148 27034 24160
rect 28166 24148 28172 24160
rect 28224 24148 28230 24200
rect 28261 24191 28319 24197
rect 28261 24157 28273 24191
rect 28307 24157 28319 24191
rect 28261 24151 28319 24157
rect 28537 24191 28595 24197
rect 28537 24157 28549 24191
rect 28583 24190 28595 24191
rect 28644 24190 28672 24228
rect 29362 24216 29368 24228
rect 29420 24216 29426 24268
rect 30024 24228 30236 24256
rect 28583 24162 28672 24190
rect 28583 24157 28595 24162
rect 28537 24151 28595 24157
rect 28276 24120 28304 24151
rect 28810 24148 28816 24200
rect 28868 24148 28874 24200
rect 28997 24191 29055 24197
rect 28997 24157 29009 24191
rect 29043 24188 29055 24191
rect 29086 24188 29092 24200
rect 29043 24160 29092 24188
rect 29043 24157 29055 24160
rect 28997 24151 29055 24157
rect 29086 24148 29092 24160
rect 29144 24188 29150 24200
rect 30024 24188 30052 24228
rect 30208 24197 30236 24228
rect 31386 24216 31392 24268
rect 31444 24216 31450 24268
rect 33042 24216 33048 24268
rect 33100 24256 33106 24268
rect 34348 24265 34376 24296
rect 34440 24296 34980 24324
rect 34333 24259 34391 24265
rect 33100 24228 33548 24256
rect 33100 24216 33106 24228
rect 29144 24160 30052 24188
rect 30096 24191 30154 24197
rect 29144 24148 29150 24160
rect 30096 24157 30108 24191
rect 30142 24157 30154 24191
rect 30096 24151 30154 24157
rect 30193 24191 30251 24197
rect 30193 24157 30205 24191
rect 30239 24157 30251 24191
rect 30193 24151 30251 24157
rect 28629 24123 28687 24129
rect 28629 24120 28641 24123
rect 26804 24092 28028 24120
rect 28276 24092 28641 24120
rect 25740 24024 26372 24052
rect 26697 24055 26755 24061
rect 25740 24012 25746 24024
rect 26697 24021 26709 24055
rect 26743 24052 26755 24055
rect 27890 24052 27896 24064
rect 26743 24024 27896 24052
rect 26743 24021 26755 24024
rect 26697 24015 26755 24021
rect 27890 24012 27896 24024
rect 27948 24012 27954 24064
rect 28000 24052 28028 24092
rect 28629 24089 28641 24092
rect 28675 24089 28687 24123
rect 28629 24083 28687 24089
rect 30006 24052 30012 24064
rect 28000 24024 30012 24052
rect 30006 24012 30012 24024
rect 30064 24012 30070 24064
rect 30111 24052 30139 24151
rect 30374 24148 30380 24200
rect 30432 24197 30438 24200
rect 30432 24191 30471 24197
rect 30459 24157 30471 24191
rect 30432 24151 30471 24157
rect 30561 24191 30619 24197
rect 30561 24157 30573 24191
rect 30607 24188 30619 24191
rect 30926 24188 30932 24200
rect 30607 24160 30932 24188
rect 30607 24157 30619 24160
rect 30561 24151 30619 24157
rect 30432 24148 30438 24151
rect 30926 24148 30932 24160
rect 30984 24148 30990 24200
rect 31018 24148 31024 24200
rect 31076 24148 31082 24200
rect 33134 24148 33140 24200
rect 33192 24148 33198 24200
rect 33520 24197 33548 24228
rect 34333 24225 34345 24259
rect 34379 24225 34391 24259
rect 34333 24219 34391 24225
rect 33230 24191 33288 24197
rect 33230 24157 33242 24191
rect 33276 24157 33288 24191
rect 33230 24151 33288 24157
rect 33505 24191 33563 24197
rect 33505 24157 33517 24191
rect 33551 24157 33563 24191
rect 33505 24151 33563 24157
rect 33643 24191 33701 24197
rect 33643 24157 33655 24191
rect 33689 24188 33701 24191
rect 33962 24188 33968 24200
rect 33689 24160 33968 24188
rect 33689 24157 33701 24160
rect 33643 24151 33701 24157
rect 30285 24123 30343 24129
rect 30285 24089 30297 24123
rect 30331 24120 30343 24123
rect 30331 24092 30880 24120
rect 30331 24089 30343 24092
rect 30285 24083 30343 24089
rect 30852 24064 30880 24092
rect 32214 24080 32220 24132
rect 32272 24080 32278 24132
rect 32674 24080 32680 24132
rect 32732 24120 32738 24132
rect 33042 24120 33048 24132
rect 32732 24092 33048 24120
rect 32732 24080 32738 24092
rect 33042 24080 33048 24092
rect 33100 24120 33106 24132
rect 33244 24120 33272 24151
rect 33962 24148 33968 24160
rect 34020 24148 34026 24200
rect 34241 24191 34299 24197
rect 34241 24157 34253 24191
rect 34287 24188 34299 24191
rect 34440 24188 34468 24296
rect 34974 24284 34980 24296
rect 35032 24284 35038 24336
rect 35250 24284 35256 24336
rect 35308 24324 35314 24336
rect 36004 24324 36032 24352
rect 36372 24336 36400 24364
rect 39942 24352 39948 24404
rect 40000 24392 40006 24404
rect 42702 24392 42708 24404
rect 40000 24364 42708 24392
rect 40000 24352 40006 24364
rect 42702 24352 42708 24364
rect 42760 24352 42766 24404
rect 43533 24395 43591 24401
rect 43533 24361 43545 24395
rect 43579 24392 43591 24395
rect 44177 24395 44235 24401
rect 44177 24392 44189 24395
rect 43579 24364 44189 24392
rect 43579 24361 43591 24364
rect 43533 24355 43591 24361
rect 44177 24361 44189 24364
rect 44223 24392 44235 24395
rect 47394 24392 47400 24404
rect 44223 24364 47400 24392
rect 44223 24361 44235 24364
rect 44177 24355 44235 24361
rect 47394 24352 47400 24364
rect 47452 24352 47458 24404
rect 48682 24392 48688 24404
rect 47504 24364 48688 24392
rect 35308 24296 36032 24324
rect 35308 24284 35314 24296
rect 34790 24216 34796 24268
rect 34848 24256 34854 24268
rect 35069 24259 35127 24265
rect 35069 24256 35081 24259
rect 34848 24228 35081 24256
rect 34848 24216 34854 24228
rect 35069 24225 35081 24228
rect 35115 24256 35127 24259
rect 35342 24256 35348 24268
rect 35115 24228 35348 24256
rect 35115 24225 35127 24228
rect 35069 24219 35127 24225
rect 35342 24216 35348 24228
rect 35400 24216 35406 24268
rect 35894 24216 35900 24268
rect 35952 24216 35958 24268
rect 36004 24256 36032 24296
rect 36354 24284 36360 24336
rect 36412 24284 36418 24336
rect 38286 24284 38292 24336
rect 38344 24324 38350 24336
rect 39209 24327 39267 24333
rect 39209 24324 39221 24327
rect 38344 24296 39221 24324
rect 38344 24284 38350 24296
rect 39209 24293 39221 24296
rect 39255 24293 39267 24327
rect 39209 24287 39267 24293
rect 39758 24284 39764 24336
rect 39816 24324 39822 24336
rect 40589 24327 40647 24333
rect 40589 24324 40601 24327
rect 39816 24296 40601 24324
rect 39816 24284 39822 24296
rect 40589 24293 40601 24296
rect 40635 24324 40647 24327
rect 41506 24324 41512 24336
rect 40635 24296 41512 24324
rect 40635 24293 40647 24296
rect 40589 24287 40647 24293
rect 41506 24284 41512 24296
rect 41564 24284 41570 24336
rect 42518 24284 42524 24336
rect 42576 24324 42582 24336
rect 47504 24324 47532 24364
rect 48682 24352 48688 24364
rect 48740 24352 48746 24404
rect 48774 24352 48780 24404
rect 48832 24392 48838 24404
rect 49053 24395 49111 24401
rect 49053 24392 49065 24395
rect 48832 24364 49065 24392
rect 48832 24352 48838 24364
rect 49053 24361 49065 24364
rect 49099 24361 49111 24395
rect 49053 24355 49111 24361
rect 49421 24395 49479 24401
rect 49421 24361 49433 24395
rect 49467 24392 49479 24395
rect 49510 24392 49516 24404
rect 49467 24364 49516 24392
rect 49467 24361 49479 24364
rect 49421 24355 49479 24361
rect 49510 24352 49516 24364
rect 49568 24352 49574 24404
rect 49694 24352 49700 24404
rect 49752 24392 49758 24404
rect 50522 24392 50528 24404
rect 49752 24364 50528 24392
rect 49752 24352 49758 24364
rect 50522 24352 50528 24364
rect 50580 24352 50586 24404
rect 50982 24352 50988 24404
rect 51040 24352 51046 24404
rect 51261 24395 51319 24401
rect 51261 24361 51273 24395
rect 51307 24392 51319 24395
rect 53929 24395 53987 24401
rect 53929 24392 53941 24395
rect 51307 24364 53941 24392
rect 51307 24361 51319 24364
rect 51261 24355 51319 24361
rect 53929 24361 53941 24364
rect 53975 24392 53987 24395
rect 54386 24392 54392 24404
rect 53975 24364 54392 24392
rect 53975 24361 53987 24364
rect 53929 24355 53987 24361
rect 42576 24296 47532 24324
rect 48041 24327 48099 24333
rect 42576 24284 42582 24296
rect 48041 24293 48053 24327
rect 48087 24324 48099 24327
rect 48087 24296 49188 24324
rect 48087 24293 48099 24296
rect 48041 24287 48099 24293
rect 36004 24228 36492 24256
rect 34287 24160 34468 24188
rect 34287 24157 34299 24160
rect 34241 24151 34299 24157
rect 34514 24148 34520 24200
rect 34572 24148 34578 24200
rect 35618 24188 35624 24200
rect 34716 24160 35624 24188
rect 34716 24129 34744 24160
rect 35618 24148 35624 24160
rect 35676 24148 35682 24200
rect 36464 24197 36492 24228
rect 36814 24216 36820 24268
rect 36872 24256 36878 24268
rect 39666 24256 39672 24268
rect 36872 24228 39672 24256
rect 36872 24216 36878 24228
rect 39666 24216 39672 24228
rect 39724 24216 39730 24268
rect 39853 24259 39911 24265
rect 39853 24225 39865 24259
rect 39899 24256 39911 24259
rect 41969 24259 42027 24265
rect 39899 24228 40816 24256
rect 39899 24225 39911 24228
rect 39853 24219 39911 24225
rect 36081 24191 36139 24197
rect 36081 24166 36093 24191
rect 36127 24166 36139 24191
rect 36173 24191 36231 24197
rect 33100 24092 33272 24120
rect 33413 24123 33471 24129
rect 33100 24080 33106 24092
rect 33413 24089 33425 24123
rect 33459 24120 33471 24123
rect 34701 24123 34759 24129
rect 34701 24120 34713 24123
rect 33459 24092 34713 24120
rect 33459 24089 33471 24092
rect 33413 24083 33471 24089
rect 34701 24089 34713 24092
rect 34747 24089 34759 24123
rect 34701 24083 34759 24089
rect 30650 24052 30656 24064
rect 30111 24024 30656 24052
rect 30650 24012 30656 24024
rect 30708 24012 30714 24064
rect 30834 24012 30840 24064
rect 30892 24012 30898 24064
rect 31478 24012 31484 24064
rect 31536 24052 31542 24064
rect 33428 24052 33456 24083
rect 35710 24080 35716 24132
rect 35768 24120 35774 24132
rect 35805 24123 35863 24129
rect 35805 24120 35817 24123
rect 35768 24092 35817 24120
rect 35768 24080 35774 24092
rect 35805 24089 35817 24092
rect 35851 24120 35863 24123
rect 35894 24120 35900 24132
rect 35851 24092 35900 24120
rect 35851 24089 35863 24092
rect 35805 24083 35863 24089
rect 35894 24080 35900 24092
rect 35952 24080 35958 24132
rect 36078 24114 36084 24166
rect 36136 24114 36142 24166
rect 36173 24157 36185 24191
rect 36219 24188 36231 24191
rect 36449 24191 36507 24197
rect 36219 24160 36308 24188
rect 36219 24157 36231 24160
rect 36173 24151 36231 24157
rect 36280 24120 36308 24160
rect 36449 24157 36461 24191
rect 36495 24157 36507 24191
rect 36449 24151 36507 24157
rect 36538 24148 36544 24200
rect 36596 24188 36602 24200
rect 36596 24160 36676 24188
rect 36596 24148 36602 24160
rect 36648 24120 36676 24160
rect 36722 24148 36728 24200
rect 36780 24148 36786 24200
rect 36906 24148 36912 24200
rect 36964 24148 36970 24200
rect 37090 24148 37096 24200
rect 37148 24148 37154 24200
rect 39393 24191 39451 24197
rect 39393 24157 39405 24191
rect 39439 24188 39451 24191
rect 39574 24188 39580 24200
rect 39439 24160 39580 24188
rect 39439 24157 39451 24160
rect 39393 24151 39451 24157
rect 39574 24148 39580 24160
rect 39632 24148 39638 24200
rect 39942 24148 39948 24200
rect 40000 24188 40006 24200
rect 40313 24191 40371 24197
rect 40313 24188 40325 24191
rect 40000 24160 40325 24188
rect 40000 24148 40006 24160
rect 40313 24157 40325 24160
rect 40359 24157 40371 24191
rect 40313 24151 40371 24157
rect 40788 24132 40816 24228
rect 41969 24225 41981 24259
rect 42015 24256 42027 24259
rect 42245 24259 42303 24265
rect 42245 24256 42257 24259
rect 42015 24228 42257 24256
rect 42015 24225 42027 24228
rect 41969 24219 42027 24225
rect 42245 24225 42257 24228
rect 42291 24256 42303 24259
rect 43073 24259 43131 24265
rect 43073 24256 43085 24259
rect 42291 24228 43085 24256
rect 42291 24225 42303 24228
rect 42245 24219 42303 24225
rect 43073 24225 43085 24228
rect 43119 24225 43131 24259
rect 43073 24219 43131 24225
rect 45646 24216 45652 24268
rect 45704 24256 45710 24268
rect 46842 24256 46848 24268
rect 45704 24228 46848 24256
rect 45704 24216 45710 24228
rect 41322 24148 41328 24200
rect 41380 24188 41386 24200
rect 41877 24191 41935 24197
rect 41877 24188 41889 24191
rect 41380 24160 41889 24188
rect 41380 24148 41386 24160
rect 41877 24157 41889 24160
rect 41923 24157 41935 24191
rect 41877 24151 41935 24157
rect 42061 24191 42119 24197
rect 42061 24157 42073 24191
rect 42107 24188 42119 24191
rect 42150 24188 42156 24200
rect 42107 24160 42156 24188
rect 42107 24157 42119 24160
rect 42061 24151 42119 24157
rect 42150 24148 42156 24160
rect 42208 24148 42214 24200
rect 42521 24191 42579 24197
rect 42521 24188 42533 24191
rect 42352 24160 42533 24188
rect 36817 24123 36875 24129
rect 36817 24120 36829 24123
rect 36280 24092 36584 24120
rect 36648 24092 36829 24120
rect 31536 24024 33456 24052
rect 31536 24012 31542 24024
rect 33962 24012 33968 24064
rect 34020 24012 34026 24064
rect 36556 24061 36584 24092
rect 36817 24089 36829 24092
rect 36863 24089 36875 24123
rect 36817 24083 36875 24089
rect 36998 24080 37004 24132
rect 37056 24120 37062 24132
rect 39482 24120 39488 24132
rect 37056 24092 39488 24120
rect 37056 24080 37062 24092
rect 39482 24080 39488 24092
rect 39540 24080 39546 24132
rect 40034 24080 40040 24132
rect 40092 24120 40098 24132
rect 40405 24123 40463 24129
rect 40405 24120 40417 24123
rect 40092 24092 40417 24120
rect 40092 24080 40098 24092
rect 40405 24089 40417 24092
rect 40451 24089 40463 24123
rect 40405 24083 40463 24089
rect 40770 24080 40776 24132
rect 40828 24080 40834 24132
rect 41414 24080 41420 24132
rect 41472 24120 41478 24132
rect 42352 24120 42380 24160
rect 42521 24157 42533 24160
rect 42567 24188 42579 24191
rect 43349 24191 43407 24197
rect 43349 24188 43361 24191
rect 42567 24160 43361 24188
rect 42567 24157 42579 24160
rect 42521 24151 42579 24157
rect 43349 24157 43361 24160
rect 43395 24188 43407 24191
rect 43714 24188 43720 24200
rect 43395 24160 43720 24188
rect 43395 24157 43407 24160
rect 43349 24151 43407 24157
rect 43714 24148 43720 24160
rect 43772 24148 43778 24200
rect 46216 24197 46244 24228
rect 46842 24216 46848 24228
rect 46900 24256 46906 24268
rect 47213 24259 47271 24265
rect 47213 24256 47225 24259
rect 46900 24228 47225 24256
rect 46900 24216 46906 24228
rect 47213 24225 47225 24228
rect 47259 24256 47271 24259
rect 48406 24256 48412 24268
rect 47259 24228 48412 24256
rect 47259 24225 47271 24228
rect 47213 24219 47271 24225
rect 48406 24216 48412 24228
rect 48464 24216 48470 24268
rect 48682 24216 48688 24268
rect 48740 24256 48746 24268
rect 48958 24256 48964 24268
rect 48740 24228 48964 24256
rect 48740 24216 48746 24228
rect 48958 24216 48964 24228
rect 49016 24216 49022 24268
rect 49160 24265 49188 24296
rect 50706 24284 50712 24336
rect 50764 24324 50770 24336
rect 51276 24324 51304 24355
rect 54386 24352 54392 24364
rect 54444 24352 54450 24404
rect 56137 24395 56195 24401
rect 56137 24361 56149 24395
rect 56183 24392 56195 24395
rect 56226 24392 56232 24404
rect 56183 24364 56232 24392
rect 56183 24361 56195 24364
rect 56137 24355 56195 24361
rect 56226 24352 56232 24364
rect 56284 24352 56290 24404
rect 50764 24296 51304 24324
rect 50764 24284 50770 24296
rect 53834 24284 53840 24336
rect 53892 24324 53898 24336
rect 57698 24324 57704 24336
rect 53892 24296 57704 24324
rect 53892 24284 53898 24296
rect 49145 24259 49203 24265
rect 49145 24225 49157 24259
rect 49191 24225 49203 24259
rect 49145 24219 49203 24225
rect 49878 24216 49884 24268
rect 49936 24216 49942 24268
rect 52362 24216 52368 24268
rect 52420 24256 52426 24268
rect 52420 24228 54064 24256
rect 52420 24216 52426 24228
rect 46201 24191 46259 24197
rect 46201 24157 46213 24191
rect 46247 24157 46259 24191
rect 47397 24191 47455 24197
rect 47397 24188 47409 24191
rect 46201 24151 46259 24157
rect 46308 24160 47409 24188
rect 41472 24092 42380 24120
rect 41472 24080 41478 24092
rect 42426 24080 42432 24132
rect 42484 24080 42490 24132
rect 42978 24080 42984 24132
rect 43036 24080 43042 24132
rect 43254 24080 43260 24132
rect 43312 24080 43318 24132
rect 45278 24080 45284 24132
rect 45336 24120 45342 24132
rect 46308 24120 46336 24160
rect 47397 24157 47409 24160
rect 47443 24157 47455 24191
rect 47397 24151 47455 24157
rect 47490 24191 47548 24197
rect 47490 24157 47502 24191
rect 47536 24157 47548 24191
rect 47490 24151 47548 24157
rect 47862 24191 47920 24197
rect 47862 24157 47874 24191
rect 47908 24157 47920 24191
rect 47862 24151 47920 24157
rect 49053 24191 49111 24197
rect 49053 24157 49065 24191
rect 49099 24188 49111 24191
rect 49418 24188 49424 24200
rect 49099 24160 49424 24188
rect 49099 24157 49111 24160
rect 49053 24151 49111 24157
rect 45336 24092 46336 24120
rect 45336 24080 45342 24092
rect 46382 24080 46388 24132
rect 46440 24080 46446 24132
rect 46934 24080 46940 24132
rect 46992 24120 46998 24132
rect 47302 24120 47308 24132
rect 46992 24092 47308 24120
rect 46992 24080 46998 24092
rect 47302 24080 47308 24092
rect 47360 24120 47366 24132
rect 47504 24120 47532 24151
rect 47360 24092 47532 24120
rect 47360 24080 47366 24092
rect 47578 24080 47584 24132
rect 47636 24120 47642 24132
rect 47673 24123 47731 24129
rect 47673 24120 47685 24123
rect 47636 24092 47685 24120
rect 47636 24080 47642 24092
rect 47673 24089 47685 24092
rect 47719 24089 47731 24123
rect 47673 24083 47731 24089
rect 47762 24080 47768 24132
rect 47820 24080 47826 24132
rect 36541 24055 36599 24061
rect 36541 24021 36553 24055
rect 36587 24021 36599 24055
rect 36541 24015 36599 24021
rect 38746 24012 38752 24064
rect 38804 24012 38810 24064
rect 39114 24012 39120 24064
rect 39172 24052 39178 24064
rect 39942 24052 39948 24064
rect 39172 24024 39948 24052
rect 39172 24012 39178 24024
rect 39942 24012 39948 24024
rect 40000 24012 40006 24064
rect 43162 24012 43168 24064
rect 43220 24052 43226 24064
rect 43901 24055 43959 24061
rect 43901 24052 43913 24055
rect 43220 24024 43913 24052
rect 43220 24012 43226 24024
rect 43901 24021 43913 24024
rect 43947 24021 43959 24055
rect 43901 24015 43959 24021
rect 44818 24012 44824 24064
rect 44876 24012 44882 24064
rect 47118 24012 47124 24064
rect 47176 24052 47182 24064
rect 47872 24052 47900 24151
rect 49418 24148 49424 24160
rect 49476 24148 49482 24200
rect 49896 24188 49924 24216
rect 54036 24200 54064 24228
rect 54110 24216 54116 24268
rect 54168 24256 54174 24268
rect 55214 24256 55220 24268
rect 54168 24228 55220 24256
rect 54168 24216 54174 24228
rect 55214 24216 55220 24228
rect 55272 24256 55278 24268
rect 56410 24256 56416 24268
rect 55272 24228 56416 24256
rect 55272 24216 55278 24228
rect 56410 24216 56416 24228
rect 56468 24256 56474 24268
rect 56612 24265 56640 24296
rect 57698 24284 57704 24296
rect 57756 24284 57762 24336
rect 56505 24259 56563 24265
rect 56505 24256 56517 24259
rect 56468 24228 56517 24256
rect 56468 24216 56474 24228
rect 56505 24225 56517 24228
rect 56551 24225 56563 24259
rect 56505 24219 56563 24225
rect 56597 24259 56655 24265
rect 56597 24225 56609 24259
rect 56643 24225 56655 24259
rect 56597 24219 56655 24225
rect 50706 24188 50712 24200
rect 49896 24160 50712 24188
rect 50706 24148 50712 24160
rect 50764 24148 50770 24200
rect 50798 24148 50804 24200
rect 50856 24148 50862 24200
rect 51077 24191 51135 24197
rect 51077 24157 51089 24191
rect 51123 24188 51135 24191
rect 51629 24191 51687 24197
rect 51629 24188 51641 24191
rect 51123 24160 51641 24188
rect 51123 24157 51135 24160
rect 51077 24151 51135 24157
rect 51629 24157 51641 24160
rect 51675 24157 51687 24191
rect 51629 24151 51687 24157
rect 52178 24148 52184 24200
rect 52236 24188 52242 24200
rect 53193 24191 53251 24197
rect 53193 24188 53205 24191
rect 52236 24160 53205 24188
rect 52236 24148 52242 24160
rect 53193 24157 53205 24160
rect 53239 24157 53251 24191
rect 53193 24151 53251 24157
rect 53558 24148 53564 24200
rect 53616 24148 53622 24200
rect 53834 24188 53840 24200
rect 53668 24160 53840 24188
rect 49970 24080 49976 24132
rect 50028 24120 50034 24132
rect 50028 24092 51764 24120
rect 50028 24080 50034 24092
rect 47176 24024 47900 24052
rect 47176 24012 47182 24024
rect 48130 24012 48136 24064
rect 48188 24012 48194 24064
rect 48314 24012 48320 24064
rect 48372 24052 48378 24064
rect 48409 24055 48467 24061
rect 48409 24052 48421 24055
rect 48372 24024 48421 24052
rect 48372 24012 48378 24024
rect 48409 24021 48421 24024
rect 48455 24052 48467 24055
rect 48590 24052 48596 24064
rect 48455 24024 48596 24052
rect 48455 24021 48467 24024
rect 48409 24015 48467 24021
rect 48590 24012 48596 24024
rect 48648 24012 48654 24064
rect 50525 24055 50583 24061
rect 50525 24021 50537 24055
rect 50571 24052 50583 24055
rect 50706 24052 50712 24064
rect 50571 24024 50712 24052
rect 50571 24021 50583 24024
rect 50525 24015 50583 24021
rect 50706 24012 50712 24024
rect 50764 24012 50770 24064
rect 51736 24052 51764 24092
rect 53374 24080 53380 24132
rect 53432 24080 53438 24132
rect 53469 24123 53527 24129
rect 53469 24089 53481 24123
rect 53515 24120 53527 24123
rect 53668 24120 53696 24160
rect 53834 24148 53840 24160
rect 53892 24148 53898 24200
rect 54018 24148 54024 24200
rect 54076 24148 54082 24200
rect 54297 24191 54355 24197
rect 54297 24157 54309 24191
rect 54343 24157 54355 24191
rect 54297 24151 54355 24157
rect 54312 24120 54340 24151
rect 54386 24148 54392 24200
rect 54444 24188 54450 24200
rect 54846 24188 54852 24200
rect 54444 24160 54852 24188
rect 54444 24148 54450 24160
rect 54846 24148 54852 24160
rect 54904 24148 54910 24200
rect 56318 24148 56324 24200
rect 56376 24148 56382 24200
rect 57422 24148 57428 24200
rect 57480 24148 57486 24200
rect 53515 24092 53696 24120
rect 53760 24092 54340 24120
rect 53515 24089 53527 24092
rect 53469 24083 53527 24089
rect 53484 24052 53512 24083
rect 53760 24061 53788 24092
rect 51736 24024 53512 24052
rect 53745 24055 53803 24061
rect 53745 24021 53757 24055
rect 53791 24021 53803 24055
rect 53745 24015 53803 24021
rect 54294 24012 54300 24064
rect 54352 24052 54358 24064
rect 54573 24055 54631 24061
rect 54573 24052 54585 24055
rect 54352 24024 54585 24052
rect 54352 24012 54358 24024
rect 54573 24021 54585 24024
rect 54619 24021 54631 24055
rect 54573 24015 54631 24021
rect 54754 24012 54760 24064
rect 54812 24052 54818 24064
rect 55769 24055 55827 24061
rect 55769 24052 55781 24055
rect 54812 24024 55781 24052
rect 54812 24012 54818 24024
rect 55769 24021 55781 24024
rect 55815 24052 55827 24055
rect 56502 24052 56508 24064
rect 55815 24024 56508 24052
rect 55815 24021 55827 24024
rect 55769 24015 55827 24021
rect 56502 24012 56508 24024
rect 56560 24012 56566 24064
rect 57609 24055 57667 24061
rect 57609 24021 57621 24055
rect 57655 24052 57667 24055
rect 58250 24052 58256 24064
rect 57655 24024 58256 24052
rect 57655 24021 57667 24024
rect 57609 24015 57667 24021
rect 58250 24012 58256 24024
rect 58308 24012 58314 24064
rect 1104 23962 58880 23984
rect 1104 23910 4874 23962
rect 4926 23910 4938 23962
rect 4990 23910 5002 23962
rect 5054 23910 5066 23962
rect 5118 23910 5130 23962
rect 5182 23910 35594 23962
rect 35646 23910 35658 23962
rect 35710 23910 35722 23962
rect 35774 23910 35786 23962
rect 35838 23910 35850 23962
rect 35902 23910 58880 23962
rect 1104 23888 58880 23910
rect 19518 23808 19524 23860
rect 19576 23848 19582 23860
rect 20073 23851 20131 23857
rect 20073 23848 20085 23851
rect 19576 23820 20085 23848
rect 19576 23808 19582 23820
rect 20073 23817 20085 23820
rect 20119 23817 20131 23851
rect 20990 23848 20996 23860
rect 20073 23811 20131 23817
rect 20364 23820 20996 23848
rect 18506 23740 18512 23792
rect 18564 23740 18570 23792
rect 20364 23789 20392 23820
rect 20990 23808 20996 23820
rect 21048 23808 21054 23860
rect 22922 23848 22928 23860
rect 21468 23820 22928 23848
rect 20349 23783 20407 23789
rect 20349 23749 20361 23783
rect 20395 23749 20407 23783
rect 20349 23743 20407 23749
rect 20441 23783 20499 23789
rect 20441 23749 20453 23783
rect 20487 23780 20499 23783
rect 20806 23780 20812 23792
rect 20487 23752 20812 23780
rect 20487 23749 20499 23752
rect 20441 23743 20499 23749
rect 20806 23740 20812 23752
rect 20864 23740 20870 23792
rect 19518 23672 19524 23724
rect 19576 23712 19582 23724
rect 19576 23684 19642 23712
rect 19576 23672 19582 23684
rect 19794 23672 19800 23724
rect 19852 23712 19858 23724
rect 20257 23715 20315 23721
rect 20257 23712 20269 23715
rect 19852 23684 20269 23712
rect 19852 23672 19858 23684
rect 20257 23681 20269 23684
rect 20303 23681 20315 23715
rect 20257 23675 20315 23681
rect 20622 23672 20628 23724
rect 20680 23712 20686 23724
rect 21468 23712 21496 23820
rect 22922 23808 22928 23820
rect 22980 23808 22986 23860
rect 23106 23808 23112 23860
rect 23164 23848 23170 23860
rect 23477 23851 23535 23857
rect 23477 23848 23489 23851
rect 23164 23820 23489 23848
rect 23164 23808 23170 23820
rect 23477 23817 23489 23820
rect 23523 23817 23535 23851
rect 23477 23811 23535 23817
rect 25038 23808 25044 23860
rect 25096 23808 25102 23860
rect 25222 23808 25228 23860
rect 25280 23848 25286 23860
rect 25501 23851 25559 23857
rect 25501 23848 25513 23851
rect 25280 23820 25513 23848
rect 25280 23808 25286 23820
rect 25501 23817 25513 23820
rect 25547 23817 25559 23851
rect 26602 23848 26608 23860
rect 25501 23811 25559 23817
rect 26344 23820 26608 23848
rect 22094 23780 22100 23792
rect 21560 23752 22100 23780
rect 21560 23721 21588 23752
rect 22094 23740 22100 23752
rect 22152 23780 22158 23792
rect 22830 23780 22836 23792
rect 22152 23752 22836 23780
rect 22152 23740 22158 23752
rect 22830 23740 22836 23752
rect 22888 23740 22894 23792
rect 24765 23783 24823 23789
rect 24765 23780 24777 23783
rect 24044 23752 24777 23780
rect 24044 23724 24072 23752
rect 24765 23749 24777 23752
rect 24811 23749 24823 23783
rect 24765 23743 24823 23749
rect 25590 23740 25596 23792
rect 25648 23780 25654 23792
rect 25648 23752 25820 23780
rect 25648 23740 25654 23752
rect 20680 23684 21496 23712
rect 21545 23715 21603 23721
rect 20680 23672 20686 23684
rect 21545 23681 21557 23715
rect 21591 23681 21603 23715
rect 21545 23675 21603 23681
rect 18233 23647 18291 23653
rect 18233 23613 18245 23647
rect 18279 23613 18291 23647
rect 18233 23607 18291 23613
rect 18248 23508 18276 23607
rect 19242 23604 19248 23656
rect 19300 23644 19306 23656
rect 21560 23644 21588 23675
rect 22002 23672 22008 23724
rect 22060 23712 22066 23724
rect 23017 23715 23075 23721
rect 23017 23712 23029 23715
rect 22060 23684 23029 23712
rect 22060 23672 22066 23684
rect 23017 23681 23029 23684
rect 23063 23681 23075 23715
rect 23017 23675 23075 23681
rect 23566 23672 23572 23724
rect 23624 23712 23630 23724
rect 23661 23715 23719 23721
rect 23661 23712 23673 23715
rect 23624 23684 23673 23712
rect 23624 23672 23630 23684
rect 23661 23681 23673 23684
rect 23707 23681 23719 23715
rect 23661 23675 23719 23681
rect 23750 23672 23756 23724
rect 23808 23672 23814 23724
rect 23842 23672 23848 23724
rect 23900 23672 23906 23724
rect 24026 23672 24032 23724
rect 24084 23672 24090 23724
rect 24489 23715 24547 23721
rect 24489 23681 24501 23715
rect 24535 23681 24547 23715
rect 24489 23675 24547 23681
rect 24673 23715 24731 23721
rect 24673 23681 24685 23715
rect 24719 23681 24731 23715
rect 24673 23675 24731 23681
rect 24857 23715 24915 23721
rect 24857 23681 24869 23715
rect 24903 23712 24915 23715
rect 25225 23715 25283 23721
rect 25225 23712 25237 23715
rect 24903 23684 25237 23712
rect 24903 23681 24915 23684
rect 24857 23675 24915 23681
rect 25225 23681 25237 23684
rect 25271 23712 25283 23715
rect 25314 23712 25320 23724
rect 25271 23684 25320 23712
rect 25271 23681 25283 23684
rect 25225 23675 25283 23681
rect 19300 23616 21588 23644
rect 19300 23604 19306 23616
rect 22278 23604 22284 23656
rect 22336 23644 22342 23656
rect 23584 23644 23612 23672
rect 22336 23616 23612 23644
rect 22336 23604 22342 23616
rect 19242 23508 19248 23520
rect 18248 23480 19248 23508
rect 19242 23468 19248 23480
rect 19300 23468 19306 23520
rect 19978 23468 19984 23520
rect 20036 23508 20042 23520
rect 24504 23508 24532 23675
rect 24688 23644 24716 23675
rect 25314 23672 25320 23684
rect 25372 23672 25378 23724
rect 25682 23672 25688 23724
rect 25740 23672 25746 23724
rect 25792 23721 25820 23752
rect 26344 23721 26372 23820
rect 26602 23808 26608 23820
rect 26660 23848 26666 23860
rect 27249 23851 27307 23857
rect 27249 23848 27261 23851
rect 26660 23820 27261 23848
rect 26660 23808 26666 23820
rect 27249 23817 27261 23820
rect 27295 23848 27307 23851
rect 31662 23848 31668 23860
rect 27295 23820 31668 23848
rect 27295 23817 27307 23820
rect 27249 23811 27307 23817
rect 31662 23808 31668 23820
rect 31720 23808 31726 23860
rect 31754 23808 31760 23860
rect 31812 23848 31818 23860
rect 32214 23848 32220 23860
rect 31812 23820 32220 23848
rect 31812 23808 31818 23820
rect 32214 23808 32220 23820
rect 32272 23808 32278 23860
rect 33134 23808 33140 23860
rect 33192 23848 33198 23860
rect 33413 23851 33471 23857
rect 33413 23848 33425 23851
rect 33192 23820 33425 23848
rect 33192 23808 33198 23820
rect 33413 23817 33425 23820
rect 33459 23817 33471 23851
rect 34793 23851 34851 23857
rect 33413 23811 33471 23817
rect 33520 23820 34284 23848
rect 26418 23740 26424 23792
rect 26476 23740 26482 23792
rect 26513 23783 26571 23789
rect 26513 23749 26525 23783
rect 26559 23780 26571 23783
rect 27062 23780 27068 23792
rect 26559 23752 27068 23780
rect 26559 23749 26571 23752
rect 26513 23743 26571 23749
rect 27062 23740 27068 23752
rect 27120 23740 27126 23792
rect 27540 23752 28028 23780
rect 25777 23715 25835 23721
rect 25777 23681 25789 23715
rect 25823 23681 25835 23715
rect 25961 23715 26019 23721
rect 25961 23712 25973 23715
rect 25777 23675 25835 23681
rect 25884 23684 25973 23712
rect 24688 23616 25452 23644
rect 20036 23480 24532 23508
rect 20036 23468 20042 23480
rect 25314 23468 25320 23520
rect 25372 23508 25378 23520
rect 25424 23517 25452 23616
rect 25884 23576 25912 23684
rect 25961 23681 25973 23684
rect 26007 23681 26019 23715
rect 25961 23675 26019 23681
rect 26053 23715 26111 23721
rect 26053 23681 26065 23715
rect 26099 23712 26111 23715
rect 26329 23715 26387 23721
rect 26099 23684 26188 23712
rect 26099 23681 26111 23684
rect 26053 23675 26111 23681
rect 26160 23585 26188 23684
rect 26329 23681 26341 23715
rect 26375 23681 26387 23715
rect 26329 23675 26387 23681
rect 26694 23672 26700 23724
rect 26752 23672 26758 23724
rect 27430 23672 27436 23724
rect 27488 23712 27494 23724
rect 27540 23721 27568 23752
rect 27525 23715 27583 23721
rect 27525 23712 27537 23715
rect 27488 23684 27537 23712
rect 27488 23672 27494 23684
rect 27525 23681 27537 23684
rect 27571 23681 27583 23715
rect 27525 23675 27583 23681
rect 27706 23672 27712 23724
rect 27764 23672 27770 23724
rect 27798 23672 27804 23724
rect 27856 23672 27862 23724
rect 27893 23715 27951 23721
rect 27893 23681 27905 23715
rect 27939 23681 27951 23715
rect 28000 23712 28028 23752
rect 28074 23740 28080 23792
rect 28132 23780 28138 23792
rect 32401 23783 32459 23789
rect 28132 23752 28764 23780
rect 28132 23740 28138 23752
rect 28258 23712 28264 23724
rect 28000 23684 28264 23712
rect 27893 23675 27951 23681
rect 27908 23644 27936 23675
rect 28258 23672 28264 23684
rect 28316 23672 28322 23724
rect 28353 23715 28411 23721
rect 28353 23681 28365 23715
rect 28399 23681 28411 23715
rect 28353 23675 28411 23681
rect 27982 23644 27988 23656
rect 27908 23616 27988 23644
rect 27982 23604 27988 23616
rect 28040 23604 28046 23656
rect 28368 23644 28396 23675
rect 28442 23672 28448 23724
rect 28500 23672 28506 23724
rect 28736 23721 28764 23752
rect 32401 23749 32413 23783
rect 32447 23780 32459 23783
rect 32582 23780 32588 23792
rect 32447 23752 32588 23780
rect 32447 23749 32459 23752
rect 32401 23743 32459 23749
rect 32582 23740 32588 23752
rect 32640 23740 32646 23792
rect 32950 23740 32956 23792
rect 33008 23780 33014 23792
rect 33520 23780 33548 23820
rect 33008 23752 33548 23780
rect 33581 23783 33639 23789
rect 33008 23740 33014 23752
rect 33581 23749 33593 23783
rect 33627 23780 33639 23783
rect 33686 23780 33692 23792
rect 33627 23752 33692 23780
rect 33627 23749 33639 23752
rect 33581 23743 33639 23749
rect 33686 23740 33692 23752
rect 33744 23740 33750 23792
rect 33781 23783 33839 23789
rect 33781 23749 33793 23783
rect 33827 23749 33839 23783
rect 33781 23743 33839 23749
rect 28537 23715 28595 23721
rect 28537 23681 28549 23715
rect 28583 23681 28595 23715
rect 28537 23675 28595 23681
rect 28721 23715 28779 23721
rect 28721 23681 28733 23715
rect 28767 23681 28779 23715
rect 28721 23675 28779 23681
rect 28552 23644 28580 23675
rect 32122 23672 32128 23724
rect 32180 23672 32186 23724
rect 32214 23672 32220 23724
rect 32272 23712 32278 23724
rect 32309 23715 32367 23721
rect 32309 23712 32321 23715
rect 32272 23684 32321 23712
rect 32272 23672 32278 23684
rect 32309 23681 32321 23684
rect 32355 23681 32367 23715
rect 32309 23675 32367 23681
rect 32493 23715 32551 23721
rect 32493 23681 32505 23715
rect 32539 23712 32551 23715
rect 33134 23712 33140 23724
rect 32539 23684 33140 23712
rect 32539 23681 32551 23684
rect 32493 23675 32551 23681
rect 33134 23672 33140 23684
rect 33192 23712 33198 23724
rect 33410 23712 33416 23724
rect 33192 23684 33416 23712
rect 33192 23672 33198 23684
rect 33410 23672 33416 23684
rect 33468 23672 33474 23724
rect 32140 23644 32168 23672
rect 33796 23644 33824 23743
rect 34256 23721 34284 23820
rect 34793 23817 34805 23851
rect 34839 23817 34851 23851
rect 34793 23811 34851 23817
rect 34330 23740 34336 23792
rect 34388 23780 34394 23792
rect 34425 23783 34483 23789
rect 34425 23780 34437 23783
rect 34388 23752 34437 23780
rect 34388 23740 34394 23752
rect 34425 23749 34437 23752
rect 34471 23749 34483 23783
rect 34425 23743 34483 23749
rect 34517 23783 34575 23789
rect 34517 23749 34529 23783
rect 34563 23780 34575 23783
rect 34808 23780 34836 23811
rect 34974 23808 34980 23860
rect 35032 23808 35038 23860
rect 35434 23808 35440 23860
rect 35492 23848 35498 23860
rect 37001 23851 37059 23857
rect 37001 23848 37013 23851
rect 35492 23820 37013 23848
rect 35492 23808 35498 23820
rect 37001 23817 37013 23820
rect 37047 23848 37059 23851
rect 37918 23848 37924 23860
rect 37047 23820 37924 23848
rect 37047 23817 37059 23820
rect 37001 23811 37059 23817
rect 37918 23808 37924 23820
rect 37976 23808 37982 23860
rect 38010 23808 38016 23860
rect 38068 23848 38074 23860
rect 38378 23848 38384 23860
rect 38068 23820 38384 23848
rect 38068 23808 38074 23820
rect 34563 23752 34744 23780
rect 34808 23752 35664 23780
rect 34563 23749 34575 23752
rect 34517 23743 34575 23749
rect 34241 23715 34299 23721
rect 34241 23681 34253 23715
rect 34287 23681 34299 23715
rect 34241 23675 34299 23681
rect 34609 23715 34667 23721
rect 34609 23681 34621 23715
rect 34655 23681 34667 23715
rect 34716 23712 34744 23752
rect 34882 23712 34888 23724
rect 34716 23684 34888 23712
rect 34609 23675 34667 23681
rect 28368 23616 28520 23644
rect 28552 23616 29040 23644
rect 32140 23616 33824 23644
rect 26145 23579 26203 23585
rect 25884 23548 26096 23576
rect 25409 23511 25467 23517
rect 25409 23508 25421 23511
rect 25372 23480 25421 23508
rect 25372 23468 25378 23480
rect 25409 23477 25421 23480
rect 25455 23508 25467 23511
rect 25958 23508 25964 23520
rect 25455 23480 25964 23508
rect 25455 23477 25467 23480
rect 25409 23471 25467 23477
rect 25958 23468 25964 23480
rect 26016 23468 26022 23520
rect 26068 23508 26096 23548
rect 26145 23545 26157 23579
rect 26191 23545 26203 23579
rect 26145 23539 26203 23545
rect 28077 23579 28135 23585
rect 28077 23545 28089 23579
rect 28123 23576 28135 23579
rect 28350 23576 28356 23588
rect 28123 23548 28356 23576
rect 28123 23545 28135 23548
rect 28077 23539 28135 23545
rect 28350 23536 28356 23548
rect 28408 23536 28414 23588
rect 28492 23576 28520 23616
rect 28902 23576 28908 23588
rect 28492 23548 28908 23576
rect 28902 23536 28908 23548
rect 28960 23536 28966 23588
rect 29012 23520 29040 23616
rect 30006 23536 30012 23588
rect 30064 23576 30070 23588
rect 34057 23579 34115 23585
rect 34057 23576 34069 23579
rect 30064 23548 34069 23576
rect 30064 23536 30070 23548
rect 34057 23545 34069 23548
rect 34103 23576 34115 23579
rect 34624 23576 34652 23675
rect 34882 23672 34888 23684
rect 34940 23672 34946 23724
rect 35158 23721 35164 23724
rect 35156 23712 35164 23721
rect 35119 23684 35164 23712
rect 35156 23675 35164 23684
rect 35158 23672 35164 23675
rect 35216 23672 35222 23724
rect 35250 23672 35256 23724
rect 35308 23672 35314 23724
rect 35345 23715 35403 23721
rect 35345 23681 35357 23715
rect 35391 23712 35403 23715
rect 35434 23712 35440 23724
rect 35391 23684 35440 23712
rect 35391 23681 35403 23684
rect 35345 23675 35403 23681
rect 35434 23672 35440 23684
rect 35492 23672 35498 23724
rect 35636 23721 35664 23752
rect 36630 23740 36636 23792
rect 36688 23740 36694 23792
rect 36814 23740 36820 23792
rect 36872 23740 36878 23792
rect 35528 23715 35586 23721
rect 35528 23681 35540 23715
rect 35574 23681 35586 23715
rect 35528 23675 35586 23681
rect 35621 23715 35679 23721
rect 35621 23681 35633 23715
rect 35667 23681 35679 23715
rect 35621 23675 35679 23681
rect 34790 23604 34796 23656
rect 34848 23644 34854 23656
rect 35268 23644 35296 23672
rect 34848 23616 35296 23644
rect 35544 23644 35572 23675
rect 38102 23672 38108 23724
rect 38160 23672 38166 23724
rect 38212 23721 38240 23820
rect 38378 23808 38384 23820
rect 38436 23848 38442 23860
rect 39850 23848 39856 23860
rect 38436 23820 39856 23848
rect 38436 23808 38442 23820
rect 39850 23808 39856 23820
rect 39908 23808 39914 23860
rect 40034 23808 40040 23860
rect 40092 23848 40098 23860
rect 45113 23851 45171 23857
rect 45113 23848 45125 23851
rect 40092 23820 45125 23848
rect 40092 23808 40098 23820
rect 38654 23740 38660 23792
rect 38712 23780 38718 23792
rect 38933 23783 38991 23789
rect 38933 23780 38945 23783
rect 38712 23752 38945 23780
rect 38712 23740 38718 23752
rect 38933 23749 38945 23752
rect 38979 23780 38991 23783
rect 39485 23783 39543 23789
rect 38979 23752 39160 23780
rect 38979 23749 38991 23752
rect 38933 23743 38991 23749
rect 38197 23715 38255 23721
rect 38197 23681 38209 23715
rect 38243 23681 38255 23715
rect 38197 23675 38255 23681
rect 38286 23672 38292 23724
rect 38344 23712 38350 23724
rect 39025 23715 39083 23721
rect 39025 23712 39037 23715
rect 38344 23684 39037 23712
rect 38344 23672 38350 23684
rect 39025 23681 39037 23684
rect 39071 23681 39083 23715
rect 39132 23712 39160 23752
rect 39485 23749 39497 23783
rect 39531 23780 39543 23783
rect 39666 23780 39672 23792
rect 39531 23752 39672 23780
rect 39531 23749 39543 23752
rect 39485 23743 39543 23749
rect 39666 23740 39672 23752
rect 39724 23740 39730 23792
rect 39758 23740 39764 23792
rect 39816 23740 39822 23792
rect 40494 23740 40500 23792
rect 40552 23780 40558 23792
rect 42518 23780 42524 23792
rect 40552 23752 42524 23780
rect 40552 23740 40558 23752
rect 42518 23740 42524 23752
rect 42576 23740 42582 23792
rect 42613 23783 42671 23789
rect 42613 23749 42625 23783
rect 42659 23780 42671 23783
rect 42886 23780 42892 23792
rect 42659 23752 42892 23780
rect 42659 23749 42671 23752
rect 42613 23743 42671 23749
rect 42886 23740 42892 23752
rect 42944 23740 42950 23792
rect 43162 23740 43168 23792
rect 43220 23780 43226 23792
rect 43901 23783 43959 23789
rect 43901 23780 43913 23783
rect 43220 23752 43913 23780
rect 43220 23740 43226 23752
rect 43901 23749 43913 23752
rect 43947 23749 43959 23783
rect 43901 23743 43959 23749
rect 39206 23712 39212 23724
rect 39132 23684 39212 23712
rect 39025 23675 39083 23681
rect 39206 23672 39212 23684
rect 39264 23712 39270 23724
rect 39853 23715 39911 23721
rect 39853 23712 39865 23715
rect 39264 23684 39865 23712
rect 39264 23672 39270 23684
rect 39853 23681 39865 23684
rect 39899 23681 39911 23715
rect 39853 23675 39911 23681
rect 42702 23672 42708 23724
rect 42760 23672 42766 23724
rect 42794 23672 42800 23724
rect 42852 23712 42858 23724
rect 44560 23721 44588 23820
rect 45113 23817 45125 23820
rect 45159 23817 45171 23851
rect 45113 23811 45171 23817
rect 45278 23808 45284 23860
rect 45336 23808 45342 23860
rect 46106 23808 46112 23860
rect 46164 23848 46170 23860
rect 46385 23851 46443 23857
rect 46385 23848 46397 23851
rect 46164 23820 46397 23848
rect 46164 23808 46170 23820
rect 46385 23817 46397 23820
rect 46431 23817 46443 23851
rect 46385 23811 46443 23817
rect 47854 23808 47860 23860
rect 47912 23848 47918 23860
rect 47912 23820 48544 23848
rect 47912 23808 47918 23820
rect 44818 23740 44824 23792
rect 44876 23780 44882 23792
rect 44913 23783 44971 23789
rect 44913 23780 44925 23783
rect 44876 23752 44925 23780
rect 44876 23740 44882 23752
rect 44913 23749 44925 23752
rect 44959 23780 44971 23783
rect 45370 23780 45376 23792
rect 44959 23752 45376 23780
rect 44959 23749 44971 23752
rect 44913 23743 44971 23749
rect 45370 23740 45376 23752
rect 45428 23780 45434 23792
rect 45557 23783 45615 23789
rect 45557 23780 45569 23783
rect 45428 23752 45569 23780
rect 45428 23740 45434 23752
rect 45557 23749 45569 23752
rect 45603 23749 45615 23783
rect 45557 23743 45615 23749
rect 46658 23740 46664 23792
rect 46716 23780 46722 23792
rect 48516 23789 48544 23820
rect 48774 23808 48780 23860
rect 48832 23808 48838 23860
rect 49142 23808 49148 23860
rect 49200 23848 49206 23860
rect 49329 23851 49387 23857
rect 49329 23848 49341 23851
rect 49200 23820 49341 23848
rect 49200 23808 49206 23820
rect 49329 23817 49341 23820
rect 49375 23848 49387 23851
rect 52178 23848 52184 23860
rect 49375 23820 50016 23848
rect 49375 23817 49387 23820
rect 49329 23811 49387 23817
rect 49988 23792 50016 23820
rect 50080 23820 52184 23848
rect 48501 23783 48559 23789
rect 46716 23752 48268 23780
rect 46716 23740 46722 23752
rect 43349 23715 43407 23721
rect 43349 23712 43361 23715
rect 42852 23684 43361 23712
rect 42852 23672 42858 23684
rect 43349 23681 43361 23684
rect 43395 23681 43407 23715
rect 43349 23675 43407 23681
rect 44545 23715 44603 23721
rect 44545 23681 44557 23715
rect 44591 23681 44603 23715
rect 44545 23675 44603 23681
rect 45186 23672 45192 23724
rect 45244 23712 45250 23724
rect 46523 23715 46581 23721
rect 46523 23712 46535 23715
rect 45244 23684 46535 23712
rect 45244 23672 45250 23684
rect 46523 23681 46535 23684
rect 46569 23681 46581 23715
rect 46523 23675 46581 23681
rect 46750 23672 46756 23724
rect 46808 23672 46814 23724
rect 46934 23672 46940 23724
rect 46992 23672 46998 23724
rect 47026 23672 47032 23724
rect 47084 23672 47090 23724
rect 47581 23715 47639 23721
rect 47581 23681 47593 23715
rect 47627 23712 47639 23715
rect 47670 23712 47676 23724
rect 47627 23684 47676 23712
rect 47627 23681 47639 23684
rect 47581 23675 47639 23681
rect 47670 23672 47676 23684
rect 47728 23672 47734 23724
rect 47762 23672 47768 23724
rect 47820 23672 47826 23724
rect 47854 23672 47860 23724
rect 47912 23672 47918 23724
rect 47946 23672 47952 23724
rect 48004 23672 48010 23724
rect 48240 23721 48268 23752
rect 48501 23749 48513 23783
rect 48547 23749 48559 23783
rect 48501 23743 48559 23749
rect 49970 23740 49976 23792
rect 50028 23740 50034 23792
rect 50080 23789 50108 23820
rect 52178 23808 52184 23820
rect 52236 23808 52242 23860
rect 53374 23808 53380 23860
rect 53432 23848 53438 23860
rect 54202 23848 54208 23860
rect 53432 23820 54208 23848
rect 53432 23808 53438 23820
rect 54202 23808 54208 23820
rect 54260 23848 54266 23860
rect 54662 23848 54668 23860
rect 54260 23820 54668 23848
rect 54260 23808 54266 23820
rect 54662 23808 54668 23820
rect 54720 23808 54726 23860
rect 55306 23808 55312 23860
rect 55364 23848 55370 23860
rect 55861 23851 55919 23857
rect 55861 23848 55873 23851
rect 55364 23820 55873 23848
rect 55364 23808 55370 23820
rect 55861 23817 55873 23820
rect 55907 23817 55919 23851
rect 55861 23811 55919 23817
rect 50065 23783 50123 23789
rect 50065 23749 50077 23783
rect 50111 23749 50123 23783
rect 50065 23743 50123 23749
rect 50706 23740 50712 23792
rect 50764 23740 50770 23792
rect 51442 23740 51448 23792
rect 51500 23740 51506 23792
rect 48225 23715 48283 23721
rect 48225 23681 48237 23715
rect 48271 23681 48283 23715
rect 48225 23675 48283 23681
rect 48409 23715 48467 23721
rect 48409 23681 48421 23715
rect 48455 23681 48467 23715
rect 48409 23675 48467 23681
rect 35802 23644 35808 23656
rect 35544 23616 35808 23644
rect 34848 23604 34854 23616
rect 35802 23604 35808 23616
rect 35860 23604 35866 23656
rect 36170 23604 36176 23656
rect 36228 23644 36234 23656
rect 36265 23647 36323 23653
rect 36265 23644 36277 23647
rect 36228 23616 36277 23644
rect 36228 23604 36234 23616
rect 36265 23613 36277 23616
rect 36311 23613 36323 23647
rect 36265 23607 36323 23613
rect 36541 23647 36599 23653
rect 36541 23613 36553 23647
rect 36587 23644 36599 23647
rect 36906 23644 36912 23656
rect 36587 23616 36912 23644
rect 36587 23613 36599 23616
rect 36541 23607 36599 23613
rect 36906 23604 36912 23616
rect 36964 23604 36970 23656
rect 37016 23616 41414 23644
rect 37016 23576 37044 23616
rect 34103 23548 34468 23576
rect 34103 23545 34115 23548
rect 34057 23539 34115 23545
rect 28169 23511 28227 23517
rect 28169 23508 28181 23511
rect 26068 23480 28181 23508
rect 28169 23477 28181 23480
rect 28215 23477 28227 23511
rect 28169 23471 28227 23477
rect 28442 23468 28448 23520
rect 28500 23508 28506 23520
rect 28626 23508 28632 23520
rect 28500 23480 28632 23508
rect 28500 23468 28506 23480
rect 28626 23468 28632 23480
rect 28684 23508 28690 23520
rect 28810 23508 28816 23520
rect 28684 23480 28816 23508
rect 28684 23468 28690 23480
rect 28810 23468 28816 23480
rect 28868 23468 28874 23520
rect 28994 23468 29000 23520
rect 29052 23468 29058 23520
rect 32214 23468 32220 23520
rect 32272 23508 32278 23520
rect 32490 23508 32496 23520
rect 32272 23480 32496 23508
rect 32272 23468 32278 23480
rect 32490 23468 32496 23480
rect 32548 23468 32554 23520
rect 32674 23468 32680 23520
rect 32732 23468 32738 23520
rect 33594 23468 33600 23520
rect 33652 23468 33658 23520
rect 34440 23508 34468 23548
rect 34624 23548 37044 23576
rect 34624 23508 34652 23548
rect 37918 23536 37924 23588
rect 37976 23576 37982 23588
rect 40126 23576 40132 23588
rect 37976 23548 40132 23576
rect 37976 23536 37982 23548
rect 40126 23536 40132 23548
rect 40184 23536 40190 23588
rect 40589 23579 40647 23585
rect 40589 23576 40601 23579
rect 40236 23548 40601 23576
rect 40236 23520 40264 23548
rect 40589 23545 40601 23548
rect 40635 23545 40647 23579
rect 41386 23576 41414 23616
rect 41506 23604 41512 23656
rect 41564 23644 41570 23656
rect 42429 23647 42487 23653
rect 42429 23644 42441 23647
rect 41564 23616 42441 23644
rect 41564 23604 41570 23616
rect 42429 23613 42441 23616
rect 42475 23644 42487 23647
rect 43254 23644 43260 23656
rect 42475 23616 43260 23644
rect 42475 23613 42487 23616
rect 42429 23607 42487 23613
rect 43254 23604 43260 23616
rect 43312 23644 43318 23656
rect 44361 23647 44419 23653
rect 44361 23644 44373 23647
rect 43312 23616 44373 23644
rect 43312 23604 43318 23616
rect 44361 23613 44373 23616
rect 44407 23613 44419 23647
rect 45741 23647 45799 23653
rect 45741 23644 45753 23647
rect 44361 23607 44419 23613
rect 44744 23616 45753 23644
rect 43806 23576 43812 23588
rect 41386 23548 43812 23576
rect 40589 23539 40647 23545
rect 34440 23480 34652 23508
rect 34882 23468 34888 23520
rect 34940 23508 34946 23520
rect 36538 23508 36544 23520
rect 34940 23480 36544 23508
rect 34940 23468 34946 23480
rect 36538 23468 36544 23480
rect 36596 23468 36602 23520
rect 38381 23511 38439 23517
rect 38381 23477 38393 23511
rect 38427 23508 38439 23511
rect 38562 23508 38568 23520
rect 38427 23480 38568 23508
rect 38427 23477 38439 23480
rect 38381 23471 38439 23477
rect 38562 23468 38568 23480
rect 38620 23468 38626 23520
rect 38749 23511 38807 23517
rect 38749 23477 38761 23511
rect 38795 23508 38807 23511
rect 38930 23508 38936 23520
rect 38795 23480 38936 23508
rect 38795 23477 38807 23480
rect 38749 23471 38807 23477
rect 38930 23468 38936 23480
rect 38988 23508 38994 23520
rect 39577 23511 39635 23517
rect 39577 23508 39589 23511
rect 38988 23480 39589 23508
rect 38988 23468 38994 23480
rect 39577 23477 39589 23480
rect 39623 23477 39635 23511
rect 39577 23471 39635 23477
rect 40037 23511 40095 23517
rect 40037 23477 40049 23511
rect 40083 23508 40095 23511
rect 40218 23508 40224 23520
rect 40083 23480 40224 23508
rect 40083 23477 40095 23480
rect 40037 23471 40095 23477
rect 40218 23468 40224 23480
rect 40276 23468 40282 23520
rect 43548 23517 43576 23548
rect 43806 23536 43812 23548
rect 43864 23576 43870 23588
rect 44085 23579 44143 23585
rect 44085 23576 44097 23579
rect 43864 23548 44097 23576
rect 43864 23536 43870 23548
rect 44085 23545 44097 23548
rect 44131 23545 44143 23579
rect 44085 23539 44143 23545
rect 43533 23511 43591 23517
rect 43533 23477 43545 23511
rect 43579 23477 43591 23511
rect 43533 23471 43591 23477
rect 44450 23468 44456 23520
rect 44508 23508 44514 23520
rect 44744 23517 44772 23616
rect 45741 23613 45753 23616
rect 45787 23613 45799 23647
rect 45741 23607 45799 23613
rect 45465 23579 45523 23585
rect 45465 23545 45477 23579
rect 45511 23576 45523 23579
rect 45646 23576 45652 23588
rect 45511 23548 45652 23576
rect 45511 23545 45523 23548
rect 45465 23539 45523 23545
rect 45646 23536 45652 23548
rect 45704 23536 45710 23588
rect 47044 23576 47072 23672
rect 47486 23604 47492 23656
rect 47544 23644 47550 23656
rect 47872 23644 47900 23672
rect 47544 23616 47900 23644
rect 47544 23604 47550 23616
rect 48130 23604 48136 23656
rect 48188 23644 48194 23656
rect 48424 23644 48452 23675
rect 48590 23672 48596 23724
rect 48648 23672 48654 23724
rect 49694 23672 49700 23724
rect 49752 23672 49758 23724
rect 49878 23721 49884 23724
rect 49845 23715 49884 23721
rect 49845 23681 49857 23715
rect 49845 23675 49884 23681
rect 49878 23672 49884 23675
rect 49936 23672 49942 23724
rect 50162 23715 50220 23721
rect 50162 23712 50174 23715
rect 50080 23684 50174 23712
rect 48188 23616 48452 23644
rect 48188 23604 48194 23616
rect 48958 23604 48964 23656
rect 49016 23604 49022 23656
rect 47044 23548 48268 23576
rect 44729 23511 44787 23517
rect 44729 23508 44741 23511
rect 44508 23480 44741 23508
rect 44508 23468 44514 23480
rect 44729 23477 44741 23480
rect 44775 23477 44787 23511
rect 44729 23471 44787 23477
rect 45094 23468 45100 23520
rect 45152 23468 45158 23520
rect 47118 23468 47124 23520
rect 47176 23508 47182 23520
rect 47213 23511 47271 23517
rect 47213 23508 47225 23511
rect 47176 23480 47225 23508
rect 47176 23468 47182 23480
rect 47213 23477 47225 23480
rect 47259 23477 47271 23511
rect 47213 23471 47271 23477
rect 48130 23468 48136 23520
rect 48188 23468 48194 23520
rect 48240 23508 48268 23548
rect 48314 23536 48320 23588
rect 48372 23576 48378 23588
rect 49513 23579 49571 23585
rect 49513 23576 49525 23579
rect 48372 23548 49525 23576
rect 48372 23536 48378 23548
rect 49513 23545 49525 23548
rect 49559 23576 49571 23579
rect 50080 23576 50108 23684
rect 50162 23681 50174 23684
rect 50208 23681 50220 23715
rect 52196 23712 52224 23808
rect 53282 23740 53288 23792
rect 53340 23780 53346 23792
rect 53837 23783 53895 23789
rect 53837 23780 53849 23783
rect 53340 23752 53849 23780
rect 53340 23740 53346 23752
rect 53837 23749 53849 23752
rect 53883 23780 53895 23783
rect 54754 23780 54760 23792
rect 53883 23752 54760 23780
rect 53883 23749 53895 23752
rect 53837 23743 53895 23749
rect 54754 23740 54760 23752
rect 54812 23740 54818 23792
rect 52733 23715 52791 23721
rect 52733 23712 52745 23715
rect 52196 23684 52745 23712
rect 50162 23675 50220 23681
rect 52733 23681 52745 23684
rect 52779 23681 52791 23715
rect 52733 23675 52791 23681
rect 52917 23715 52975 23721
rect 52917 23681 52929 23715
rect 52963 23712 52975 23715
rect 53558 23712 53564 23724
rect 52963 23684 53564 23712
rect 52963 23681 52975 23684
rect 52917 23675 52975 23681
rect 50433 23647 50491 23653
rect 50433 23613 50445 23647
rect 50479 23613 50491 23647
rect 50433 23607 50491 23613
rect 49559 23548 50108 23576
rect 49559 23545 49571 23548
rect 49513 23539 49571 23545
rect 50338 23536 50344 23588
rect 50396 23536 50402 23588
rect 49142 23508 49148 23520
rect 48240 23480 49148 23508
rect 49142 23468 49148 23480
rect 49200 23468 49206 23520
rect 49234 23468 49240 23520
rect 49292 23508 49298 23520
rect 50448 23508 50476 23607
rect 52638 23604 52644 23656
rect 52696 23644 52702 23656
rect 52932 23644 52960 23675
rect 53558 23672 53564 23684
rect 53616 23672 53622 23724
rect 55876 23712 55904 23811
rect 56229 23715 56287 23721
rect 56229 23712 56241 23715
rect 55876 23684 56241 23712
rect 56229 23681 56241 23684
rect 56275 23681 56287 23715
rect 56229 23675 56287 23681
rect 56321 23715 56379 23721
rect 56321 23681 56333 23715
rect 56367 23712 56379 23715
rect 56965 23715 57023 23721
rect 56965 23712 56977 23715
rect 56367 23684 56977 23712
rect 56367 23681 56379 23684
rect 56321 23675 56379 23681
rect 56965 23681 56977 23684
rect 57011 23681 57023 23715
rect 56965 23675 57023 23681
rect 58250 23672 58256 23724
rect 58308 23672 58314 23724
rect 52696 23616 52960 23644
rect 52696 23604 52702 23616
rect 53926 23604 53932 23656
rect 53984 23644 53990 23656
rect 54021 23647 54079 23653
rect 54021 23644 54033 23647
rect 53984 23616 54033 23644
rect 53984 23604 53990 23616
rect 54021 23613 54033 23616
rect 54067 23613 54079 23647
rect 54021 23607 54079 23613
rect 54294 23604 54300 23656
rect 54352 23604 54358 23656
rect 56686 23604 56692 23656
rect 56744 23604 56750 23656
rect 57422 23604 57428 23656
rect 57480 23644 57486 23656
rect 57517 23647 57575 23653
rect 57517 23644 57529 23647
rect 57480 23616 57529 23644
rect 57480 23604 57486 23616
rect 57517 23613 57529 23616
rect 57563 23613 57575 23647
rect 57517 23607 57575 23613
rect 49292 23480 50476 23508
rect 53101 23511 53159 23517
rect 49292 23468 49298 23480
rect 53101 23477 53113 23511
rect 53147 23508 53159 23511
rect 53742 23508 53748 23520
rect 53147 23480 53748 23508
rect 53147 23477 53159 23480
rect 53101 23471 53159 23477
rect 53742 23468 53748 23480
rect 53800 23468 53806 23520
rect 54018 23468 54024 23520
rect 54076 23508 54082 23520
rect 55398 23508 55404 23520
rect 54076 23480 55404 23508
rect 54076 23468 54082 23480
rect 55398 23468 55404 23480
rect 55456 23508 55462 23520
rect 55769 23511 55827 23517
rect 55769 23508 55781 23511
rect 55456 23480 55781 23508
rect 55456 23468 55462 23480
rect 55769 23477 55781 23480
rect 55815 23477 55827 23511
rect 55769 23471 55827 23477
rect 55950 23468 55956 23520
rect 56008 23508 56014 23520
rect 56045 23511 56103 23517
rect 56045 23508 56057 23511
rect 56008 23480 56057 23508
rect 56008 23468 56014 23480
rect 56045 23477 56057 23480
rect 56091 23477 56103 23511
rect 56045 23471 56103 23477
rect 58434 23468 58440 23520
rect 58492 23468 58498 23520
rect 1104 23418 58880 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 58880 23418
rect 1104 23344 58880 23366
rect 20990 23264 20996 23316
rect 21048 23264 21054 23316
rect 22186 23264 22192 23316
rect 22244 23264 22250 23316
rect 22462 23264 22468 23316
rect 22520 23304 22526 23316
rect 23658 23304 23664 23316
rect 22520 23276 23664 23304
rect 22520 23264 22526 23276
rect 23658 23264 23664 23276
rect 23716 23304 23722 23316
rect 23845 23307 23903 23313
rect 23845 23304 23857 23307
rect 23716 23276 23857 23304
rect 23716 23264 23722 23276
rect 23845 23273 23857 23276
rect 23891 23273 23903 23307
rect 23845 23267 23903 23273
rect 22204 23236 22232 23264
rect 21744 23208 22232 23236
rect 19242 23128 19248 23180
rect 19300 23128 19306 23180
rect 21542 23128 21548 23180
rect 21600 23128 21606 23180
rect 17954 23060 17960 23112
rect 18012 23100 18018 23112
rect 21744 23109 21772 23208
rect 22094 23128 22100 23180
rect 22152 23128 22158 23180
rect 22370 23128 22376 23180
rect 22428 23128 22434 23180
rect 18141 23103 18199 23109
rect 18141 23100 18153 23103
rect 18012 23072 18153 23100
rect 18012 23060 18018 23072
rect 18141 23069 18153 23072
rect 18187 23069 18199 23103
rect 21453 23103 21511 23109
rect 21453 23100 21465 23103
rect 18141 23063 18199 23069
rect 20916 23072 21465 23100
rect 18598 22992 18604 23044
rect 18656 23032 18662 23044
rect 19521 23035 19579 23041
rect 19521 23032 19533 23035
rect 18656 23004 19533 23032
rect 18656 22992 18662 23004
rect 19521 23001 19533 23004
rect 19567 23001 19579 23035
rect 19521 22995 19579 23001
rect 19610 22992 19616 23044
rect 19668 23032 19674 23044
rect 19668 23004 20010 23032
rect 19668 22992 19674 23004
rect 19886 22924 19892 22976
rect 19944 22964 19950 22976
rect 20916 22964 20944 23072
rect 21453 23069 21465 23072
rect 21499 23069 21511 23103
rect 21453 23063 21511 23069
rect 21729 23103 21787 23109
rect 21729 23069 21741 23103
rect 21775 23069 21787 23103
rect 21729 23063 21787 23069
rect 21468 23032 21496 23063
rect 21818 23060 21824 23112
rect 21876 23060 21882 23112
rect 23860 23100 23888 23267
rect 28810 23264 28816 23316
rect 28868 23304 28874 23316
rect 29273 23307 29331 23313
rect 29273 23304 29285 23307
rect 28868 23276 29285 23304
rect 28868 23264 28874 23276
rect 29273 23273 29285 23276
rect 29319 23304 29331 23307
rect 30374 23304 30380 23316
rect 29319 23276 30380 23304
rect 29319 23273 29331 23276
rect 29273 23267 29331 23273
rect 30374 23264 30380 23276
rect 30432 23264 30438 23316
rect 34790 23264 34796 23316
rect 34848 23304 34854 23316
rect 34931 23307 34989 23313
rect 34931 23304 34943 23307
rect 34848 23276 34943 23304
rect 34848 23264 34854 23276
rect 34931 23273 34943 23276
rect 34977 23273 34989 23307
rect 34931 23267 34989 23273
rect 35268 23276 38056 23304
rect 26694 23236 26700 23248
rect 25792 23208 26700 23236
rect 25792 23109 25820 23208
rect 26694 23196 26700 23208
rect 26752 23196 26758 23248
rect 32324 23208 33640 23236
rect 28810 23168 28816 23180
rect 26068 23140 28816 23168
rect 26068 23109 26096 23140
rect 28810 23128 28816 23140
rect 28868 23128 28874 23180
rect 31018 23128 31024 23180
rect 31076 23168 31082 23180
rect 32324 23177 32352 23208
rect 32309 23171 32367 23177
rect 32309 23168 32321 23171
rect 31076 23140 32321 23168
rect 31076 23128 31082 23140
rect 32309 23137 32321 23140
rect 32355 23137 32367 23171
rect 32309 23131 32367 23137
rect 32858 23128 32864 23180
rect 32916 23128 32922 23180
rect 25777 23103 25835 23109
rect 25777 23100 25789 23103
rect 23860 23072 25789 23100
rect 25777 23069 25789 23072
rect 25823 23069 25835 23103
rect 25777 23063 25835 23069
rect 26053 23103 26111 23109
rect 26053 23069 26065 23103
rect 26099 23069 26111 23103
rect 26053 23063 26111 23069
rect 26145 23103 26203 23109
rect 26145 23069 26157 23103
rect 26191 23100 26203 23103
rect 26191 23072 27476 23100
rect 26191 23069 26203 23072
rect 26145 23063 26203 23069
rect 21468 23004 22784 23032
rect 19944 22936 20944 22964
rect 22005 22967 22063 22973
rect 19944 22924 19950 22936
rect 22005 22933 22017 22967
rect 22051 22964 22063 22967
rect 22186 22964 22192 22976
rect 22051 22936 22192 22964
rect 22051 22933 22063 22936
rect 22005 22927 22063 22933
rect 22186 22924 22192 22936
rect 22244 22924 22250 22976
rect 22756 22964 22784 23004
rect 22830 22992 22836 23044
rect 22888 22992 22894 23044
rect 24854 22992 24860 23044
rect 24912 23032 24918 23044
rect 25961 23035 26019 23041
rect 25961 23032 25973 23035
rect 24912 23004 25973 23032
rect 24912 22992 24918 23004
rect 25961 23001 25973 23004
rect 26007 23032 26019 23035
rect 26007 23004 26096 23032
rect 26007 23001 26019 23004
rect 25961 22995 26019 23001
rect 26068 22976 26096 23004
rect 23658 22964 23664 22976
rect 22756 22936 23664 22964
rect 23658 22924 23664 22936
rect 23716 22964 23722 22976
rect 24026 22964 24032 22976
rect 23716 22936 24032 22964
rect 23716 22924 23722 22936
rect 24026 22924 24032 22936
rect 24084 22924 24090 22976
rect 26050 22924 26056 22976
rect 26108 22924 26114 22976
rect 26326 22924 26332 22976
rect 26384 22924 26390 22976
rect 27448 22964 27476 23072
rect 27522 23060 27528 23112
rect 27580 23060 27586 23112
rect 31941 23103 31999 23109
rect 31941 23069 31953 23103
rect 31987 23100 31999 23103
rect 32401 23103 32459 23109
rect 32401 23100 32413 23103
rect 31987 23072 32413 23100
rect 31987 23069 31999 23072
rect 31941 23063 31999 23069
rect 32401 23069 32413 23072
rect 32447 23069 32459 23103
rect 32401 23063 32459 23069
rect 32582 23060 32588 23112
rect 32640 23060 32646 23112
rect 32674 23060 32680 23112
rect 32732 23060 32738 23112
rect 32953 23103 33011 23109
rect 32953 23069 32965 23103
rect 32999 23100 33011 23103
rect 33042 23100 33048 23112
rect 32999 23072 33048 23100
rect 32999 23069 33011 23072
rect 32953 23063 33011 23069
rect 27801 23035 27859 23041
rect 27801 23001 27813 23035
rect 27847 23032 27859 23035
rect 28074 23032 28080 23044
rect 27847 23004 28080 23032
rect 27847 23001 27859 23004
rect 27801 22995 27859 23001
rect 28074 22992 28080 23004
rect 28132 22992 28138 23044
rect 28442 22992 28448 23044
rect 28500 22992 28506 23044
rect 31570 22992 31576 23044
rect 31628 22992 31634 23044
rect 32968 23032 32996 23063
rect 33042 23060 33048 23072
rect 33100 23060 33106 23112
rect 33612 23100 33640 23208
rect 33686 23128 33692 23180
rect 33744 23168 33750 23180
rect 35268 23168 35296 23276
rect 33744 23140 35296 23168
rect 33744 23128 33750 23140
rect 35342 23128 35348 23180
rect 35400 23168 35406 23180
rect 36725 23171 36783 23177
rect 36725 23168 36737 23171
rect 35400 23140 36737 23168
rect 35400 23128 35406 23140
rect 36725 23137 36737 23140
rect 36771 23168 36783 23171
rect 37458 23168 37464 23180
rect 36771 23140 37464 23168
rect 36771 23137 36783 23140
rect 36725 23131 36783 23137
rect 37458 23128 37464 23140
rect 37516 23128 37522 23180
rect 35360 23100 35388 23128
rect 33612 23072 35388 23100
rect 36262 23060 36268 23112
rect 36320 23100 36326 23112
rect 36357 23103 36415 23109
rect 36357 23100 36369 23103
rect 36320 23072 36369 23100
rect 36320 23060 36326 23072
rect 36357 23069 36369 23072
rect 36403 23069 36415 23103
rect 36357 23063 36415 23069
rect 36446 23060 36452 23112
rect 36504 23100 36510 23112
rect 36630 23100 36636 23112
rect 36504 23072 36636 23100
rect 36504 23060 36510 23072
rect 36630 23060 36636 23072
rect 36688 23060 36694 23112
rect 38028 23100 38056 23276
rect 39206 23264 39212 23316
rect 39264 23264 39270 23316
rect 39574 23264 39580 23316
rect 39632 23304 39638 23316
rect 39669 23307 39727 23313
rect 39669 23304 39681 23307
rect 39632 23276 39681 23304
rect 39632 23264 39638 23276
rect 39669 23273 39681 23276
rect 39715 23273 39727 23307
rect 39669 23267 39727 23273
rect 40126 23264 40132 23316
rect 40184 23304 40190 23316
rect 40497 23307 40555 23313
rect 40497 23304 40509 23307
rect 40184 23276 40509 23304
rect 40184 23264 40190 23276
rect 40497 23273 40509 23276
rect 40543 23273 40555 23307
rect 40497 23267 40555 23273
rect 40586 23264 40592 23316
rect 40644 23304 40650 23316
rect 41141 23307 41199 23313
rect 41141 23304 41153 23307
rect 40644 23276 41153 23304
rect 40644 23264 40650 23276
rect 41141 23273 41153 23276
rect 41187 23304 41199 23307
rect 41693 23307 41751 23313
rect 41693 23304 41705 23307
rect 41187 23276 41705 23304
rect 41187 23273 41199 23276
rect 41141 23267 41199 23273
rect 41693 23273 41705 23276
rect 41739 23273 41751 23307
rect 41693 23267 41751 23273
rect 43438 23264 43444 23316
rect 43496 23304 43502 23316
rect 43809 23307 43867 23313
rect 43809 23304 43821 23307
rect 43496 23276 43821 23304
rect 43496 23264 43502 23276
rect 43809 23273 43821 23276
rect 43855 23304 43867 23307
rect 44174 23304 44180 23316
rect 43855 23276 44180 23304
rect 43855 23273 43867 23276
rect 43809 23267 43867 23273
rect 44174 23264 44180 23276
rect 44232 23264 44238 23316
rect 44269 23307 44327 23313
rect 44269 23273 44281 23307
rect 44315 23304 44327 23307
rect 44729 23307 44787 23313
rect 44729 23304 44741 23307
rect 44315 23276 44741 23304
rect 44315 23273 44327 23276
rect 44269 23267 44327 23273
rect 44729 23273 44741 23276
rect 44775 23304 44787 23307
rect 45462 23304 45468 23316
rect 44775 23276 45468 23304
rect 44775 23273 44787 23276
rect 44729 23267 44787 23273
rect 45462 23264 45468 23276
rect 45520 23304 45526 23316
rect 45830 23304 45836 23316
rect 45520 23276 45836 23304
rect 45520 23264 45526 23276
rect 45830 23264 45836 23276
rect 45888 23264 45894 23316
rect 46658 23264 46664 23316
rect 46716 23264 46722 23316
rect 47762 23264 47768 23316
rect 47820 23304 47826 23316
rect 48498 23304 48504 23316
rect 47820 23276 48504 23304
rect 47820 23264 47826 23276
rect 48498 23264 48504 23276
rect 48556 23264 48562 23316
rect 49234 23304 49240 23316
rect 48608 23276 49240 23304
rect 38841 23239 38899 23245
rect 38841 23205 38853 23239
rect 38887 23236 38899 23239
rect 38930 23236 38936 23248
rect 38887 23208 38936 23236
rect 38887 23205 38899 23208
rect 38841 23199 38899 23205
rect 38930 23196 38936 23208
rect 38988 23196 38994 23248
rect 41598 23236 41604 23248
rect 39500 23208 41604 23236
rect 38286 23128 38292 23180
rect 38344 23168 38350 23180
rect 38344 23140 39252 23168
rect 38344 23128 38350 23140
rect 38473 23103 38531 23109
rect 38473 23100 38485 23103
rect 38028 23072 38485 23100
rect 38473 23069 38485 23072
rect 38519 23100 38531 23103
rect 39114 23100 39120 23112
rect 38519 23072 39120 23100
rect 38519 23069 38531 23072
rect 38473 23063 38531 23069
rect 39114 23060 39120 23072
rect 39172 23060 39178 23112
rect 32324 23004 32996 23032
rect 32324 22976 32352 23004
rect 35618 22992 35624 23044
rect 35676 22992 35682 23044
rect 39224 23041 39252 23140
rect 39390 23060 39396 23112
rect 39448 23100 39454 23112
rect 39500 23109 39528 23208
rect 41598 23196 41604 23208
rect 41656 23196 41662 23248
rect 41785 23239 41843 23245
rect 41785 23205 41797 23239
rect 41831 23236 41843 23239
rect 43625 23239 43683 23245
rect 43625 23236 43637 23239
rect 41831 23208 43637 23236
rect 41831 23205 41843 23208
rect 41785 23199 41843 23205
rect 43625 23205 43637 23208
rect 43671 23236 43683 23239
rect 46014 23236 46020 23248
rect 43671 23208 46020 23236
rect 43671 23205 43683 23208
rect 43625 23199 43683 23205
rect 46014 23196 46020 23208
rect 46072 23196 46078 23248
rect 39758 23168 39764 23180
rect 39684 23140 39764 23168
rect 39684 23109 39712 23140
rect 39758 23128 39764 23140
rect 39816 23168 39822 23180
rect 39853 23171 39911 23177
rect 39853 23168 39865 23171
rect 39816 23140 39865 23168
rect 39816 23128 39822 23140
rect 39853 23137 39865 23140
rect 39899 23137 39911 23171
rect 39853 23131 39911 23137
rect 40126 23128 40132 23180
rect 40184 23168 40190 23180
rect 41690 23168 41696 23180
rect 40184 23140 41696 23168
rect 40184 23128 40190 23140
rect 41690 23128 41696 23140
rect 41748 23128 41754 23180
rect 42426 23168 42432 23180
rect 41800 23140 42432 23168
rect 39485 23103 39543 23109
rect 39485 23100 39497 23103
rect 39448 23072 39497 23100
rect 39448 23060 39454 23072
rect 39485 23069 39497 23072
rect 39531 23069 39543 23103
rect 39485 23063 39543 23069
rect 39669 23103 39727 23109
rect 39669 23069 39681 23103
rect 39715 23069 39727 23103
rect 39669 23063 39727 23069
rect 39942 23060 39948 23112
rect 40000 23060 40006 23112
rect 41414 23060 41420 23112
rect 41472 23060 41478 23112
rect 41598 23060 41604 23112
rect 41656 23060 41662 23112
rect 39209 23035 39267 23041
rect 39209 23001 39221 23035
rect 39255 23032 39267 23035
rect 41800 23032 41828 23140
rect 42426 23128 42432 23140
rect 42484 23168 42490 23180
rect 42521 23171 42579 23177
rect 42521 23168 42533 23171
rect 42484 23140 42533 23168
rect 42484 23128 42490 23140
rect 42521 23137 42533 23140
rect 42567 23137 42579 23171
rect 42521 23131 42579 23137
rect 44821 23171 44879 23177
rect 44821 23137 44833 23171
rect 44867 23168 44879 23171
rect 45741 23171 45799 23177
rect 45741 23168 45753 23171
rect 44867 23140 45753 23168
rect 44867 23137 44879 23140
rect 44821 23131 44879 23137
rect 45741 23137 45753 23140
rect 45787 23137 45799 23171
rect 47486 23168 47492 23180
rect 45741 23131 45799 23137
rect 46308 23140 47492 23168
rect 46308 23112 46336 23140
rect 47486 23128 47492 23140
rect 47544 23128 47550 23180
rect 48406 23128 48412 23180
rect 48464 23168 48470 23180
rect 48608 23168 48636 23276
rect 49234 23264 49240 23276
rect 49292 23264 49298 23316
rect 49329 23307 49387 23313
rect 49329 23273 49341 23307
rect 49375 23304 49387 23307
rect 49694 23304 49700 23316
rect 49375 23276 49700 23304
rect 49375 23273 49387 23276
rect 49329 23267 49387 23273
rect 49694 23264 49700 23276
rect 49752 23264 49758 23316
rect 49878 23264 49884 23316
rect 49936 23304 49942 23316
rect 49936 23276 50660 23304
rect 49936 23264 49942 23276
rect 50632 23236 50660 23276
rect 50798 23264 50804 23316
rect 50856 23304 50862 23316
rect 50893 23307 50951 23313
rect 50893 23304 50905 23307
rect 50856 23276 50905 23304
rect 50856 23264 50862 23276
rect 50893 23273 50905 23276
rect 50939 23273 50951 23307
rect 50893 23267 50951 23273
rect 53834 23264 53840 23316
rect 53892 23304 53898 23316
rect 54021 23307 54079 23313
rect 54021 23304 54033 23307
rect 53892 23276 54033 23304
rect 53892 23264 53898 23276
rect 54021 23273 54033 23276
rect 54067 23273 54079 23307
rect 54021 23267 54079 23273
rect 52362 23236 52368 23248
rect 50632 23208 52368 23236
rect 48464 23140 48636 23168
rect 48792 23140 50384 23168
rect 48464 23128 48470 23140
rect 41877 23103 41935 23109
rect 41877 23069 41889 23103
rect 41923 23069 41935 23103
rect 41877 23063 41935 23069
rect 42613 23103 42671 23109
rect 42613 23069 42625 23103
rect 42659 23100 42671 23103
rect 42794 23100 42800 23112
rect 42659 23072 42800 23100
rect 42659 23069 42671 23072
rect 42613 23063 42671 23069
rect 39255 23004 41828 23032
rect 39255 23001 39267 23004
rect 39209 22995 39267 23001
rect 27982 22964 27988 22976
rect 27448 22936 27988 22964
rect 27982 22924 27988 22936
rect 28040 22924 28046 22976
rect 30515 22967 30573 22973
rect 30515 22933 30527 22967
rect 30561 22964 30573 22967
rect 32306 22964 32312 22976
rect 30561 22936 32312 22964
rect 30561 22933 30573 22936
rect 30515 22927 30573 22933
rect 32306 22924 32312 22936
rect 32364 22924 32370 22976
rect 33962 22924 33968 22976
rect 34020 22964 34026 22976
rect 36814 22964 36820 22976
rect 34020 22936 36820 22964
rect 34020 22924 34026 22936
rect 36814 22924 36820 22936
rect 36872 22924 36878 22976
rect 38654 22924 38660 22976
rect 38712 22924 38718 22976
rect 39393 22967 39451 22973
rect 39393 22933 39405 22967
rect 39439 22964 39451 22967
rect 39574 22964 39580 22976
rect 39439 22936 39580 22964
rect 39439 22933 39451 22936
rect 39393 22927 39451 22933
rect 39574 22924 39580 22936
rect 39632 22924 39638 22976
rect 39758 22924 39764 22976
rect 39816 22964 39822 22976
rect 41233 22967 41291 22973
rect 41233 22964 41245 22967
rect 39816 22936 41245 22964
rect 39816 22924 39822 22936
rect 41233 22933 41245 22936
rect 41279 22964 41291 22967
rect 41892 22964 41920 23063
rect 42794 23060 42800 23072
rect 42852 23100 42858 23112
rect 43165 23103 43223 23109
rect 43165 23100 43177 23103
rect 42852 23072 43177 23100
rect 42852 23060 42858 23072
rect 43165 23069 43177 23072
rect 43211 23069 43223 23103
rect 43165 23063 43223 23069
rect 43438 23060 43444 23112
rect 43496 23060 43502 23112
rect 45186 23109 45192 23112
rect 44545 23103 44603 23109
rect 44545 23069 44557 23103
rect 44591 23069 44603 23103
rect 45184 23100 45192 23109
rect 45147 23072 45192 23100
rect 44545 23063 44603 23069
rect 45184 23063 45192 23072
rect 42150 22992 42156 23044
rect 42208 22992 42214 23044
rect 42334 22992 42340 23044
rect 42392 23032 42398 23044
rect 43073 23035 43131 23041
rect 43073 23032 43085 23035
rect 42392 23004 43085 23032
rect 42392 22992 42398 23004
rect 43073 23001 43085 23004
rect 43119 23032 43131 23035
rect 44560 23032 44588 23063
rect 45186 23060 45192 23063
rect 45244 23060 45250 23112
rect 45556 23103 45614 23109
rect 45556 23069 45568 23103
rect 45602 23069 45614 23103
rect 45556 23063 45614 23069
rect 43119 23004 43944 23032
rect 44560 23004 45048 23032
rect 43119 23001 43131 23004
rect 43073 22995 43131 23001
rect 43916 22976 43944 23004
rect 41279 22936 41920 22964
rect 41279 22933 41291 22936
rect 41233 22927 41291 22933
rect 42242 22924 42248 22976
rect 42300 22964 42306 22976
rect 43257 22967 43315 22973
rect 43257 22964 43269 22967
rect 42300 22936 43269 22964
rect 42300 22924 42306 22936
rect 43257 22933 43269 22936
rect 43303 22933 43315 22967
rect 43257 22927 43315 22933
rect 43898 22924 43904 22976
rect 43956 22924 43962 22976
rect 44358 22924 44364 22976
rect 44416 22924 44422 22976
rect 45020 22973 45048 23004
rect 45278 22992 45284 23044
rect 45336 22992 45342 23044
rect 45373 23035 45431 23041
rect 45373 23001 45385 23035
rect 45419 23001 45431 23035
rect 45572 23032 45600 23063
rect 45646 23060 45652 23112
rect 45704 23060 45710 23112
rect 46290 23060 46296 23112
rect 46348 23060 46354 23112
rect 48792 23109 48820 23140
rect 48777 23103 48835 23109
rect 48777 23069 48789 23103
rect 48823 23069 48835 23103
rect 48777 23063 48835 23069
rect 49145 23103 49203 23109
rect 49145 23069 49157 23103
rect 49191 23100 49203 23103
rect 49421 23103 49479 23109
rect 49421 23100 49433 23103
rect 49191 23072 49433 23100
rect 49191 23069 49203 23072
rect 49145 23063 49203 23069
rect 49421 23069 49433 23072
rect 49467 23100 49479 23103
rect 49878 23100 49884 23112
rect 49467 23072 49884 23100
rect 49467 23069 49479 23072
rect 49421 23063 49479 23069
rect 49878 23060 49884 23072
rect 49936 23060 49942 23112
rect 50356 23109 50384 23140
rect 50632 23109 50660 23208
rect 52362 23196 52368 23208
rect 52420 23196 52426 23248
rect 50341 23103 50399 23109
rect 50341 23069 50353 23103
rect 50387 23069 50399 23103
rect 50341 23063 50399 23069
rect 50617 23103 50675 23109
rect 50617 23069 50629 23103
rect 50663 23069 50675 23103
rect 50617 23063 50675 23069
rect 46658 23032 46664 23044
rect 45572 23004 46664 23032
rect 45373 22995 45431 23001
rect 45005 22967 45063 22973
rect 45005 22933 45017 22967
rect 45051 22933 45063 22967
rect 45388 22964 45416 22995
rect 46658 22992 46664 23004
rect 46716 22992 46722 23044
rect 47578 22992 47584 23044
rect 47636 22992 47642 23044
rect 48133 23035 48191 23041
rect 48133 23001 48145 23035
rect 48179 23032 48191 23035
rect 48866 23032 48872 23044
rect 48179 23004 48872 23032
rect 48179 23001 48191 23004
rect 48133 22995 48191 23001
rect 48866 22992 48872 23004
rect 48924 22992 48930 23044
rect 48958 22992 48964 23044
rect 49016 22992 49022 23044
rect 49053 23035 49111 23041
rect 49053 23001 49065 23035
rect 49099 23001 49111 23035
rect 49053 22995 49111 23001
rect 45554 22964 45560 22976
rect 45388 22936 45560 22964
rect 45005 22927 45063 22933
rect 45554 22924 45560 22936
rect 45612 22964 45618 22976
rect 46750 22964 46756 22976
rect 45612 22936 46756 22964
rect 45612 22924 45618 22936
rect 46750 22924 46756 22936
rect 46808 22924 46814 22976
rect 47210 22924 47216 22976
rect 47268 22964 47274 22976
rect 48593 22967 48651 22973
rect 48593 22964 48605 22967
rect 47268 22936 48605 22964
rect 47268 22924 47274 22936
rect 48593 22933 48605 22936
rect 48639 22964 48651 22967
rect 49068 22964 49096 22995
rect 48639 22936 49096 22964
rect 50356 22964 50384 23063
rect 50706 23060 50712 23112
rect 50764 23060 50770 23112
rect 53653 23103 53711 23109
rect 53653 23069 53665 23103
rect 53699 23100 53711 23103
rect 53926 23100 53932 23112
rect 53699 23072 53932 23100
rect 53699 23069 53711 23072
rect 53653 23063 53711 23069
rect 50525 23035 50583 23041
rect 50525 23001 50537 23035
rect 50571 23032 50583 23035
rect 50798 23032 50804 23044
rect 50571 23004 50804 23032
rect 50571 23001 50583 23004
rect 50525 22995 50583 23001
rect 50798 22992 50804 23004
rect 50856 22992 50862 23044
rect 52914 22992 52920 23044
rect 52972 22992 52978 23044
rect 53374 22992 53380 23044
rect 53432 22992 53438 23044
rect 53668 23032 53696 23063
rect 53926 23060 53932 23072
rect 53984 23060 53990 23112
rect 54036 23100 54064 23267
rect 57422 23264 57428 23316
rect 57480 23264 57486 23316
rect 55950 23128 55956 23180
rect 56008 23128 56014 23180
rect 54205 23103 54263 23109
rect 54205 23100 54217 23103
rect 54036 23072 54217 23100
rect 54205 23069 54217 23072
rect 54251 23069 54263 23103
rect 55582 23100 55588 23112
rect 54205 23063 54263 23069
rect 54956 23072 55588 23100
rect 53576 23004 53696 23032
rect 53944 23032 53972 23060
rect 54956 23041 54984 23072
rect 55582 23060 55588 23072
rect 55640 23100 55646 23112
rect 55677 23103 55735 23109
rect 55677 23100 55689 23103
rect 55640 23072 55689 23100
rect 55640 23060 55646 23072
rect 55677 23069 55689 23072
rect 55723 23069 55735 23103
rect 55677 23063 55735 23069
rect 54941 23035 54999 23041
rect 54941 23032 54953 23035
rect 53944 23004 54953 23032
rect 51902 22964 51908 22976
rect 50356 22936 51908 22964
rect 48639 22933 48651 22936
rect 48593 22927 48651 22933
rect 51902 22924 51908 22936
rect 51960 22924 51966 22976
rect 52454 22924 52460 22976
rect 52512 22964 52518 22976
rect 53576 22964 53604 23004
rect 54941 23001 54953 23004
rect 54987 23001 54999 23035
rect 54941 22995 54999 23001
rect 55048 23004 56442 23032
rect 52512 22936 53604 22964
rect 52512 22924 52518 22936
rect 53650 22924 53656 22976
rect 53708 22964 53714 22976
rect 55048 22964 55076 23004
rect 53708 22936 55076 22964
rect 56336 22964 56364 23004
rect 56594 22964 56600 22976
rect 56336 22936 56600 22964
rect 53708 22924 53714 22936
rect 56594 22924 56600 22936
rect 56652 22924 56658 22976
rect 1104 22874 58880 22896
rect 1104 22822 4874 22874
rect 4926 22822 4938 22874
rect 4990 22822 5002 22874
rect 5054 22822 5066 22874
rect 5118 22822 5130 22874
rect 5182 22822 35594 22874
rect 35646 22822 35658 22874
rect 35710 22822 35722 22874
rect 35774 22822 35786 22874
rect 35838 22822 35850 22874
rect 35902 22822 58880 22874
rect 1104 22800 58880 22822
rect 19429 22763 19487 22769
rect 19429 22729 19441 22763
rect 19475 22760 19487 22763
rect 22002 22760 22008 22772
rect 19475 22732 22008 22760
rect 19475 22729 19487 22732
rect 19429 22723 19487 22729
rect 17954 22652 17960 22704
rect 18012 22692 18018 22704
rect 19061 22695 19119 22701
rect 19061 22692 19073 22695
rect 18012 22664 19073 22692
rect 18012 22652 18018 22664
rect 19061 22661 19073 22664
rect 19107 22692 19119 22695
rect 19242 22692 19248 22704
rect 19107 22664 19248 22692
rect 19107 22661 19119 22664
rect 19061 22655 19119 22661
rect 19242 22652 19248 22664
rect 19300 22652 19306 22704
rect 18322 22584 18328 22636
rect 18380 22624 18386 22636
rect 19444 22624 19472 22723
rect 22002 22720 22008 22732
rect 22060 22720 22066 22772
rect 22830 22760 22836 22772
rect 22480 22732 22836 22760
rect 22094 22692 22100 22704
rect 21836 22664 22100 22692
rect 19794 22633 19800 22636
rect 19792 22624 19800 22633
rect 18380 22596 19472 22624
rect 19755 22596 19800 22624
rect 18380 22584 18386 22596
rect 19792 22587 19800 22596
rect 19794 22584 19800 22587
rect 19852 22584 19858 22636
rect 19886 22584 19892 22636
rect 19944 22584 19950 22636
rect 19978 22584 19984 22636
rect 20036 22584 20042 22636
rect 20070 22584 20076 22636
rect 20128 22633 20134 22636
rect 21836 22633 21864 22664
rect 22094 22652 22100 22664
rect 22152 22652 22158 22704
rect 22480 22692 22508 22732
rect 22830 22720 22836 22732
rect 22888 22720 22894 22772
rect 23569 22763 23627 22769
rect 23569 22729 23581 22763
rect 23615 22760 23627 22763
rect 23658 22760 23664 22772
rect 23615 22732 23664 22760
rect 23615 22729 23627 22732
rect 23569 22723 23627 22729
rect 23658 22720 23664 22732
rect 23716 22720 23722 22772
rect 27430 22760 27436 22772
rect 25792 22732 27436 22760
rect 22554 22692 22560 22704
rect 22480 22664 22560 22692
rect 22554 22652 22560 22664
rect 22612 22652 22618 22704
rect 20128 22627 20167 22633
rect 20155 22593 20167 22627
rect 20128 22587 20167 22593
rect 20257 22627 20315 22633
rect 20257 22593 20269 22627
rect 20303 22624 20315 22627
rect 21821 22627 21879 22633
rect 20303 22596 20484 22624
rect 20303 22593 20315 22596
rect 20257 22587 20315 22593
rect 20128 22584 20134 22587
rect 19812 22556 19840 22584
rect 20346 22556 20352 22568
rect 19812 22528 20352 22556
rect 20346 22516 20352 22528
rect 20404 22516 20410 22568
rect 20456 22432 20484 22596
rect 21821 22593 21833 22627
rect 21867 22593 21879 22627
rect 21821 22587 21879 22593
rect 23750 22584 23756 22636
rect 23808 22624 23814 22636
rect 25590 22624 25596 22636
rect 23808 22596 25596 22624
rect 23808 22584 23814 22596
rect 25590 22584 25596 22596
rect 25648 22624 25654 22636
rect 25792 22633 25820 22732
rect 27430 22720 27436 22732
rect 27488 22720 27494 22772
rect 28074 22720 28080 22772
rect 28132 22720 28138 22772
rect 34606 22720 34612 22772
rect 34664 22760 34670 22772
rect 34664 22732 35848 22760
rect 34664 22720 34670 22732
rect 35820 22704 35848 22732
rect 35986 22720 35992 22772
rect 36044 22720 36050 22772
rect 36173 22763 36231 22769
rect 36173 22729 36185 22763
rect 36219 22760 36231 22763
rect 36219 22732 36584 22760
rect 36219 22729 36231 22732
rect 36173 22723 36231 22729
rect 26326 22692 26332 22704
rect 26068 22664 26332 22692
rect 26068 22633 26096 22664
rect 26326 22652 26332 22664
rect 26384 22652 26390 22704
rect 28534 22692 28540 22704
rect 28276 22664 28540 22692
rect 28276 22636 28304 22664
rect 28534 22652 28540 22664
rect 28592 22692 28598 22704
rect 28721 22695 28779 22701
rect 28721 22692 28733 22695
rect 28592 22664 28733 22692
rect 28592 22652 28598 22664
rect 28721 22661 28733 22664
rect 28767 22661 28779 22695
rect 28721 22655 28779 22661
rect 32122 22652 32128 22704
rect 32180 22692 32186 22704
rect 32180 22664 32720 22692
rect 32180 22652 32186 22664
rect 32692 22636 32720 22664
rect 34790 22652 34796 22704
rect 34848 22692 34854 22704
rect 34848 22664 35664 22692
rect 34848 22652 34854 22664
rect 25777 22627 25835 22633
rect 25777 22624 25789 22627
rect 25648 22596 25789 22624
rect 25648 22584 25654 22596
rect 25777 22593 25789 22596
rect 25823 22593 25835 22627
rect 25777 22587 25835 22593
rect 26053 22627 26111 22633
rect 26053 22593 26065 22627
rect 26099 22593 26111 22627
rect 26053 22587 26111 22593
rect 26145 22627 26203 22633
rect 26145 22593 26157 22627
rect 26191 22624 26203 22627
rect 26970 22624 26976 22636
rect 26191 22596 26976 22624
rect 26191 22593 26203 22596
rect 26145 22587 26203 22593
rect 22097 22559 22155 22565
rect 22097 22525 22109 22559
rect 22143 22556 22155 22559
rect 22186 22556 22192 22568
rect 22143 22528 22192 22556
rect 22143 22525 22155 22528
rect 22097 22519 22155 22525
rect 22186 22516 22192 22528
rect 22244 22516 22250 22568
rect 26160 22556 26188 22587
rect 26970 22584 26976 22596
rect 27028 22584 27034 22636
rect 28258 22584 28264 22636
rect 28316 22584 28322 22636
rect 28350 22584 28356 22636
rect 28408 22584 28414 22636
rect 28442 22584 28448 22636
rect 28500 22624 28506 22636
rect 28629 22627 28687 22633
rect 28629 22624 28641 22627
rect 28500 22596 28641 22624
rect 28500 22584 28506 22596
rect 28629 22593 28641 22596
rect 28675 22624 28687 22627
rect 28810 22624 28816 22636
rect 28675 22596 28816 22624
rect 28675 22593 28687 22596
rect 28629 22587 28687 22593
rect 28810 22584 28816 22596
rect 28868 22584 28874 22636
rect 32309 22627 32367 22633
rect 32309 22593 32321 22627
rect 32355 22593 32367 22627
rect 32309 22587 32367 22593
rect 25792 22528 26188 22556
rect 19610 22380 19616 22432
rect 19668 22380 19674 22432
rect 20438 22380 20444 22432
rect 20496 22380 20502 22432
rect 21818 22380 21824 22432
rect 21876 22420 21882 22432
rect 25792 22420 25820 22528
rect 31570 22516 31576 22568
rect 31628 22556 31634 22568
rect 32324 22556 32352 22587
rect 32398 22584 32404 22636
rect 32456 22584 32462 22636
rect 32674 22584 32680 22636
rect 32732 22584 32738 22636
rect 32769 22627 32827 22633
rect 32769 22593 32781 22627
rect 32815 22624 32827 22627
rect 34698 22624 34704 22636
rect 32815 22596 34704 22624
rect 32815 22593 32827 22596
rect 32769 22587 32827 22593
rect 34698 22584 34704 22596
rect 34756 22584 34762 22636
rect 35161 22627 35219 22633
rect 35161 22593 35173 22627
rect 35207 22624 35219 22627
rect 35207 22596 35241 22624
rect 35207 22593 35219 22596
rect 35161 22587 35219 22593
rect 33226 22556 33232 22568
rect 31628 22528 33232 22556
rect 31628 22516 31634 22528
rect 33226 22516 33232 22528
rect 33284 22516 33290 22568
rect 25866 22448 25872 22500
rect 25924 22488 25930 22500
rect 26234 22488 26240 22500
rect 25924 22460 26240 22488
rect 25924 22448 25930 22460
rect 26234 22448 26240 22460
rect 26292 22448 26298 22500
rect 28537 22491 28595 22497
rect 28537 22457 28549 22491
rect 28583 22488 28595 22491
rect 30006 22488 30012 22500
rect 28583 22460 30012 22488
rect 28583 22457 28595 22460
rect 28537 22451 28595 22457
rect 30006 22448 30012 22460
rect 30064 22448 30070 22500
rect 32766 22448 32772 22500
rect 32824 22488 32830 22500
rect 34422 22488 34428 22500
rect 32824 22460 34428 22488
rect 32824 22448 32830 22460
rect 34422 22448 34428 22460
rect 34480 22448 34486 22500
rect 34716 22488 34744 22584
rect 34977 22559 35035 22565
rect 34977 22525 34989 22559
rect 35023 22556 35035 22559
rect 35176 22556 35204 22587
rect 35342 22584 35348 22636
rect 35400 22624 35406 22636
rect 35636 22633 35664 22664
rect 35802 22652 35808 22704
rect 35860 22652 35866 22704
rect 35897 22695 35955 22701
rect 35897 22661 35909 22695
rect 35943 22692 35955 22695
rect 36004 22692 36032 22720
rect 35943 22664 36032 22692
rect 35943 22661 35955 22664
rect 35897 22655 35955 22661
rect 35529 22627 35587 22633
rect 35529 22624 35541 22627
rect 35400 22596 35541 22624
rect 35400 22584 35406 22596
rect 35529 22593 35541 22596
rect 35575 22593 35587 22627
rect 35529 22587 35587 22593
rect 35621 22627 35679 22633
rect 35621 22593 35633 22627
rect 35667 22593 35679 22627
rect 35621 22587 35679 22593
rect 35989 22627 36047 22633
rect 35989 22593 36001 22627
rect 36035 22624 36047 22627
rect 36078 22624 36084 22636
rect 36035 22596 36084 22624
rect 36035 22593 36047 22596
rect 35989 22587 36047 22593
rect 35894 22556 35900 22568
rect 35023 22528 35900 22556
rect 35023 22525 35035 22528
rect 34977 22519 35035 22525
rect 35894 22516 35900 22528
rect 35952 22516 35958 22568
rect 36004 22488 36032 22587
rect 36078 22584 36084 22596
rect 36136 22584 36142 22636
rect 36265 22627 36323 22633
rect 36265 22593 36277 22627
rect 36311 22624 36323 22627
rect 36446 22624 36452 22636
rect 36311 22596 36452 22624
rect 36311 22593 36323 22596
rect 36265 22587 36323 22593
rect 36446 22584 36452 22596
rect 36504 22584 36510 22636
rect 36556 22633 36584 22732
rect 37826 22720 37832 22772
rect 37884 22720 37890 22772
rect 38654 22720 38660 22772
rect 38712 22760 38718 22772
rect 38841 22763 38899 22769
rect 38841 22760 38853 22763
rect 38712 22732 38853 22760
rect 38712 22720 38718 22732
rect 38841 22729 38853 22732
rect 38887 22729 38899 22763
rect 38841 22723 38899 22729
rect 39390 22720 39396 22772
rect 39448 22720 39454 22772
rect 42334 22760 42340 22772
rect 39500 22732 42340 22760
rect 36541 22627 36599 22633
rect 36541 22593 36553 22627
rect 36587 22593 36599 22627
rect 36541 22587 36599 22593
rect 36630 22584 36636 22636
rect 36688 22584 36694 22636
rect 37550 22584 37556 22636
rect 37608 22624 37614 22636
rect 37844 22624 37872 22720
rect 38289 22695 38347 22701
rect 38289 22661 38301 22695
rect 38335 22692 38347 22695
rect 39408 22692 39436 22720
rect 38335 22664 39436 22692
rect 38335 22661 38347 22664
rect 38289 22655 38347 22661
rect 38105 22627 38163 22633
rect 38105 22624 38117 22627
rect 37608 22596 38117 22624
rect 37608 22584 37614 22596
rect 38105 22593 38117 22596
rect 38151 22593 38163 22627
rect 38105 22587 38163 22593
rect 38378 22584 38384 22636
rect 38436 22584 38442 22636
rect 39114 22584 39120 22636
rect 39172 22624 39178 22636
rect 39301 22627 39359 22633
rect 39301 22624 39313 22627
rect 39172 22596 39313 22624
rect 39172 22584 39178 22596
rect 39301 22593 39313 22596
rect 39347 22593 39359 22627
rect 39301 22587 39359 22593
rect 36354 22516 36360 22568
rect 36412 22516 36418 22568
rect 36648 22488 36676 22584
rect 36814 22516 36820 22568
rect 36872 22556 36878 22568
rect 39500 22556 39528 22732
rect 42334 22720 42340 22732
rect 42392 22720 42398 22772
rect 42429 22763 42487 22769
rect 42429 22729 42441 22763
rect 42475 22729 42487 22763
rect 42429 22723 42487 22729
rect 42444 22692 42472 22723
rect 42702 22720 42708 22772
rect 42760 22760 42766 22772
rect 42760 22732 44496 22760
rect 42760 22720 42766 22732
rect 41432 22664 42472 22692
rect 42797 22695 42855 22701
rect 39574 22584 39580 22636
rect 39632 22624 39638 22636
rect 39942 22624 39948 22636
rect 39632 22596 39948 22624
rect 39632 22584 39638 22596
rect 39942 22584 39948 22596
rect 40000 22584 40006 22636
rect 41432 22633 41460 22664
rect 42797 22661 42809 22695
rect 42843 22692 42855 22695
rect 43530 22692 43536 22704
rect 42843 22664 43536 22692
rect 42843 22661 42855 22664
rect 42797 22655 42855 22661
rect 43530 22652 43536 22664
rect 43588 22652 43594 22704
rect 44358 22652 44364 22704
rect 44416 22652 44422 22704
rect 44468 22692 44496 22732
rect 48866 22720 48872 22772
rect 48924 22720 48930 22772
rect 49050 22720 49056 22772
rect 49108 22760 49114 22772
rect 49605 22763 49663 22769
rect 49605 22760 49617 22763
rect 49108 22732 49617 22760
rect 49108 22720 49114 22732
rect 49605 22729 49617 22732
rect 49651 22760 49663 22763
rect 49694 22760 49700 22772
rect 49651 22732 49700 22760
rect 49651 22729 49663 22732
rect 49605 22723 49663 22729
rect 49694 22720 49700 22732
rect 49752 22760 49758 22772
rect 53282 22760 53288 22772
rect 49752 22732 53288 22760
rect 49752 22720 49758 22732
rect 53282 22720 53288 22732
rect 53340 22720 53346 22772
rect 53374 22720 53380 22772
rect 53432 22760 53438 22772
rect 54021 22763 54079 22769
rect 54021 22760 54033 22763
rect 53432 22732 54033 22760
rect 53432 22720 53438 22732
rect 54021 22729 54033 22732
rect 54067 22729 54079 22763
rect 54021 22723 54079 22729
rect 44468 22664 44850 22692
rect 48130 22652 48136 22704
rect 48188 22692 48194 22704
rect 48188 22664 48636 22692
rect 48188 22652 48194 22664
rect 41325 22627 41383 22633
rect 41325 22593 41337 22627
rect 41371 22593 41383 22627
rect 41325 22587 41383 22593
rect 41417 22627 41475 22633
rect 41417 22593 41429 22627
rect 41463 22593 41475 22627
rect 41417 22587 41475 22593
rect 36872 22528 39528 22556
rect 41340 22556 41368 22587
rect 41598 22584 41604 22636
rect 41656 22624 41662 22636
rect 41693 22627 41751 22633
rect 41693 22624 41705 22627
rect 41656 22596 41705 22624
rect 41656 22584 41662 22596
rect 41693 22593 41705 22596
rect 41739 22624 41751 22627
rect 41785 22627 41843 22633
rect 41785 22624 41797 22627
rect 41739 22596 41797 22624
rect 41739 22593 41751 22596
rect 41693 22587 41751 22593
rect 41785 22593 41797 22596
rect 41831 22624 41843 22627
rect 42242 22624 42248 22636
rect 41831 22596 42248 22624
rect 41831 22593 41843 22596
rect 41785 22587 41843 22593
rect 42242 22584 42248 22596
rect 42300 22584 42306 22636
rect 42610 22584 42616 22636
rect 42668 22584 42674 22636
rect 42705 22627 42763 22633
rect 42705 22593 42717 22627
rect 42751 22593 42763 22627
rect 42705 22587 42763 22593
rect 41506 22556 41512 22568
rect 41340 22528 41512 22556
rect 36872 22516 36878 22528
rect 41506 22516 41512 22528
rect 41564 22516 41570 22568
rect 42518 22516 42524 22568
rect 42576 22556 42582 22568
rect 42720 22556 42748 22587
rect 42978 22584 42984 22636
rect 43036 22584 43042 22636
rect 46658 22584 46664 22636
rect 46716 22624 46722 22636
rect 48608 22633 48636 22664
rect 53650 22652 53656 22704
rect 53708 22692 53714 22704
rect 53708 22664 54694 22692
rect 53708 22652 53714 22664
rect 55582 22652 55588 22704
rect 55640 22692 55646 22704
rect 55640 22664 56180 22692
rect 55640 22652 55646 22664
rect 56152 22636 56180 22664
rect 47581 22627 47639 22633
rect 47581 22624 47593 22627
rect 46716 22596 47593 22624
rect 46716 22584 46722 22596
rect 47581 22593 47593 22596
rect 47627 22593 47639 22627
rect 47581 22587 47639 22593
rect 48225 22627 48283 22633
rect 48225 22593 48237 22627
rect 48271 22624 48283 22627
rect 48317 22627 48375 22633
rect 48317 22624 48329 22627
rect 48271 22596 48329 22624
rect 48271 22593 48283 22596
rect 48225 22587 48283 22593
rect 48317 22593 48329 22596
rect 48363 22593 48375 22627
rect 48317 22587 48375 22593
rect 48593 22627 48651 22633
rect 48593 22593 48605 22627
rect 48639 22593 48651 22627
rect 48593 22587 48651 22593
rect 48685 22627 48743 22633
rect 48685 22593 48697 22627
rect 48731 22593 48743 22627
rect 48685 22587 48743 22593
rect 42576 22528 43208 22556
rect 42576 22516 42582 22528
rect 43180 22497 43208 22528
rect 43990 22516 43996 22568
rect 44048 22556 44054 22568
rect 44085 22559 44143 22565
rect 44085 22556 44097 22559
rect 44048 22528 44097 22556
rect 44048 22516 44054 22528
rect 44085 22525 44097 22528
rect 44131 22525 44143 22559
rect 47210 22556 47216 22568
rect 44085 22519 44143 22525
rect 44192 22528 47216 22556
rect 34716 22460 36032 22488
rect 36096 22460 36676 22488
rect 41049 22491 41107 22497
rect 21876 22392 25820 22420
rect 21876 22380 21882 22392
rect 26326 22380 26332 22432
rect 26384 22380 26390 22432
rect 32122 22380 32128 22432
rect 32180 22380 32186 22432
rect 32585 22423 32643 22429
rect 32585 22389 32597 22423
rect 32631 22420 32643 22423
rect 32858 22420 32864 22432
rect 32631 22392 32864 22420
rect 32631 22389 32643 22392
rect 32585 22383 32643 22389
rect 32858 22380 32864 22392
rect 32916 22380 32922 22432
rect 32953 22423 33011 22429
rect 32953 22389 32965 22423
rect 32999 22420 33011 22423
rect 33134 22420 33140 22432
rect 32999 22392 33140 22420
rect 32999 22389 33011 22392
rect 32953 22383 33011 22389
rect 33134 22380 33140 22392
rect 33192 22420 33198 22432
rect 33594 22420 33600 22432
rect 33192 22392 33600 22420
rect 33192 22380 33198 22392
rect 33594 22380 33600 22392
rect 33652 22380 33658 22432
rect 35342 22380 35348 22432
rect 35400 22420 35406 22432
rect 36096 22420 36124 22460
rect 41049 22457 41061 22491
rect 41095 22488 41107 22491
rect 43165 22491 43223 22497
rect 41095 22460 41644 22488
rect 41095 22457 41107 22460
rect 41049 22451 41107 22457
rect 35400 22392 36124 22420
rect 36817 22423 36875 22429
rect 35400 22380 35406 22392
rect 36817 22389 36829 22423
rect 36863 22420 36875 22423
rect 37642 22420 37648 22432
rect 36863 22392 37648 22420
rect 36863 22389 36875 22392
rect 36817 22383 36875 22389
rect 37642 22380 37648 22392
rect 37700 22380 37706 22432
rect 37826 22380 37832 22432
rect 37884 22420 37890 22432
rect 37921 22423 37979 22429
rect 37921 22420 37933 22423
rect 37884 22392 37933 22420
rect 37884 22380 37890 22392
rect 37921 22389 37933 22392
rect 37967 22389 37979 22423
rect 37921 22383 37979 22389
rect 39758 22380 39764 22432
rect 39816 22420 39822 22432
rect 39853 22423 39911 22429
rect 39853 22420 39865 22423
rect 39816 22392 39865 22420
rect 39816 22380 39822 22392
rect 39853 22389 39865 22392
rect 39899 22389 39911 22423
rect 39853 22383 39911 22389
rect 41138 22380 41144 22432
rect 41196 22380 41202 22432
rect 41616 22429 41644 22460
rect 43165 22457 43177 22491
rect 43211 22488 43223 22491
rect 44192 22488 44220 22528
rect 47210 22516 47216 22528
rect 47268 22516 47274 22568
rect 47397 22559 47455 22565
rect 47397 22525 47409 22559
rect 47443 22556 47455 22559
rect 47670 22556 47676 22568
rect 47443 22528 47676 22556
rect 47443 22525 47455 22528
rect 47397 22519 47455 22525
rect 47670 22516 47676 22528
rect 47728 22556 47734 22568
rect 48700 22556 48728 22587
rect 49234 22584 49240 22636
rect 49292 22624 49298 22636
rect 49329 22627 49387 22633
rect 49329 22624 49341 22627
rect 49292 22596 49341 22624
rect 49292 22584 49298 22596
rect 49329 22593 49341 22596
rect 49375 22593 49387 22627
rect 49329 22587 49387 22593
rect 51902 22584 51908 22636
rect 51960 22624 51966 22636
rect 52733 22627 52791 22633
rect 52733 22624 52745 22627
rect 51960 22596 52745 22624
rect 51960 22584 51966 22596
rect 52733 22593 52745 22596
rect 52779 22593 52791 22627
rect 52733 22587 52791 22593
rect 53377 22627 53435 22633
rect 53377 22593 53389 22627
rect 53423 22624 53435 22627
rect 53469 22627 53527 22633
rect 53469 22624 53481 22627
rect 53423 22596 53481 22624
rect 53423 22593 53435 22596
rect 53377 22587 53435 22593
rect 53469 22593 53481 22596
rect 53515 22593 53527 22627
rect 53469 22587 53527 22593
rect 53742 22584 53748 22636
rect 53800 22584 53806 22636
rect 53837 22627 53895 22633
rect 53837 22593 53849 22627
rect 53883 22593 53895 22627
rect 53837 22587 53895 22593
rect 53852 22556 53880 22587
rect 56134 22584 56140 22636
rect 56192 22584 56198 22636
rect 58250 22584 58256 22636
rect 58308 22584 58314 22636
rect 54113 22559 54171 22565
rect 54113 22556 54125 22559
rect 47728 22528 54125 22556
rect 47728 22516 47734 22528
rect 54113 22525 54125 22528
rect 54159 22525 54171 22559
rect 54113 22519 54171 22525
rect 55858 22516 55864 22568
rect 55916 22516 55922 22568
rect 50982 22488 50988 22500
rect 43211 22460 44220 22488
rect 48424 22460 50988 22488
rect 43211 22457 43223 22460
rect 43165 22451 43223 22457
rect 41601 22423 41659 22429
rect 41601 22389 41613 22423
rect 41647 22420 41659 22423
rect 42150 22420 42156 22432
rect 41647 22392 42156 22420
rect 41647 22389 41659 22392
rect 41601 22383 41659 22389
rect 42150 22380 42156 22392
rect 42208 22380 42214 22432
rect 42978 22380 42984 22432
rect 43036 22420 43042 22432
rect 45833 22423 45891 22429
rect 45833 22420 45845 22423
rect 43036 22392 45845 22420
rect 43036 22380 43042 22392
rect 45833 22389 45845 22392
rect 45879 22420 45891 22423
rect 46290 22420 46296 22432
rect 45879 22392 46296 22420
rect 45879 22389 45891 22392
rect 45833 22383 45891 22389
rect 46290 22380 46296 22392
rect 46348 22380 46354 22432
rect 48038 22380 48044 22432
rect 48096 22420 48102 22432
rect 48424 22429 48452 22460
rect 50982 22448 50988 22460
rect 51040 22448 51046 22500
rect 58434 22448 58440 22500
rect 58492 22448 58498 22500
rect 48409 22423 48467 22429
rect 48409 22420 48421 22423
rect 48096 22392 48421 22420
rect 48096 22380 48102 22392
rect 48409 22389 48421 22392
rect 48455 22389 48467 22423
rect 48409 22383 48467 22389
rect 48682 22380 48688 22432
rect 48740 22420 48746 22432
rect 48866 22420 48872 22432
rect 48740 22392 48872 22420
rect 48740 22380 48746 22392
rect 48866 22380 48872 22392
rect 48924 22380 48930 22432
rect 53558 22380 53564 22432
rect 53616 22380 53622 22432
rect 54386 22380 54392 22432
rect 54444 22380 54450 22432
rect 1104 22330 58880 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 58880 22330
rect 1104 22256 58880 22278
rect 18598 22176 18604 22228
rect 18656 22176 18662 22228
rect 20438 22176 20444 22228
rect 20496 22216 20502 22228
rect 22738 22216 22744 22228
rect 20496 22188 22744 22216
rect 20496 22176 20502 22188
rect 22738 22176 22744 22188
rect 22796 22216 22802 22228
rect 24854 22216 24860 22228
rect 22796 22188 24860 22216
rect 22796 22176 22802 22188
rect 24854 22176 24860 22188
rect 24912 22176 24918 22228
rect 25590 22176 25596 22228
rect 25648 22176 25654 22228
rect 25866 22176 25872 22228
rect 25924 22176 25930 22228
rect 26326 22176 26332 22228
rect 26384 22216 26390 22228
rect 27077 22219 27135 22225
rect 27077 22216 27089 22219
rect 26384 22188 27089 22216
rect 26384 22176 26390 22188
rect 27077 22185 27089 22188
rect 27123 22185 27135 22219
rect 27077 22179 27135 22185
rect 28166 22176 28172 22228
rect 28224 22216 28230 22228
rect 28994 22216 29000 22228
rect 28224 22188 29000 22216
rect 28224 22176 28230 22188
rect 28994 22176 29000 22188
rect 29052 22216 29058 22228
rect 30282 22216 30288 22228
rect 29052 22188 30288 22216
rect 29052 22176 29058 22188
rect 30282 22176 30288 22188
rect 30340 22176 30346 22228
rect 32674 22176 32680 22228
rect 32732 22216 32738 22228
rect 32999 22219 33057 22225
rect 32999 22216 33011 22219
rect 32732 22188 33011 22216
rect 32732 22176 32738 22188
rect 32999 22185 33011 22188
rect 33045 22185 33057 22219
rect 32999 22179 33057 22185
rect 25884 22148 25912 22176
rect 25792 22120 25912 22148
rect 19610 22080 19616 22092
rect 18800 22052 19616 22080
rect 18800 22021 18828 22052
rect 19610 22040 19616 22052
rect 19668 22040 19674 22092
rect 20990 22080 20996 22092
rect 19812 22052 20996 22080
rect 18785 22015 18843 22021
rect 18785 21981 18797 22015
rect 18831 21981 18843 22015
rect 18785 21975 18843 21981
rect 18969 22015 19027 22021
rect 18969 21981 18981 22015
rect 19015 21981 19027 22015
rect 18969 21975 19027 21981
rect 19061 22015 19119 22021
rect 19061 21981 19073 22015
rect 19107 22012 19119 22015
rect 19812 22012 19840 22052
rect 20990 22040 20996 22052
rect 21048 22040 21054 22092
rect 19107 21984 19840 22012
rect 19107 21981 19119 21984
rect 19061 21975 19119 21981
rect 18984 21944 19012 21975
rect 19886 21972 19892 22024
rect 19944 21972 19950 22024
rect 23569 22015 23627 22021
rect 23569 21981 23581 22015
rect 23615 22012 23627 22015
rect 25792 22012 25820 22120
rect 27982 22108 27988 22160
rect 28040 22148 28046 22160
rect 28040 22120 29408 22148
rect 28040 22108 28046 22120
rect 27341 22083 27399 22089
rect 27341 22049 27353 22083
rect 27387 22080 27399 22083
rect 27522 22080 27528 22092
rect 27387 22052 27528 22080
rect 27387 22049 27399 22052
rect 27341 22043 27399 22049
rect 27522 22040 27528 22052
rect 27580 22040 27586 22092
rect 29086 22040 29092 22092
rect 29144 22080 29150 22092
rect 29380 22080 29408 22120
rect 29144 22052 29408 22080
rect 29144 22040 29150 22052
rect 27893 22015 27951 22021
rect 27893 22012 27905 22015
rect 23615 21984 25820 22012
rect 27356 21984 27905 22012
rect 23615 21981 23627 21984
rect 23569 21975 23627 21981
rect 19334 21944 19340 21956
rect 18984 21916 19340 21944
rect 19334 21904 19340 21916
rect 19392 21904 19398 21956
rect 19797 21947 19855 21953
rect 19797 21913 19809 21947
rect 19843 21944 19855 21947
rect 19904 21944 19932 21972
rect 20530 21944 20536 21956
rect 19843 21916 19932 21944
rect 19996 21916 20536 21944
rect 19843 21913 19855 21916
rect 19797 21907 19855 21913
rect 19426 21836 19432 21888
rect 19484 21876 19490 21888
rect 19996 21876 20024 21916
rect 20530 21904 20536 21916
rect 20588 21904 20594 21956
rect 20898 21904 20904 21956
rect 20956 21944 20962 21956
rect 24210 21944 24216 21956
rect 20956 21916 24216 21944
rect 20956 21904 20962 21916
rect 24210 21904 24216 21916
rect 24268 21904 24274 21956
rect 27356 21944 27384 21984
rect 27893 21981 27905 21984
rect 27939 22012 27951 22015
rect 28534 22012 28540 22024
rect 27939 21984 28540 22012
rect 27939 21981 27951 21984
rect 27893 21975 27951 21981
rect 28534 21972 28540 21984
rect 28592 21972 28598 22024
rect 29380 22012 29408 22052
rect 31573 22083 31631 22089
rect 31573 22049 31585 22083
rect 31619 22080 31631 22083
rect 32122 22080 32128 22092
rect 31619 22052 32128 22080
rect 31619 22049 31631 22052
rect 31573 22043 31631 22049
rect 32122 22040 32128 22052
rect 32180 22040 32186 22092
rect 33014 22080 33042 22179
rect 34422 22176 34428 22228
rect 34480 22216 34486 22228
rect 35618 22216 35624 22228
rect 34480 22188 35624 22216
rect 34480 22176 34486 22188
rect 35618 22176 35624 22188
rect 35676 22176 35682 22228
rect 35710 22176 35716 22228
rect 35768 22216 35774 22228
rect 35986 22216 35992 22228
rect 35768 22188 35992 22216
rect 35768 22176 35774 22188
rect 35986 22176 35992 22188
rect 36044 22176 36050 22228
rect 36262 22225 36268 22228
rect 36219 22219 36268 22225
rect 36219 22185 36231 22219
rect 36265 22185 36268 22219
rect 36219 22179 36268 22185
rect 36262 22176 36268 22179
rect 36320 22216 36326 22228
rect 36446 22216 36452 22228
rect 36320 22188 36452 22216
rect 36320 22176 36326 22188
rect 36446 22176 36452 22188
rect 36504 22176 36510 22228
rect 40668 22219 40726 22225
rect 40668 22185 40680 22219
rect 40714 22216 40726 22219
rect 41138 22216 41144 22228
rect 40714 22188 41144 22216
rect 40714 22185 40726 22188
rect 40668 22179 40726 22185
rect 41138 22176 41144 22188
rect 41196 22176 41202 22228
rect 43530 22176 43536 22228
rect 43588 22216 43594 22228
rect 45554 22216 45560 22228
rect 43588 22188 45560 22216
rect 43588 22176 43594 22188
rect 45554 22176 45560 22188
rect 45612 22176 45618 22228
rect 47854 22176 47860 22228
rect 47912 22216 47918 22228
rect 48314 22216 48320 22228
rect 47912 22188 48320 22216
rect 47912 22176 47918 22188
rect 48314 22176 48320 22188
rect 48372 22176 48378 22228
rect 49694 22176 49700 22228
rect 49752 22176 49758 22228
rect 33134 22108 33140 22160
rect 33192 22108 33198 22160
rect 42242 22108 42248 22160
rect 42300 22148 42306 22160
rect 45278 22148 45284 22160
rect 42300 22120 45284 22148
rect 42300 22108 42306 22120
rect 45278 22108 45284 22120
rect 45336 22108 45342 22160
rect 47765 22151 47823 22157
rect 47765 22117 47777 22151
rect 47811 22148 47823 22151
rect 48038 22148 48044 22160
rect 47811 22120 48044 22148
rect 47811 22117 47823 22120
rect 47765 22111 47823 22117
rect 48038 22108 48044 22120
rect 48096 22108 48102 22160
rect 52914 22108 52920 22160
rect 52972 22148 52978 22160
rect 53650 22148 53656 22160
rect 52972 22120 53656 22148
rect 52972 22108 52978 22120
rect 53650 22108 53656 22120
rect 53708 22108 53714 22160
rect 33014 22052 33548 22080
rect 29549 22015 29607 22021
rect 29549 22012 29561 22015
rect 29380 21984 29561 22012
rect 29549 21981 29561 21984
rect 29595 21981 29607 22015
rect 29549 21975 29607 21981
rect 31202 21972 31208 22024
rect 31260 21972 31266 22024
rect 33520 22021 33548 22052
rect 34716 22052 35571 22080
rect 33321 22015 33379 22021
rect 33321 21981 33333 22015
rect 33367 21981 33379 22015
rect 33321 21975 33379 21981
rect 33505 22015 33563 22021
rect 33505 21981 33517 22015
rect 33551 21981 33563 22015
rect 33505 21975 33563 21981
rect 26634 21916 27384 21944
rect 27430 21904 27436 21956
rect 27488 21944 27494 21956
rect 27525 21947 27583 21953
rect 27525 21944 27537 21947
rect 27488 21916 27537 21944
rect 27488 21904 27494 21916
rect 27525 21913 27537 21916
rect 27571 21944 27583 21947
rect 27982 21944 27988 21956
rect 27571 21916 27988 21944
rect 27571 21913 27583 21916
rect 27525 21907 27583 21913
rect 27982 21904 27988 21916
rect 28040 21904 28046 21956
rect 31938 21944 31944 21956
rect 31864 21916 31944 21944
rect 19484 21848 20024 21876
rect 19484 21836 19490 21848
rect 20070 21836 20076 21888
rect 20128 21876 20134 21888
rect 20346 21876 20352 21888
rect 20128 21848 20352 21876
rect 20128 21836 20134 21848
rect 20346 21836 20352 21848
rect 20404 21836 20410 21888
rect 21542 21836 21548 21888
rect 21600 21876 21606 21888
rect 22278 21876 22284 21888
rect 21600 21848 22284 21876
rect 21600 21836 21606 21848
rect 22278 21836 22284 21848
rect 22336 21876 22342 21888
rect 23290 21876 23296 21888
rect 22336 21848 23296 21876
rect 22336 21836 22342 21848
rect 23290 21836 23296 21848
rect 23348 21876 23354 21888
rect 23753 21879 23811 21885
rect 23753 21876 23765 21879
rect 23348 21848 23765 21876
rect 23348 21836 23354 21848
rect 23753 21845 23765 21848
rect 23799 21876 23811 21879
rect 24026 21876 24032 21888
rect 23799 21848 24032 21876
rect 23799 21845 23811 21848
rect 23753 21839 23811 21845
rect 24026 21836 24032 21848
rect 24084 21836 24090 21888
rect 28718 21836 28724 21888
rect 28776 21876 28782 21888
rect 29733 21879 29791 21885
rect 29733 21876 29745 21879
rect 28776 21848 29745 21876
rect 28776 21836 28782 21848
rect 29733 21845 29745 21848
rect 29779 21845 29791 21879
rect 29733 21839 29791 21845
rect 31018 21836 31024 21888
rect 31076 21876 31082 21888
rect 31662 21876 31668 21888
rect 31076 21848 31668 21876
rect 31076 21836 31082 21848
rect 31662 21836 31668 21848
rect 31720 21876 31726 21888
rect 31864 21876 31892 21916
rect 31938 21904 31944 21916
rect 31996 21904 32002 21956
rect 33336 21944 33364 21975
rect 33594 21972 33600 22024
rect 33652 22012 33658 22024
rect 34606 22012 34612 22024
rect 33652 21984 34612 22012
rect 33652 21972 33658 21984
rect 34606 21972 34612 21984
rect 34664 21972 34670 22024
rect 34716 21956 34744 22052
rect 35342 21972 35348 22024
rect 35400 21972 35406 22024
rect 35437 22015 35495 22021
rect 35437 21981 35449 22015
rect 35483 21981 35495 22015
rect 35437 21975 35495 21981
rect 34698 21944 34704 21956
rect 33336 21916 34704 21944
rect 31720 21848 31892 21876
rect 31720 21836 31726 21848
rect 32214 21836 32220 21888
rect 32272 21876 32278 21888
rect 33336 21876 33364 21916
rect 34698 21904 34704 21916
rect 34756 21904 34762 21956
rect 32272 21848 33364 21876
rect 32272 21836 32278 21848
rect 35066 21836 35072 21888
rect 35124 21836 35130 21888
rect 35158 21836 35164 21888
rect 35216 21836 35222 21888
rect 35342 21836 35348 21888
rect 35400 21876 35406 21888
rect 35452 21876 35480 21975
rect 35400 21848 35480 21876
rect 35543 21876 35571 22052
rect 37458 22040 37464 22092
rect 37516 22080 37522 22092
rect 38013 22083 38071 22089
rect 38013 22080 38025 22083
rect 37516 22052 38025 22080
rect 37516 22040 37522 22052
rect 38013 22049 38025 22052
rect 38059 22049 38071 22083
rect 38013 22043 38071 22049
rect 44174 22040 44180 22092
rect 44232 22080 44238 22092
rect 46842 22080 46848 22092
rect 44232 22052 46848 22080
rect 44232 22040 44238 22052
rect 46842 22040 46848 22052
rect 46900 22040 46906 22092
rect 50246 22080 50252 22092
rect 48424 22052 50252 22080
rect 35710 21972 35716 22024
rect 35768 21972 35774 22024
rect 35802 21972 35808 22024
rect 35860 21972 35866 22024
rect 37642 21972 37648 22024
rect 37700 21972 37706 22024
rect 40402 21972 40408 22024
rect 40460 21972 40466 22024
rect 44450 21972 44456 22024
rect 44508 22012 44514 22024
rect 45005 22015 45063 22021
rect 45005 22012 45017 22015
rect 44508 21984 45017 22012
rect 44508 21972 44514 21984
rect 45005 21981 45017 21984
rect 45051 21981 45063 22015
rect 45186 22012 45192 22024
rect 45005 21975 45063 21981
rect 45112 21984 45192 22012
rect 37274 21904 37280 21956
rect 37332 21944 37338 21956
rect 42702 21944 42708 21956
rect 37332 21916 37412 21944
rect 41906 21916 42708 21944
rect 37332 21904 37338 21916
rect 35989 21879 36047 21885
rect 35989 21876 36001 21879
rect 35543 21848 36001 21876
rect 35400 21836 35406 21848
rect 35989 21845 36001 21848
rect 36035 21845 36047 21879
rect 37384 21876 37412 21916
rect 42702 21904 42708 21916
rect 42760 21904 42766 21956
rect 44818 21904 44824 21956
rect 44876 21944 44882 21956
rect 45112 21944 45140 21984
rect 45186 21972 45192 21984
rect 45244 21972 45250 22024
rect 47210 21972 47216 22024
rect 47268 22012 47274 22024
rect 47397 22015 47455 22021
rect 47397 22012 47409 22015
rect 47268 21984 47409 22012
rect 47268 21972 47274 21984
rect 47397 21981 47409 21984
rect 47443 22012 47455 22015
rect 47581 22015 47639 22021
rect 47581 22012 47593 22015
rect 47443 21984 47593 22012
rect 47443 21981 47455 21984
rect 47397 21975 47455 21981
rect 47581 21981 47593 21984
rect 47627 21981 47639 22015
rect 47581 21975 47639 21981
rect 47946 21972 47952 22024
rect 48004 22012 48010 22024
rect 48133 22015 48191 22021
rect 48133 22012 48145 22015
rect 48004 21984 48145 22012
rect 48004 21972 48010 21984
rect 48133 21981 48145 21984
rect 48179 21981 48191 22015
rect 48133 21975 48191 21981
rect 44876 21916 45140 21944
rect 45204 21916 45508 21944
rect 44876 21904 44882 21916
rect 38470 21876 38476 21888
rect 37384 21848 38476 21876
rect 35989 21839 36047 21845
rect 38470 21836 38476 21848
rect 38528 21836 38534 21888
rect 41598 21836 41604 21888
rect 41656 21876 41662 21888
rect 42153 21879 42211 21885
rect 42153 21876 42165 21879
rect 41656 21848 42165 21876
rect 41656 21836 41662 21848
rect 42153 21845 42165 21848
rect 42199 21876 42211 21879
rect 42337 21879 42395 21885
rect 42337 21876 42349 21879
rect 42199 21848 42349 21876
rect 42199 21845 42211 21848
rect 42153 21839 42211 21845
rect 42337 21845 42349 21848
rect 42383 21845 42395 21879
rect 42337 21839 42395 21845
rect 43898 21836 43904 21888
rect 43956 21876 43962 21888
rect 45204 21876 45232 21916
rect 43956 21848 45232 21876
rect 43956 21836 43962 21848
rect 45278 21836 45284 21888
rect 45336 21876 45342 21888
rect 45373 21879 45431 21885
rect 45373 21876 45385 21879
rect 45336 21848 45385 21876
rect 45336 21836 45342 21848
rect 45373 21845 45385 21848
rect 45419 21845 45431 21879
rect 45480 21876 45508 21916
rect 45554 21904 45560 21956
rect 45612 21944 45618 21956
rect 46474 21944 46480 21956
rect 45612 21916 46480 21944
rect 45612 21904 45618 21916
rect 46474 21904 46480 21916
rect 46532 21944 46538 21956
rect 47854 21944 47860 21956
rect 46532 21916 47860 21944
rect 46532 21904 46538 21916
rect 47854 21904 47860 21916
rect 47912 21904 47918 21956
rect 47302 21876 47308 21888
rect 45480 21848 47308 21876
rect 45373 21839 45431 21845
rect 47302 21836 47308 21848
rect 47360 21836 47366 21888
rect 47762 21836 47768 21888
rect 47820 21876 47826 21888
rect 47949 21879 48007 21885
rect 47949 21876 47961 21879
rect 47820 21848 47961 21876
rect 47820 21836 47826 21848
rect 47949 21845 47961 21848
rect 47995 21845 48007 21879
rect 48148 21876 48176 21975
rect 48314 21972 48320 22024
rect 48372 21972 48378 22024
rect 48225 21947 48283 21953
rect 48225 21913 48237 21947
rect 48271 21944 48283 21947
rect 48424 21944 48452 22052
rect 50246 22040 50252 22052
rect 50304 22040 50310 22092
rect 53101 22083 53159 22089
rect 53101 22080 53113 22083
rect 52380 22052 53113 22080
rect 48501 22015 48559 22021
rect 48501 21981 48513 22015
rect 48547 22012 48559 22015
rect 48682 22012 48688 22024
rect 48547 21984 48688 22012
rect 48547 21981 48559 21984
rect 48501 21975 48559 21981
rect 48682 21972 48688 21984
rect 48740 21972 48746 22024
rect 48961 22015 49019 22021
rect 48961 21981 48973 22015
rect 49007 22012 49019 22015
rect 49050 22012 49056 22024
rect 49007 21984 49056 22012
rect 49007 21981 49019 21984
rect 48961 21975 49019 21981
rect 49050 21972 49056 21984
rect 49108 21972 49114 22024
rect 49145 22015 49203 22021
rect 49145 21981 49157 22015
rect 49191 22012 49203 22015
rect 49326 22012 49332 22024
rect 49191 21984 49332 22012
rect 49191 21981 49203 21984
rect 49145 21975 49203 21981
rect 49326 21972 49332 21984
rect 49384 22012 49390 22024
rect 52380 22021 52408 22052
rect 53101 22049 53113 22052
rect 53147 22080 53159 22083
rect 55674 22080 55680 22092
rect 53147 22052 55680 22080
rect 53147 22049 53159 22052
rect 53101 22043 53159 22049
rect 55674 22040 55680 22052
rect 55732 22040 55738 22092
rect 49513 22015 49571 22021
rect 49513 22012 49525 22015
rect 49384 21984 49525 22012
rect 49384 21972 49390 21984
rect 49513 21981 49525 21984
rect 49559 21981 49571 22015
rect 49513 21975 49571 21981
rect 52365 22015 52423 22021
rect 52365 21981 52377 22015
rect 52411 21981 52423 22015
rect 52365 21975 52423 21981
rect 54021 22015 54079 22021
rect 54021 21981 54033 22015
rect 54067 22012 54079 22015
rect 54478 22012 54484 22024
rect 54067 21984 54484 22012
rect 54067 21981 54079 21984
rect 54021 21975 54079 21981
rect 48271 21916 48452 21944
rect 49528 21944 49556 21975
rect 54478 21972 54484 21984
rect 54536 21972 54542 22024
rect 56134 21972 56140 22024
rect 56192 22012 56198 22024
rect 56873 22015 56931 22021
rect 56873 22012 56885 22015
rect 56192 21984 56885 22012
rect 56192 21972 56198 21984
rect 56873 21981 56885 21984
rect 56919 21981 56931 22015
rect 56873 21975 56931 21981
rect 52549 21947 52607 21953
rect 52549 21944 52561 21947
rect 49528 21916 52561 21944
rect 48271 21913 48283 21916
rect 48225 21907 48283 21913
rect 52549 21913 52561 21916
rect 52595 21944 52607 21947
rect 52825 21947 52883 21953
rect 52825 21944 52837 21947
rect 52595 21916 52837 21944
rect 52595 21913 52607 21916
rect 52549 21907 52607 21913
rect 52825 21913 52837 21916
rect 52871 21913 52883 21947
rect 52825 21907 52883 21913
rect 55398 21904 55404 21956
rect 55456 21944 55462 21956
rect 55677 21947 55735 21953
rect 55677 21944 55689 21947
rect 55456 21916 55689 21944
rect 55456 21904 55462 21916
rect 55677 21913 55689 21916
rect 55723 21913 55735 21947
rect 55677 21907 55735 21913
rect 57140 21947 57198 21953
rect 57140 21913 57152 21947
rect 57186 21944 57198 21947
rect 57514 21944 57520 21956
rect 57186 21916 57520 21944
rect 57186 21913 57198 21916
rect 57140 21907 57198 21913
rect 57514 21904 57520 21916
rect 57572 21904 57578 21956
rect 48498 21876 48504 21888
rect 48148 21848 48504 21876
rect 47949 21839 48007 21845
rect 48498 21836 48504 21848
rect 48556 21836 48562 21888
rect 48866 21836 48872 21888
rect 48924 21836 48930 21888
rect 49050 21836 49056 21888
rect 49108 21876 49114 21888
rect 49329 21879 49387 21885
rect 49329 21876 49341 21879
rect 49108 21848 49341 21876
rect 49108 21836 49114 21848
rect 49329 21845 49341 21848
rect 49375 21876 49387 21879
rect 49786 21876 49792 21888
rect 49375 21848 49792 21876
rect 49375 21845 49387 21848
rect 49329 21839 49387 21845
rect 49786 21836 49792 21848
rect 49844 21836 49850 21888
rect 50893 21879 50951 21885
rect 50893 21845 50905 21879
rect 50939 21876 50951 21879
rect 51350 21876 51356 21888
rect 50939 21848 51356 21876
rect 50939 21845 50951 21848
rect 50893 21839 50951 21845
rect 51350 21836 51356 21848
rect 51408 21836 51414 21888
rect 52086 21836 52092 21888
rect 52144 21876 52150 21888
rect 52181 21879 52239 21885
rect 52181 21876 52193 21879
rect 52144 21848 52193 21876
rect 52144 21836 52150 21848
rect 52181 21845 52193 21848
rect 52227 21845 52239 21879
rect 52181 21839 52239 21845
rect 52638 21836 52644 21888
rect 52696 21836 52702 21888
rect 53374 21836 53380 21888
rect 53432 21836 53438 21888
rect 55306 21836 55312 21888
rect 55364 21876 55370 21888
rect 55493 21879 55551 21885
rect 55493 21876 55505 21879
rect 55364 21848 55505 21876
rect 55364 21836 55370 21848
rect 55493 21845 55505 21848
rect 55539 21845 55551 21879
rect 55493 21839 55551 21845
rect 58250 21836 58256 21888
rect 58308 21876 58314 21888
rect 58434 21876 58440 21888
rect 58308 21848 58440 21876
rect 58308 21836 58314 21848
rect 58434 21836 58440 21848
rect 58492 21836 58498 21888
rect 1104 21786 58880 21808
rect 1104 21734 4874 21786
rect 4926 21734 4938 21786
rect 4990 21734 5002 21786
rect 5054 21734 5066 21786
rect 5118 21734 5130 21786
rect 5182 21734 35594 21786
rect 35646 21734 35658 21786
rect 35710 21734 35722 21786
rect 35774 21734 35786 21786
rect 35838 21734 35850 21786
rect 35902 21734 58880 21786
rect 1104 21712 58880 21734
rect 19429 21675 19487 21681
rect 19429 21641 19441 21675
rect 19475 21641 19487 21675
rect 19429 21635 19487 21641
rect 19061 21539 19119 21545
rect 19061 21505 19073 21539
rect 19107 21536 19119 21539
rect 19444 21536 19472 21635
rect 19978 21632 19984 21684
rect 20036 21632 20042 21684
rect 20162 21632 20168 21684
rect 20220 21632 20226 21684
rect 20438 21632 20444 21684
rect 20496 21672 20502 21684
rect 20898 21672 20904 21684
rect 20496 21644 20576 21672
rect 20496 21632 20502 21644
rect 19797 21607 19855 21613
rect 19797 21573 19809 21607
rect 19843 21604 19855 21607
rect 19996 21604 20024 21632
rect 20548 21613 20576 21644
rect 20640 21644 20904 21672
rect 20533 21607 20591 21613
rect 20533 21604 20545 21607
rect 19843 21576 20545 21604
rect 19843 21573 19855 21576
rect 19797 21567 19855 21573
rect 20533 21573 20545 21576
rect 20579 21573 20591 21607
rect 20533 21567 20591 21573
rect 19107 21508 19472 21536
rect 19608 21539 19666 21545
rect 19107 21505 19119 21508
rect 19061 21499 19119 21505
rect 19608 21505 19620 21539
rect 19654 21505 19666 21539
rect 19608 21499 19666 21505
rect 19337 21471 19395 21477
rect 19337 21437 19349 21471
rect 19383 21468 19395 21471
rect 19426 21468 19432 21480
rect 19383 21440 19432 21468
rect 19383 21437 19395 21440
rect 19337 21431 19395 21437
rect 19426 21428 19432 21440
rect 19484 21428 19490 21480
rect 19628 21400 19656 21499
rect 19702 21496 19708 21548
rect 19760 21496 19766 21548
rect 19978 21536 19984 21548
rect 19939 21508 19984 21536
rect 19978 21496 19984 21508
rect 20036 21496 20042 21548
rect 20073 21539 20131 21545
rect 20073 21505 20085 21539
rect 20119 21505 20131 21539
rect 20073 21499 20131 21505
rect 20088 21468 20116 21499
rect 20254 21496 20260 21548
rect 20312 21536 20318 21548
rect 20349 21539 20407 21545
rect 20349 21536 20361 21539
rect 20312 21508 20361 21536
rect 20312 21496 20318 21508
rect 20349 21505 20361 21508
rect 20395 21505 20407 21539
rect 20349 21499 20407 21505
rect 20438 21496 20444 21548
rect 20496 21496 20502 21548
rect 20640 21468 20668 21644
rect 20898 21632 20904 21644
rect 20956 21632 20962 21684
rect 23566 21632 23572 21684
rect 23624 21632 23630 21684
rect 26050 21672 26056 21684
rect 24504 21644 26056 21672
rect 23584 21604 23612 21632
rect 23661 21607 23719 21613
rect 23661 21604 23673 21607
rect 22388 21576 23673 21604
rect 22388 21548 22416 21576
rect 23661 21573 23673 21576
rect 23707 21573 23719 21607
rect 24394 21604 24400 21616
rect 23661 21567 23719 21573
rect 23952 21576 24400 21604
rect 20717 21539 20775 21545
rect 20717 21505 20729 21539
rect 20763 21536 20775 21539
rect 22370 21536 22376 21548
rect 20763 21508 22376 21536
rect 20763 21505 20775 21508
rect 20717 21499 20775 21505
rect 22370 21496 22376 21508
rect 22428 21496 22434 21548
rect 23564 21539 23622 21545
rect 23564 21505 23576 21539
rect 23610 21536 23622 21539
rect 23753 21539 23811 21545
rect 23610 21508 23704 21536
rect 23610 21505 23622 21508
rect 23564 21499 23622 21505
rect 23676 21480 23704 21508
rect 23753 21505 23765 21539
rect 23799 21536 23811 21539
rect 23842 21536 23848 21548
rect 23799 21508 23848 21536
rect 23799 21505 23811 21508
rect 23753 21499 23811 21505
rect 23658 21468 23664 21480
rect 20088 21440 20668 21468
rect 20824 21440 23664 21468
rect 20254 21400 20260 21412
rect 19628 21372 20260 21400
rect 20254 21360 20260 21372
rect 20312 21400 20318 21412
rect 20824 21400 20852 21440
rect 23658 21428 23664 21440
rect 23716 21428 23722 21480
rect 20312 21372 20852 21400
rect 23768 21400 23796 21499
rect 23842 21496 23848 21508
rect 23900 21496 23906 21548
rect 23952 21545 23980 21576
rect 24394 21564 24400 21576
rect 24452 21564 24458 21616
rect 23936 21539 23994 21545
rect 23936 21505 23948 21539
rect 23982 21505 23994 21539
rect 23936 21499 23994 21505
rect 24029 21539 24087 21545
rect 24029 21505 24041 21539
rect 24075 21505 24087 21539
rect 24029 21499 24087 21505
rect 24044 21468 24072 21499
rect 24118 21496 24124 21548
rect 24176 21496 24182 21548
rect 24504 21545 24532 21644
rect 26050 21632 26056 21644
rect 26108 21632 26114 21684
rect 27982 21632 27988 21684
rect 28040 21672 28046 21684
rect 30653 21675 30711 21681
rect 30653 21672 30665 21675
rect 28040 21644 30665 21672
rect 28040 21632 28046 21644
rect 30653 21641 30665 21644
rect 30699 21641 30711 21675
rect 30653 21635 30711 21641
rect 24578 21564 24584 21616
rect 24636 21604 24642 21616
rect 27522 21604 27528 21616
rect 24636 21576 26372 21604
rect 24636 21564 24642 21576
rect 24489 21539 24547 21545
rect 24489 21505 24501 21539
rect 24535 21505 24547 21539
rect 24489 21499 24547 21505
rect 24854 21496 24860 21548
rect 24912 21496 24918 21548
rect 26344 21545 26372 21576
rect 26988 21576 27528 21604
rect 26237 21539 26295 21545
rect 26237 21536 26249 21539
rect 26160 21508 26249 21536
rect 24872 21468 24900 21496
rect 25866 21468 25872 21480
rect 24044 21440 25872 21468
rect 25866 21428 25872 21440
rect 25924 21428 25930 21480
rect 23768 21372 24716 21400
rect 20312 21360 20318 21372
rect 18782 21292 18788 21344
rect 18840 21332 18846 21344
rect 18877 21335 18935 21341
rect 18877 21332 18889 21335
rect 18840 21304 18889 21332
rect 18840 21292 18846 21304
rect 18877 21301 18889 21304
rect 18923 21301 18935 21335
rect 18877 21295 18935 21301
rect 18966 21292 18972 21344
rect 19024 21332 19030 21344
rect 19245 21335 19303 21341
rect 19245 21332 19257 21335
rect 19024 21304 19257 21332
rect 19024 21292 19030 21304
rect 19245 21301 19257 21304
rect 19291 21332 19303 21335
rect 19334 21332 19340 21344
rect 19291 21304 19340 21332
rect 19291 21301 19303 21304
rect 19245 21295 19303 21301
rect 19334 21292 19340 21304
rect 19392 21332 19398 21344
rect 21542 21332 21548 21344
rect 19392 21304 21548 21332
rect 19392 21292 19398 21304
rect 21542 21292 21548 21304
rect 21600 21292 21606 21344
rect 23385 21335 23443 21341
rect 23385 21301 23397 21335
rect 23431 21332 23443 21335
rect 23842 21332 23848 21344
rect 23431 21304 23848 21332
rect 23431 21301 23443 21304
rect 23385 21295 23443 21301
rect 23842 21292 23848 21304
rect 23900 21292 23906 21344
rect 23934 21292 23940 21344
rect 23992 21332 23998 21344
rect 24305 21335 24363 21341
rect 24305 21332 24317 21335
rect 23992 21304 24317 21332
rect 23992 21292 23998 21304
rect 24305 21301 24317 21304
rect 24351 21332 24363 21335
rect 24578 21332 24584 21344
rect 24351 21304 24584 21332
rect 24351 21301 24363 21304
rect 24305 21295 24363 21301
rect 24578 21292 24584 21304
rect 24636 21292 24642 21344
rect 24688 21341 24716 21372
rect 24673 21335 24731 21341
rect 24673 21301 24685 21335
rect 24719 21332 24731 21335
rect 25590 21332 25596 21344
rect 24719 21304 25596 21332
rect 24719 21301 24731 21304
rect 24673 21295 24731 21301
rect 25590 21292 25596 21304
rect 25648 21292 25654 21344
rect 25869 21335 25927 21341
rect 25869 21301 25881 21335
rect 25915 21332 25927 21335
rect 26160 21332 26188 21508
rect 26237 21505 26249 21508
rect 26283 21505 26295 21539
rect 26237 21499 26295 21505
rect 26329 21539 26387 21545
rect 26329 21505 26341 21539
rect 26375 21505 26387 21539
rect 26329 21499 26387 21505
rect 26344 21468 26372 21499
rect 26602 21496 26608 21548
rect 26660 21496 26666 21548
rect 26988 21545 27016 21576
rect 27522 21564 27528 21576
rect 27580 21564 27586 21616
rect 28626 21604 28632 21616
rect 28474 21576 28632 21604
rect 28626 21564 28632 21576
rect 28684 21564 28690 21616
rect 29270 21564 29276 21616
rect 29328 21604 29334 21616
rect 29328 21576 29868 21604
rect 29328 21564 29334 21576
rect 29840 21545 29868 21576
rect 26973 21539 27031 21545
rect 26973 21505 26985 21539
rect 27019 21505 27031 21539
rect 26973 21499 27031 21505
rect 29457 21539 29515 21545
rect 29457 21505 29469 21539
rect 29503 21536 29515 21539
rect 29549 21539 29607 21545
rect 29549 21536 29561 21539
rect 29503 21508 29561 21536
rect 29503 21505 29515 21508
rect 29457 21499 29515 21505
rect 29549 21505 29561 21508
rect 29595 21505 29607 21539
rect 29549 21499 29607 21505
rect 29825 21539 29883 21545
rect 29825 21505 29837 21539
rect 29871 21505 29883 21539
rect 29825 21499 29883 21505
rect 29914 21496 29920 21548
rect 29972 21496 29978 21548
rect 30469 21539 30527 21545
rect 30469 21505 30481 21539
rect 30515 21505 30527 21539
rect 30668 21536 30696 21635
rect 31018 21632 31024 21684
rect 31076 21632 31082 21684
rect 32306 21632 32312 21684
rect 32364 21632 32370 21684
rect 32490 21632 32496 21684
rect 32548 21672 32554 21684
rect 32677 21675 32735 21681
rect 32677 21672 32689 21675
rect 32548 21644 32689 21672
rect 32548 21632 32554 21644
rect 32677 21641 32689 21644
rect 32723 21641 32735 21675
rect 32677 21635 32735 21641
rect 32858 21632 32864 21684
rect 32916 21672 32922 21684
rect 32953 21675 33011 21681
rect 32953 21672 32965 21675
rect 32916 21644 32965 21672
rect 32916 21632 32922 21644
rect 32953 21641 32965 21644
rect 32999 21641 33011 21675
rect 32953 21635 33011 21641
rect 34514 21632 34520 21684
rect 34572 21672 34578 21684
rect 34701 21675 34759 21681
rect 34701 21672 34713 21675
rect 34572 21644 34713 21672
rect 34572 21632 34578 21644
rect 34701 21641 34713 21644
rect 34747 21641 34759 21675
rect 34701 21635 34759 21641
rect 36722 21632 36728 21684
rect 36780 21672 36786 21684
rect 42886 21672 42892 21684
rect 36780 21644 42892 21672
rect 36780 21632 36786 21644
rect 42886 21632 42892 21644
rect 42944 21632 42950 21684
rect 43990 21632 43996 21684
rect 44048 21672 44054 21684
rect 44634 21672 44640 21684
rect 44048 21644 44640 21672
rect 44048 21632 44054 21644
rect 44634 21632 44640 21644
rect 44692 21672 44698 21684
rect 45554 21672 45560 21684
rect 44692 21644 45560 21672
rect 44692 21632 44698 21644
rect 45554 21632 45560 21644
rect 45612 21632 45618 21684
rect 46017 21675 46075 21681
rect 46017 21641 46029 21675
rect 46063 21672 46075 21675
rect 48682 21672 48688 21684
rect 46063 21644 48688 21672
rect 46063 21641 46075 21644
rect 46017 21635 46075 21641
rect 32324 21604 32352 21632
rect 32401 21607 32459 21613
rect 32401 21604 32413 21607
rect 31680 21576 31892 21604
rect 32324 21576 32413 21604
rect 30837 21539 30895 21545
rect 30837 21536 30849 21539
rect 30668 21508 30849 21536
rect 30469 21499 30527 21505
rect 30837 21505 30849 21508
rect 30883 21505 30895 21539
rect 30837 21499 30895 21505
rect 26789 21471 26847 21477
rect 26344 21440 26740 21468
rect 26234 21360 26240 21412
rect 26292 21400 26298 21412
rect 26421 21403 26479 21409
rect 26421 21400 26433 21403
rect 26292 21372 26433 21400
rect 26292 21360 26298 21372
rect 26421 21369 26433 21372
rect 26467 21369 26479 21403
rect 26421 21363 26479 21369
rect 26326 21332 26332 21344
rect 25915 21304 26332 21332
rect 25915 21301 25927 21304
rect 25869 21295 25927 21301
rect 26326 21292 26332 21304
rect 26384 21292 26390 21344
rect 26712 21332 26740 21440
rect 26789 21437 26801 21471
rect 26835 21468 26847 21471
rect 27249 21471 27307 21477
rect 27249 21468 27261 21471
rect 26835 21440 27261 21468
rect 26835 21437 26847 21440
rect 26789 21431 26847 21437
rect 27249 21437 27261 21440
rect 27295 21437 27307 21471
rect 27249 21431 27307 21437
rect 27706 21428 27712 21480
rect 27764 21468 27770 21480
rect 28813 21471 28871 21477
rect 28813 21468 28825 21471
rect 27764 21440 28825 21468
rect 27764 21428 27770 21440
rect 28813 21437 28825 21440
rect 28859 21437 28871 21471
rect 30484 21468 30512 21499
rect 31570 21496 31576 21548
rect 31628 21496 31634 21548
rect 31680 21545 31708 21576
rect 31665 21539 31723 21545
rect 31665 21505 31677 21539
rect 31711 21505 31723 21539
rect 31665 21499 31723 21505
rect 31202 21468 31208 21480
rect 30484 21440 31208 21468
rect 28813 21431 28871 21437
rect 31202 21428 31208 21440
rect 31260 21428 31266 21480
rect 30006 21400 30012 21412
rect 29656 21372 30012 21400
rect 28534 21332 28540 21344
rect 26712 21304 28540 21332
rect 28534 21292 28540 21304
rect 28592 21332 28598 21344
rect 29656 21341 29684 21372
rect 30006 21360 30012 21372
rect 30064 21400 30070 21412
rect 31864 21400 31892 21576
rect 32401 21573 32413 21576
rect 32447 21573 32459 21607
rect 33594 21604 33600 21616
rect 32401 21567 32459 21573
rect 32508 21576 33600 21604
rect 31941 21539 31999 21545
rect 31941 21505 31953 21539
rect 31987 21536 31999 21539
rect 32125 21539 32183 21545
rect 32125 21536 32137 21539
rect 31987 21508 32137 21536
rect 31987 21505 31999 21508
rect 31941 21499 31999 21505
rect 32125 21505 32137 21508
rect 32171 21505 32183 21539
rect 32125 21499 32183 21505
rect 32140 21468 32168 21499
rect 32214 21496 32220 21548
rect 32272 21536 32278 21548
rect 32508 21545 32536 21576
rect 33594 21564 33600 21576
rect 33652 21564 33658 21616
rect 36170 21564 36176 21616
rect 36228 21604 36234 21616
rect 37274 21604 37280 21616
rect 36228 21576 37280 21604
rect 36228 21564 36234 21576
rect 37274 21564 37280 21576
rect 37332 21564 37338 21616
rect 39298 21564 39304 21616
rect 39356 21604 39362 21616
rect 46860 21604 46888 21644
rect 48682 21632 48688 21644
rect 48740 21632 48746 21684
rect 48866 21632 48872 21684
rect 48924 21672 48930 21684
rect 50798 21672 50804 21684
rect 48924 21644 49188 21672
rect 48924 21632 48930 21644
rect 39356 21576 45034 21604
rect 46768 21576 46888 21604
rect 47397 21607 47455 21613
rect 39356 21564 39362 21576
rect 32309 21539 32367 21545
rect 32309 21536 32321 21539
rect 32272 21508 32321 21536
rect 32272 21496 32278 21508
rect 32309 21505 32321 21508
rect 32355 21505 32367 21539
rect 32309 21499 32367 21505
rect 32493 21539 32551 21545
rect 32493 21505 32505 21539
rect 32539 21505 32551 21539
rect 32493 21499 32551 21505
rect 32766 21496 32772 21548
rect 32824 21496 32830 21548
rect 34054 21496 34060 21548
rect 34112 21496 34118 21548
rect 34146 21496 34152 21548
rect 34204 21496 34210 21548
rect 34333 21539 34391 21545
rect 34333 21505 34345 21539
rect 34379 21505 34391 21539
rect 34333 21499 34391 21505
rect 34164 21468 34192 21496
rect 32140 21440 34192 21468
rect 34348 21412 34376 21499
rect 34422 21496 34428 21548
rect 34480 21496 34486 21548
rect 34514 21496 34520 21548
rect 34572 21545 34578 21548
rect 34572 21536 34580 21545
rect 34572 21508 34617 21536
rect 34572 21499 34580 21508
rect 34572 21496 34578 21499
rect 35158 21496 35164 21548
rect 35216 21496 35222 21548
rect 41506 21496 41512 21548
rect 41564 21536 41570 21548
rect 41874 21536 41880 21548
rect 41564 21508 41880 21536
rect 41564 21496 41570 21508
rect 41874 21496 41880 21508
rect 41932 21496 41938 21548
rect 41969 21539 42027 21545
rect 41969 21505 41981 21539
rect 42015 21505 42027 21539
rect 41969 21499 42027 21505
rect 42245 21539 42303 21545
rect 42245 21505 42257 21539
rect 42291 21536 42303 21539
rect 42978 21536 42984 21548
rect 42291 21508 42984 21536
rect 42291 21505 42303 21508
rect 42245 21499 42303 21505
rect 34793 21471 34851 21477
rect 34793 21437 34805 21471
rect 34839 21468 34851 21471
rect 35434 21468 35440 21480
rect 34839 21440 35440 21468
rect 34839 21437 34851 21440
rect 34793 21431 34851 21437
rect 35434 21428 35440 21440
rect 35492 21428 35498 21480
rect 35894 21428 35900 21480
rect 35952 21468 35958 21480
rect 36078 21468 36084 21480
rect 35952 21440 36084 21468
rect 35952 21428 35958 21440
rect 36078 21428 36084 21440
rect 36136 21428 36142 21480
rect 41984 21468 42012 21499
rect 42978 21496 42984 21508
rect 43036 21496 43042 21548
rect 46768 21545 46796 21576
rect 47397 21573 47409 21607
rect 47443 21604 47455 21607
rect 47946 21604 47952 21616
rect 47443 21576 47952 21604
rect 47443 21573 47455 21576
rect 47397 21567 47455 21573
rect 47946 21564 47952 21576
rect 48004 21564 48010 21616
rect 49160 21604 49188 21644
rect 49344 21644 50804 21672
rect 49344 21616 49372 21644
rect 50798 21632 50804 21644
rect 50856 21672 50862 21684
rect 51994 21672 52000 21684
rect 50856 21644 52000 21672
rect 50856 21632 50862 21644
rect 51994 21632 52000 21644
rect 52052 21632 52058 21684
rect 53374 21672 53380 21684
rect 52104 21644 53380 21672
rect 49082 21590 49188 21604
rect 49068 21576 49188 21590
rect 46753 21539 46811 21545
rect 46753 21505 46765 21539
rect 46799 21505 46811 21539
rect 46753 21499 46811 21505
rect 46842 21496 46848 21548
rect 46900 21536 46906 21548
rect 47581 21539 47639 21545
rect 47581 21536 47593 21539
rect 46900 21508 47593 21536
rect 46900 21496 46906 21508
rect 47581 21505 47593 21508
rect 47627 21505 47639 21539
rect 49068 21536 49096 21576
rect 49326 21564 49332 21616
rect 49384 21564 49390 21616
rect 51442 21604 51448 21616
rect 51290 21576 51448 21604
rect 51442 21564 51448 21576
rect 51500 21564 51506 21616
rect 52104 21545 52132 21644
rect 53374 21632 53380 21644
rect 53432 21632 53438 21684
rect 54386 21632 54392 21684
rect 54444 21672 54450 21684
rect 55030 21672 55036 21684
rect 54444 21644 55036 21672
rect 54444 21632 54450 21644
rect 55030 21632 55036 21644
rect 55088 21632 55094 21684
rect 55769 21675 55827 21681
rect 55769 21641 55781 21675
rect 55815 21672 55827 21675
rect 55858 21672 55864 21684
rect 55815 21644 55864 21672
rect 55815 21641 55827 21644
rect 55769 21635 55827 21641
rect 55858 21632 55864 21644
rect 55916 21632 55922 21684
rect 57514 21632 57520 21684
rect 57572 21632 57578 21684
rect 52549 21607 52607 21613
rect 52549 21573 52561 21607
rect 52595 21604 52607 21607
rect 53009 21607 53067 21613
rect 53009 21604 53021 21607
rect 52595 21576 53021 21604
rect 52595 21573 52607 21576
rect 52549 21567 52607 21573
rect 53009 21573 53021 21576
rect 53055 21573 53067 21607
rect 53009 21567 53067 21573
rect 53650 21564 53656 21616
rect 53708 21564 53714 21616
rect 54662 21564 54668 21616
rect 54720 21604 54726 21616
rect 54757 21607 54815 21613
rect 54757 21604 54769 21607
rect 54720 21576 54769 21604
rect 54720 21564 54726 21576
rect 54757 21573 54769 21576
rect 54803 21604 54815 21607
rect 55122 21604 55128 21616
rect 54803 21576 55128 21604
rect 54803 21573 54815 21576
rect 54757 21567 54815 21573
rect 55122 21564 55128 21576
rect 55180 21604 55186 21616
rect 55953 21607 56011 21613
rect 55953 21604 55965 21607
rect 55180 21576 55965 21604
rect 55180 21564 55186 21576
rect 55953 21573 55965 21576
rect 55999 21573 56011 21607
rect 55953 21567 56011 21573
rect 56686 21564 56692 21616
rect 56744 21604 56750 21616
rect 56962 21604 56968 21616
rect 56744 21576 56968 21604
rect 56744 21564 56750 21576
rect 56962 21564 56968 21576
rect 57020 21604 57026 21616
rect 57020 21576 57192 21604
rect 57020 21564 57026 21576
rect 52089 21539 52147 21545
rect 49068 21508 50379 21536
rect 47581 21499 47639 21505
rect 43070 21468 43076 21480
rect 41984 21440 43076 21468
rect 43070 21428 43076 21440
rect 43128 21428 43134 21480
rect 44174 21428 44180 21480
rect 44232 21468 44238 21480
rect 44269 21471 44327 21477
rect 44269 21468 44281 21471
rect 44232 21440 44281 21468
rect 44232 21428 44238 21440
rect 44269 21437 44281 21440
rect 44315 21437 44327 21471
rect 44269 21431 44327 21437
rect 44545 21471 44603 21477
rect 44545 21437 44557 21471
rect 44591 21468 44603 21471
rect 45002 21468 45008 21480
rect 44591 21440 45008 21468
rect 44591 21437 44603 21440
rect 44545 21431 44603 21437
rect 45002 21428 45008 21440
rect 45060 21428 45066 21480
rect 47486 21428 47492 21480
rect 47544 21468 47550 21480
rect 47857 21471 47915 21477
rect 47857 21468 47869 21471
rect 47544 21440 47869 21468
rect 47544 21428 47550 21440
rect 47857 21437 47869 21440
rect 47903 21437 47915 21471
rect 47857 21431 47915 21437
rect 47946 21428 47952 21480
rect 48004 21468 48010 21480
rect 48866 21468 48872 21480
rect 48004 21440 48872 21468
rect 48004 21428 48010 21440
rect 48866 21428 48872 21440
rect 48924 21428 48930 21480
rect 49418 21468 49424 21480
rect 48976 21440 49424 21468
rect 33134 21400 33140 21412
rect 30064 21372 31754 21400
rect 31864 21372 33140 21400
rect 30064 21360 30070 21372
rect 28721 21335 28779 21341
rect 28721 21332 28733 21335
rect 28592 21304 28733 21332
rect 28592 21292 28598 21304
rect 28721 21301 28733 21304
rect 28767 21301 28779 21335
rect 28721 21295 28779 21301
rect 29641 21335 29699 21341
rect 29641 21301 29653 21335
rect 29687 21301 29699 21335
rect 29641 21295 29699 21301
rect 30098 21292 30104 21344
rect 30156 21292 30162 21344
rect 31389 21335 31447 21341
rect 31389 21301 31401 21335
rect 31435 21332 31447 21335
rect 31570 21332 31576 21344
rect 31435 21304 31576 21332
rect 31435 21301 31447 21304
rect 31389 21295 31447 21301
rect 31570 21292 31576 21304
rect 31628 21292 31634 21344
rect 31726 21332 31754 21372
rect 33134 21360 33140 21372
rect 33192 21360 33198 21412
rect 34330 21360 34336 21412
rect 34388 21400 34394 21412
rect 39666 21400 39672 21412
rect 34388 21372 34744 21400
rect 34388 21360 34394 21372
rect 31849 21335 31907 21341
rect 31849 21332 31861 21335
rect 31726 21304 31861 21332
rect 31849 21301 31861 21304
rect 31895 21332 31907 21335
rect 32858 21332 32864 21344
rect 31895 21304 32864 21332
rect 31895 21301 31907 21304
rect 31849 21295 31907 21301
rect 32858 21292 32864 21304
rect 32916 21292 32922 21344
rect 34716 21332 34744 21372
rect 35912 21372 39672 21400
rect 35066 21332 35072 21344
rect 34716 21304 35072 21332
rect 35066 21292 35072 21304
rect 35124 21332 35130 21344
rect 35912 21332 35940 21372
rect 39666 21360 39672 21372
rect 39724 21400 39730 21412
rect 40310 21400 40316 21412
rect 39724 21372 40316 21400
rect 39724 21360 39730 21372
rect 40310 21360 40316 21372
rect 40368 21360 40374 21412
rect 41230 21360 41236 21412
rect 41288 21400 41294 21412
rect 41601 21403 41659 21409
rect 41601 21400 41613 21403
rect 41288 21372 41613 21400
rect 41288 21360 41294 21372
rect 41601 21369 41613 21372
rect 41647 21400 41659 21403
rect 42150 21400 42156 21412
rect 41647 21372 42156 21400
rect 41647 21369 41659 21372
rect 41601 21363 41659 21369
rect 42150 21360 42156 21372
rect 42208 21360 42214 21412
rect 46032 21372 47716 21400
rect 35124 21304 35940 21332
rect 35124 21292 35130 21304
rect 36078 21292 36084 21344
rect 36136 21332 36142 21344
rect 36587 21335 36645 21341
rect 36587 21332 36599 21335
rect 36136 21304 36599 21332
rect 36136 21292 36142 21304
rect 36587 21301 36599 21304
rect 36633 21301 36645 21335
rect 36587 21295 36645 21301
rect 41690 21292 41696 21344
rect 41748 21292 41754 21344
rect 44542 21292 44548 21344
rect 44600 21332 44606 21344
rect 46032 21332 46060 21372
rect 44600 21304 46060 21332
rect 44600 21292 44606 21304
rect 46106 21292 46112 21344
rect 46164 21292 46170 21344
rect 47688 21332 47716 21372
rect 48976 21332 49004 21440
rect 49418 21428 49424 21440
rect 49476 21468 49482 21480
rect 49973 21471 50031 21477
rect 49973 21468 49985 21471
rect 49476 21440 49985 21468
rect 49476 21428 49482 21440
rect 49973 21437 49985 21440
rect 50019 21437 50031 21471
rect 49973 21431 50031 21437
rect 50246 21428 50252 21480
rect 50304 21428 50310 21480
rect 49050 21360 49056 21412
rect 49108 21400 49114 21412
rect 49108 21372 49464 21400
rect 49108 21360 49114 21372
rect 49436 21341 49464 21372
rect 49329 21335 49387 21341
rect 49329 21332 49341 21335
rect 47688 21304 49341 21332
rect 49329 21301 49341 21304
rect 49375 21301 49387 21335
rect 49329 21295 49387 21301
rect 49421 21335 49479 21341
rect 49421 21301 49433 21335
rect 49467 21301 49479 21335
rect 50351 21332 50379 21508
rect 52089 21505 52101 21539
rect 52135 21505 52147 21539
rect 52089 21499 52147 21505
rect 52365 21539 52423 21545
rect 52365 21505 52377 21539
rect 52411 21536 52423 21539
rect 52454 21536 52460 21548
rect 52411 21508 52460 21536
rect 52411 21505 52423 21508
rect 52365 21499 52423 21505
rect 52454 21496 52460 21508
rect 52512 21496 52518 21548
rect 54478 21496 54484 21548
rect 54536 21536 54542 21548
rect 54573 21539 54631 21545
rect 54573 21536 54585 21539
rect 54536 21508 54585 21536
rect 54536 21496 54542 21508
rect 54573 21505 54585 21508
rect 54619 21505 54631 21539
rect 54573 21499 54631 21505
rect 54849 21539 54907 21545
rect 54849 21505 54861 21539
rect 54895 21505 54907 21539
rect 54849 21499 54907 21505
rect 50982 21428 50988 21480
rect 51040 21468 51046 21480
rect 51721 21471 51779 21477
rect 51721 21468 51733 21471
rect 51040 21440 51733 21468
rect 51040 21428 51046 21440
rect 51721 21437 51733 21440
rect 51767 21437 51779 21471
rect 51997 21471 52055 21477
rect 51997 21468 52009 21471
rect 51721 21431 51779 21437
rect 51920 21440 52009 21468
rect 51920 21400 51948 21440
rect 51997 21437 52009 21440
rect 52043 21437 52055 21471
rect 51997 21431 52055 21437
rect 52733 21471 52791 21477
rect 52733 21437 52745 21471
rect 52779 21437 52791 21471
rect 54864 21468 54892 21499
rect 54938 21496 54944 21548
rect 54996 21496 55002 21548
rect 55030 21496 55036 21548
rect 55088 21536 55094 21548
rect 55217 21539 55275 21545
rect 55217 21536 55229 21539
rect 55088 21508 55229 21536
rect 55088 21496 55094 21508
rect 55217 21505 55229 21508
rect 55263 21505 55275 21539
rect 55217 21499 55275 21505
rect 55493 21539 55551 21545
rect 55493 21505 55505 21539
rect 55539 21505 55551 21539
rect 55493 21499 55551 21505
rect 55508 21468 55536 21499
rect 55582 21496 55588 21548
rect 55640 21496 55646 21548
rect 56137 21539 56195 21545
rect 56137 21505 56149 21539
rect 56183 21505 56195 21539
rect 56137 21499 56195 21505
rect 52733 21431 52791 21437
rect 54588 21440 54892 21468
rect 55140 21440 55536 21468
rect 52362 21400 52368 21412
rect 51920 21372 52368 21400
rect 51534 21332 51540 21344
rect 50351 21304 51540 21332
rect 49421 21295 49479 21301
rect 51534 21292 51540 21304
rect 51592 21292 51598 21344
rect 51718 21292 51724 21344
rect 51776 21332 51782 21344
rect 51920 21332 51948 21372
rect 52362 21360 52368 21372
rect 52420 21400 52426 21412
rect 52748 21400 52776 21431
rect 54588 21412 54616 21440
rect 52420 21372 52776 21400
rect 52420 21360 52426 21372
rect 54570 21360 54576 21412
rect 54628 21360 54634 21412
rect 55140 21409 55168 21440
rect 55125 21403 55183 21409
rect 55125 21369 55137 21403
rect 55171 21369 55183 21403
rect 55125 21363 55183 21369
rect 51776 21304 51948 21332
rect 51776 21292 51782 21304
rect 52178 21292 52184 21344
rect 52236 21332 52242 21344
rect 53558 21332 53564 21344
rect 52236 21304 53564 21332
rect 52236 21292 52242 21304
rect 53558 21292 53564 21304
rect 53616 21292 53622 21344
rect 54478 21292 54484 21344
rect 54536 21292 54542 21344
rect 55306 21292 55312 21344
rect 55364 21292 55370 21344
rect 55674 21292 55680 21344
rect 55732 21332 55738 21344
rect 56152 21332 56180 21499
rect 56870 21496 56876 21548
rect 56928 21496 56934 21548
rect 57164 21545 57192 21576
rect 57057 21539 57115 21545
rect 57057 21505 57069 21539
rect 57103 21505 57115 21539
rect 57057 21499 57115 21505
rect 57149 21539 57207 21545
rect 57149 21505 57161 21539
rect 57195 21505 57207 21539
rect 57149 21499 57207 21505
rect 57241 21539 57299 21545
rect 57241 21505 57253 21539
rect 57287 21536 57299 21539
rect 57885 21539 57943 21545
rect 57885 21536 57897 21539
rect 57287 21508 57897 21536
rect 57287 21505 57299 21508
rect 57241 21499 57299 21505
rect 57885 21505 57897 21508
rect 57931 21505 57943 21539
rect 57885 21499 57943 21505
rect 56686 21428 56692 21480
rect 56744 21468 56750 21480
rect 57072 21468 57100 21499
rect 58434 21496 58440 21548
rect 58492 21496 58498 21548
rect 56744 21440 57100 21468
rect 56744 21428 56750 21440
rect 56321 21335 56379 21341
rect 56321 21332 56333 21335
rect 55732 21304 56333 21332
rect 55732 21292 55738 21304
rect 56321 21301 56333 21304
rect 56367 21301 56379 21335
rect 56321 21295 56379 21301
rect 1104 21242 58880 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 58880 21242
rect 1104 21168 58880 21190
rect 20162 21128 20168 21140
rect 18800 21100 20168 21128
rect 18800 20933 18828 21100
rect 20162 21088 20168 21100
rect 20220 21088 20226 21140
rect 25133 21131 25191 21137
rect 25133 21128 25145 21131
rect 22020 21100 25145 21128
rect 18966 21020 18972 21072
rect 19024 21020 19030 21072
rect 19076 21032 19380 21060
rect 19076 20933 19104 21032
rect 19242 20952 19248 21004
rect 19300 20952 19306 21004
rect 19352 20992 19380 21032
rect 19978 20992 19984 21004
rect 19352 20964 19984 20992
rect 19978 20952 19984 20964
rect 20036 20952 20042 21004
rect 22020 20992 22048 21100
rect 25133 21097 25145 21100
rect 25179 21097 25191 21131
rect 25133 21091 25191 21097
rect 25866 21088 25872 21140
rect 25924 21088 25930 21140
rect 26053 21131 26111 21137
rect 26053 21097 26065 21131
rect 26099 21128 26111 21131
rect 26602 21128 26608 21140
rect 26099 21100 26608 21128
rect 26099 21097 26111 21100
rect 26053 21091 26111 21097
rect 26602 21088 26608 21100
rect 26660 21088 26666 21140
rect 29107 21131 29165 21137
rect 29107 21097 29119 21131
rect 29153 21128 29165 21131
rect 30098 21128 30104 21140
rect 29153 21100 30104 21128
rect 29153 21097 29165 21100
rect 29107 21091 29165 21097
rect 30098 21088 30104 21100
rect 30156 21088 30162 21140
rect 30282 21088 30288 21140
rect 30340 21128 30346 21140
rect 32999 21131 33057 21137
rect 30340 21100 32720 21128
rect 30340 21088 30346 21100
rect 22094 21020 22100 21072
rect 22152 21060 22158 21072
rect 22152 21032 22508 21060
rect 22152 21020 22158 21032
rect 22020 20964 22140 20992
rect 18693 20927 18751 20933
rect 18693 20924 18705 20927
rect 18432 20896 18705 20924
rect 18432 20788 18460 20896
rect 18693 20893 18705 20896
rect 18739 20893 18751 20927
rect 18693 20887 18751 20893
rect 18785 20927 18843 20933
rect 18785 20893 18797 20927
rect 18831 20893 18843 20927
rect 18785 20887 18843 20893
rect 19061 20927 19119 20933
rect 19061 20893 19073 20927
rect 19107 20893 19119 20927
rect 21818 20924 21824 20936
rect 19061 20887 19119 20893
rect 20916 20896 21824 20924
rect 18509 20859 18567 20865
rect 18509 20825 18521 20859
rect 18555 20856 18567 20859
rect 19521 20859 19579 20865
rect 19521 20856 19533 20859
rect 18555 20828 19533 20856
rect 18555 20825 18567 20828
rect 18509 20819 18567 20825
rect 19521 20825 19533 20828
rect 19567 20825 19579 20859
rect 19521 20819 19579 20825
rect 19794 20816 19800 20868
rect 19852 20856 19858 20868
rect 19852 20828 20010 20856
rect 19852 20816 19858 20828
rect 20916 20788 20944 20896
rect 21818 20884 21824 20896
rect 21876 20924 21882 20936
rect 22112 20933 22140 20964
rect 22278 20952 22284 21004
rect 22336 20952 22342 21004
rect 22480 21001 22508 21032
rect 24118 21020 24124 21072
rect 24176 21060 24182 21072
rect 24176 21032 26004 21060
rect 24176 21020 24182 21032
rect 22465 20995 22523 21001
rect 22465 20961 22477 20995
rect 22511 20961 22523 20995
rect 22465 20955 22523 20961
rect 24213 20995 24271 21001
rect 24213 20961 24225 20995
rect 24259 20992 24271 20995
rect 24949 20995 25007 21001
rect 24949 20992 24961 20995
rect 24259 20964 24961 20992
rect 24259 20961 24271 20964
rect 24213 20955 24271 20961
rect 24949 20961 24961 20964
rect 24995 20992 25007 20995
rect 25498 20992 25504 21004
rect 24995 20964 25504 20992
rect 24995 20961 25007 20964
rect 24949 20955 25007 20961
rect 25498 20952 25504 20964
rect 25556 20992 25562 21004
rect 25556 20964 25728 20992
rect 25556 20952 25562 20964
rect 22005 20927 22063 20933
rect 22005 20924 22017 20927
rect 21876 20896 22017 20924
rect 21876 20884 21882 20896
rect 22005 20893 22017 20896
rect 22051 20893 22063 20927
rect 22005 20887 22063 20893
rect 22097 20927 22155 20933
rect 22097 20893 22109 20927
rect 22143 20893 22155 20927
rect 22097 20887 22155 20893
rect 22370 20884 22376 20936
rect 22428 20884 22434 20936
rect 24578 20884 24584 20936
rect 24636 20924 24642 20936
rect 25700 20933 25728 20964
rect 25317 20927 25375 20933
rect 25317 20924 25329 20927
rect 24636 20896 25329 20924
rect 24636 20884 24642 20896
rect 25317 20893 25329 20896
rect 25363 20893 25375 20927
rect 25317 20887 25375 20893
rect 25685 20927 25743 20933
rect 25685 20893 25697 20927
rect 25731 20893 25743 20927
rect 25976 20924 26004 21032
rect 26234 21020 26240 21072
rect 26292 21060 26298 21072
rect 26881 21063 26939 21069
rect 26881 21060 26893 21063
rect 26292 21032 26893 21060
rect 26292 21020 26298 21032
rect 26881 21029 26893 21032
rect 26927 21029 26939 21063
rect 26881 21023 26939 21029
rect 26050 20952 26056 21004
rect 26108 20992 26114 21004
rect 26108 20964 26464 20992
rect 26108 20952 26114 20964
rect 26436 20933 26464 20964
rect 26528 20964 26740 20992
rect 26191 20927 26249 20933
rect 26191 20924 26203 20927
rect 25976 20896 26203 20924
rect 25685 20887 25743 20893
rect 26191 20893 26203 20896
rect 26237 20893 26249 20927
rect 26191 20887 26249 20893
rect 26421 20927 26479 20933
rect 26421 20893 26433 20927
rect 26467 20893 26479 20927
rect 26421 20887 26479 20893
rect 22741 20859 22799 20865
rect 22741 20825 22753 20859
rect 22787 20825 22799 20859
rect 22741 20819 22799 20825
rect 18432 20760 20944 20788
rect 20990 20748 20996 20800
rect 21048 20748 21054 20800
rect 21821 20791 21879 20797
rect 21821 20757 21833 20791
rect 21867 20788 21879 20791
rect 22186 20788 22192 20800
rect 21867 20760 22192 20788
rect 21867 20757 21879 20760
rect 21821 20751 21879 20757
rect 22186 20748 22192 20760
rect 22244 20748 22250 20800
rect 22756 20788 22784 20819
rect 23198 20816 23204 20868
rect 23256 20816 23262 20868
rect 24118 20816 24124 20868
rect 24176 20856 24182 20868
rect 24397 20859 24455 20865
rect 24397 20856 24409 20859
rect 24176 20828 24409 20856
rect 24176 20816 24182 20828
rect 24397 20825 24409 20828
rect 24443 20825 24455 20859
rect 24397 20819 24455 20825
rect 24854 20816 24860 20868
rect 24912 20856 24918 20868
rect 25409 20859 25467 20865
rect 25409 20856 25421 20859
rect 24912 20828 25421 20856
rect 24912 20816 24918 20828
rect 25409 20825 25421 20828
rect 25455 20825 25467 20859
rect 25409 20819 25467 20825
rect 25501 20859 25559 20865
rect 25501 20825 25513 20859
rect 25547 20856 25559 20859
rect 25590 20856 25596 20868
rect 25547 20828 25596 20856
rect 25547 20825 25559 20828
rect 25501 20819 25559 20825
rect 25590 20816 25596 20828
rect 25648 20816 25654 20868
rect 25700 20856 25728 20887
rect 26329 20859 26387 20865
rect 26329 20856 26341 20859
rect 25700 20828 26341 20856
rect 26329 20825 26341 20828
rect 26375 20825 26387 20859
rect 26329 20819 26387 20825
rect 23658 20788 23664 20800
rect 22756 20760 23664 20788
rect 23658 20748 23664 20760
rect 23716 20748 23722 20800
rect 25866 20748 25872 20800
rect 25924 20788 25930 20800
rect 26528 20788 26556 20964
rect 26712 20933 26740 20964
rect 27522 20952 27528 21004
rect 27580 20992 27586 21004
rect 27580 20964 29408 20992
rect 27580 20952 27586 20964
rect 26604 20927 26662 20933
rect 26604 20893 26616 20927
rect 26650 20893 26662 20927
rect 26604 20887 26662 20893
rect 26697 20927 26755 20933
rect 26697 20893 26709 20927
rect 26743 20893 26755 20927
rect 26697 20887 26755 20893
rect 27065 20927 27123 20933
rect 27065 20893 27077 20927
rect 27111 20924 27123 20927
rect 27154 20924 27160 20936
rect 27111 20896 27160 20924
rect 27111 20893 27123 20896
rect 27065 20887 27123 20893
rect 26620 20856 26648 20887
rect 27154 20884 27160 20896
rect 27212 20884 27218 20936
rect 29380 20933 29408 20964
rect 30006 20952 30012 21004
rect 30064 20952 30070 21004
rect 31570 20952 31576 21004
rect 31628 20952 31634 21004
rect 32692 20992 32720 21100
rect 32999 21097 33011 21131
rect 33045 21128 33057 21131
rect 34146 21128 34152 21140
rect 33045 21100 34152 21128
rect 33045 21097 33057 21100
rect 32999 21091 33057 21097
rect 34146 21088 34152 21100
rect 34204 21088 34210 21140
rect 34422 21088 34428 21140
rect 34480 21128 34486 21140
rect 35158 21128 35164 21140
rect 34480 21100 35164 21128
rect 34480 21088 34486 21100
rect 35158 21088 35164 21100
rect 35216 21088 35222 21140
rect 35342 21088 35348 21140
rect 35400 21128 35406 21140
rect 35621 21131 35679 21137
rect 35621 21128 35633 21131
rect 35400 21100 35633 21128
rect 35400 21088 35406 21100
rect 35621 21097 35633 21100
rect 35667 21097 35679 21131
rect 35621 21091 35679 21097
rect 36265 21131 36323 21137
rect 36265 21097 36277 21131
rect 36311 21128 36323 21131
rect 36633 21131 36691 21137
rect 36633 21128 36645 21131
rect 36311 21100 36645 21128
rect 36311 21097 36323 21100
rect 36265 21091 36323 21097
rect 36633 21097 36645 21100
rect 36679 21128 36691 21131
rect 36722 21128 36728 21140
rect 36679 21100 36728 21128
rect 36679 21097 36691 21100
rect 36633 21091 36691 21097
rect 36722 21088 36728 21100
rect 36780 21088 36786 21140
rect 38654 21088 38660 21140
rect 38712 21128 38718 21140
rect 38712 21100 42196 21128
rect 38712 21088 38718 21100
rect 40586 21060 40592 21072
rect 39592 21032 40592 21060
rect 34330 20992 34336 21004
rect 32692 20964 34336 20992
rect 34330 20952 34336 20964
rect 34388 20952 34394 21004
rect 34698 20952 34704 21004
rect 34756 20952 34762 21004
rect 36262 20992 36268 21004
rect 35084 20964 36268 20992
rect 29365 20927 29423 20933
rect 29365 20893 29377 20927
rect 29411 20924 29423 20927
rect 29638 20924 29644 20936
rect 29411 20896 29644 20924
rect 29411 20893 29423 20896
rect 29365 20887 29423 20893
rect 29638 20884 29644 20896
rect 29696 20884 29702 20936
rect 29730 20884 29736 20936
rect 29788 20884 29794 20936
rect 29822 20884 29828 20936
rect 29880 20884 29886 20936
rect 30101 20927 30159 20933
rect 30101 20893 30113 20927
rect 30147 20924 30159 20927
rect 30469 20927 30527 20933
rect 30469 20924 30481 20927
rect 30147 20896 30481 20924
rect 30147 20893 30159 20896
rect 30101 20887 30159 20893
rect 30469 20893 30481 20896
rect 30515 20893 30527 20927
rect 30469 20887 30527 20893
rect 31021 20927 31079 20933
rect 31021 20893 31033 20927
rect 31067 20893 31079 20927
rect 31021 20887 31079 20893
rect 27798 20856 27804 20868
rect 26620 20828 27804 20856
rect 27798 20816 27804 20828
rect 27856 20816 27862 20868
rect 28626 20816 28632 20868
rect 28684 20816 28690 20868
rect 28810 20816 28816 20868
rect 28868 20856 28874 20868
rect 31036 20856 31064 20887
rect 31202 20884 31208 20936
rect 31260 20884 31266 20936
rect 31110 20856 31116 20868
rect 28868 20828 31116 20856
rect 28868 20816 28874 20828
rect 31110 20816 31116 20828
rect 31168 20816 31174 20868
rect 31938 20856 31944 20868
rect 31864 20828 31944 20856
rect 25924 20760 26556 20788
rect 27617 20791 27675 20797
rect 25924 20748 25930 20760
rect 27617 20757 27629 20791
rect 27663 20788 27675 20791
rect 27706 20788 27712 20800
rect 27663 20760 27712 20788
rect 27663 20757 27675 20760
rect 27617 20751 27675 20757
rect 27706 20748 27712 20760
rect 27764 20748 27770 20800
rect 29549 20791 29607 20797
rect 29549 20757 29561 20791
rect 29595 20788 29607 20791
rect 29914 20788 29920 20800
rect 29595 20760 29920 20788
rect 29595 20757 29607 20760
rect 29549 20751 29607 20757
rect 29914 20748 29920 20760
rect 29972 20748 29978 20800
rect 31294 20748 31300 20800
rect 31352 20788 31358 20800
rect 31864 20788 31892 20828
rect 31938 20816 31944 20828
rect 31996 20816 32002 20868
rect 34716 20856 34744 20952
rect 35084 20933 35112 20964
rect 36262 20952 36268 20964
rect 36320 20952 36326 21004
rect 36354 20952 36360 21004
rect 36412 20992 36418 21004
rect 39592 20992 39620 21032
rect 40586 21020 40592 21032
rect 40644 21060 40650 21072
rect 40862 21060 40868 21072
rect 40644 21032 40868 21060
rect 40644 21020 40650 21032
rect 40862 21020 40868 21032
rect 40920 21020 40926 21072
rect 42168 21060 42196 21100
rect 42886 21088 42892 21140
rect 42944 21128 42950 21140
rect 43165 21131 43223 21137
rect 43165 21128 43177 21131
rect 42944 21100 43177 21128
rect 42944 21088 42950 21100
rect 43165 21097 43177 21100
rect 43211 21128 43223 21131
rect 44082 21128 44088 21140
rect 43211 21100 44088 21128
rect 43211 21097 43223 21100
rect 43165 21091 43223 21097
rect 44082 21088 44088 21100
rect 44140 21088 44146 21140
rect 45002 21088 45008 21140
rect 45060 21088 45066 21140
rect 45462 21088 45468 21140
rect 45520 21128 45526 21140
rect 45649 21131 45707 21137
rect 45649 21128 45661 21131
rect 45520 21100 45661 21128
rect 45520 21088 45526 21100
rect 45649 21097 45661 21100
rect 45695 21097 45707 21131
rect 45649 21091 45707 21097
rect 47486 21088 47492 21140
rect 47544 21088 47550 21140
rect 47946 21088 47952 21140
rect 48004 21088 48010 21140
rect 48314 21088 48320 21140
rect 48372 21128 48378 21140
rect 49326 21128 49332 21140
rect 48372 21100 49332 21128
rect 48372 21088 48378 21100
rect 49326 21088 49332 21100
rect 49384 21128 49390 21140
rect 49789 21131 49847 21137
rect 49384 21100 49464 21128
rect 49384 21088 49390 21100
rect 43990 21060 43996 21072
rect 42168 21032 43996 21060
rect 43990 21020 43996 21032
rect 44048 21020 44054 21072
rect 44266 21060 44272 21072
rect 44100 21032 44272 21060
rect 36412 20964 39620 20992
rect 39669 20995 39727 21001
rect 36412 20952 36418 20964
rect 39669 20961 39681 20995
rect 39715 20992 39727 20995
rect 40034 20992 40040 21004
rect 39715 20964 40040 20992
rect 39715 20961 39727 20964
rect 39669 20955 39727 20961
rect 40034 20952 40040 20964
rect 40092 20992 40098 21004
rect 40405 20995 40463 21001
rect 40405 20992 40417 20995
rect 40092 20964 40417 20992
rect 40092 20952 40098 20964
rect 40405 20961 40417 20964
rect 40451 20961 40463 20995
rect 40405 20955 40463 20961
rect 41141 20995 41199 21001
rect 41141 20961 41153 20995
rect 41187 20992 41199 20995
rect 41690 20992 41696 21004
rect 41187 20964 41696 20992
rect 41187 20961 41199 20964
rect 41141 20955 41199 20961
rect 41690 20952 41696 20964
rect 41748 20952 41754 21004
rect 41874 20952 41880 21004
rect 41932 20992 41938 21004
rect 41932 20964 43116 20992
rect 41932 20952 41938 20964
rect 35069 20927 35127 20933
rect 35069 20893 35081 20927
rect 35115 20893 35127 20927
rect 35069 20887 35127 20893
rect 35158 20884 35164 20936
rect 35216 20924 35222 20936
rect 35345 20927 35403 20933
rect 35345 20924 35357 20927
rect 35216 20896 35357 20924
rect 35216 20884 35222 20896
rect 35345 20893 35357 20896
rect 35391 20893 35403 20927
rect 35345 20887 35403 20893
rect 35437 20927 35495 20933
rect 35437 20893 35449 20927
rect 35483 20924 35495 20927
rect 35802 20924 35808 20936
rect 35483 20896 35808 20924
rect 35483 20893 35495 20896
rect 35437 20887 35495 20893
rect 35802 20884 35808 20896
rect 35860 20884 35866 20936
rect 37918 20884 37924 20936
rect 37976 20884 37982 20936
rect 39298 20884 39304 20936
rect 39356 20884 39362 20936
rect 40494 20884 40500 20936
rect 40552 20924 40558 20936
rect 40865 20927 40923 20933
rect 40865 20924 40877 20927
rect 40552 20896 40877 20924
rect 40552 20884 40558 20896
rect 40865 20893 40877 20896
rect 40911 20893 40923 20927
rect 40865 20887 40923 20893
rect 42886 20884 42892 20936
rect 42944 20884 42950 20936
rect 35253 20859 35311 20865
rect 35253 20856 35265 20859
rect 34716 20828 35265 20856
rect 35253 20825 35265 20828
rect 35299 20825 35311 20859
rect 35253 20819 35311 20825
rect 36357 20859 36415 20865
rect 36357 20825 36369 20859
rect 36403 20856 36415 20859
rect 36814 20856 36820 20868
rect 36403 20828 36820 20856
rect 36403 20825 36415 20828
rect 36357 20819 36415 20825
rect 36814 20816 36820 20828
rect 36872 20816 36878 20868
rect 38194 20816 38200 20868
rect 38252 20816 38258 20868
rect 31352 20760 31892 20788
rect 31352 20748 31358 20760
rect 34514 20748 34520 20800
rect 34572 20788 34578 20800
rect 34698 20788 34704 20800
rect 34572 20760 34704 20788
rect 34572 20748 34578 20760
rect 34698 20748 34704 20760
rect 34756 20788 34762 20800
rect 34793 20791 34851 20797
rect 34793 20788 34805 20791
rect 34756 20760 34805 20788
rect 34756 20748 34762 20760
rect 34793 20757 34805 20760
rect 34839 20757 34851 20791
rect 34793 20751 34851 20757
rect 38470 20748 38476 20800
rect 38528 20788 38534 20800
rect 39316 20788 39344 20884
rect 42702 20856 42708 20868
rect 42366 20828 42708 20856
rect 42702 20816 42708 20828
rect 42760 20816 42766 20868
rect 38528 20760 39344 20788
rect 38528 20748 38534 20760
rect 39850 20748 39856 20800
rect 39908 20748 39914 20800
rect 42613 20791 42671 20797
rect 42613 20757 42625 20791
rect 42659 20788 42671 20791
rect 42978 20788 42984 20800
rect 42659 20760 42984 20788
rect 42659 20757 42671 20760
rect 42613 20751 42671 20757
rect 42978 20748 42984 20760
rect 43036 20748 43042 20800
rect 43088 20788 43116 20964
rect 44100 20933 44128 21032
rect 44266 21020 44272 21032
rect 44324 21020 44330 21072
rect 44729 21063 44787 21069
rect 44729 21029 44741 21063
rect 44775 21060 44787 21063
rect 47578 21060 47584 21072
rect 44775 21032 47584 21060
rect 44775 21029 44787 21032
rect 44729 21023 44787 21029
rect 47578 21020 47584 21032
rect 47636 21020 47642 21072
rect 48406 21060 48412 21072
rect 47688 21032 48412 21060
rect 46753 20995 46811 21001
rect 46753 20961 46765 20995
rect 46799 20992 46811 20995
rect 47688 20992 47716 21032
rect 48406 21020 48412 21032
rect 48464 21020 48470 21072
rect 48866 20992 48872 21004
rect 46799 20964 47716 20992
rect 48056 20964 48872 20992
rect 46799 20961 46811 20964
rect 46753 20955 46811 20961
rect 44266 20933 44272 20936
rect 44085 20927 44143 20933
rect 44085 20893 44097 20927
rect 44131 20893 44143 20927
rect 44085 20887 44143 20893
rect 44233 20927 44272 20933
rect 44233 20893 44245 20927
rect 44233 20887 44272 20893
rect 44266 20884 44272 20887
rect 44324 20884 44330 20936
rect 44450 20884 44456 20936
rect 44508 20884 44514 20936
rect 44634 20933 44640 20936
rect 44591 20927 44640 20933
rect 44591 20893 44603 20927
rect 44637 20893 44640 20927
rect 44591 20887 44640 20893
rect 44634 20884 44640 20887
rect 44692 20884 44698 20936
rect 44726 20884 44732 20936
rect 44784 20924 44790 20936
rect 45189 20927 45247 20933
rect 45189 20924 45201 20927
rect 44784 20896 45201 20924
rect 44784 20884 44790 20896
rect 45189 20893 45201 20896
rect 45235 20893 45247 20927
rect 45189 20887 45247 20893
rect 45278 20884 45284 20936
rect 45336 20884 45342 20936
rect 45557 20927 45615 20933
rect 45557 20893 45569 20927
rect 45603 20924 45615 20927
rect 46106 20924 46112 20936
rect 45603 20896 46112 20924
rect 45603 20893 45615 20896
rect 45557 20887 45615 20893
rect 46106 20884 46112 20896
rect 46164 20884 46170 20936
rect 46842 20884 46848 20936
rect 46900 20884 46906 20936
rect 47228 20933 47256 20964
rect 47121 20927 47179 20933
rect 47121 20924 47133 20927
rect 46951 20896 47133 20924
rect 44358 20816 44364 20868
rect 44416 20856 44422 20868
rect 44416 20828 44864 20856
rect 44416 20816 44422 20828
rect 44726 20788 44732 20800
rect 43088 20760 44732 20788
rect 44726 20748 44732 20760
rect 44784 20748 44790 20800
rect 44836 20788 44864 20828
rect 44910 20816 44916 20868
rect 44968 20856 44974 20868
rect 46951 20856 46979 20896
rect 47121 20893 47133 20896
rect 47167 20893 47179 20927
rect 47121 20887 47179 20893
rect 47213 20927 47271 20933
rect 47213 20893 47225 20927
rect 47259 20893 47271 20927
rect 47213 20887 47271 20893
rect 47486 20884 47492 20936
rect 47544 20924 47550 20936
rect 47670 20924 47676 20936
rect 47544 20896 47676 20924
rect 47544 20884 47550 20896
rect 47670 20884 47676 20896
rect 47728 20884 47734 20936
rect 47762 20884 47768 20936
rect 47820 20884 47826 20936
rect 48056 20933 48084 20964
rect 48866 20952 48872 20964
rect 48924 20952 48930 21004
rect 48590 20933 48596 20936
rect 48041 20927 48099 20933
rect 48041 20893 48053 20927
rect 48087 20893 48099 20927
rect 48588 20924 48596 20933
rect 48551 20896 48596 20924
rect 48041 20887 48099 20893
rect 48588 20887 48596 20896
rect 48590 20884 48596 20887
rect 48648 20884 48654 20936
rect 48682 20884 48688 20936
rect 48740 20884 48746 20936
rect 48774 20884 48780 20936
rect 48832 20884 48838 20936
rect 48958 20884 48964 20936
rect 49016 20884 49022 20936
rect 49050 20884 49056 20936
rect 49108 20884 49114 20936
rect 49142 20884 49148 20936
rect 49200 20884 49206 20936
rect 49326 20933 49332 20936
rect 49293 20927 49332 20933
rect 49293 20893 49305 20927
rect 49293 20887 49332 20893
rect 49326 20884 49332 20887
rect 49384 20884 49390 20936
rect 49436 20933 49464 21100
rect 49789 21097 49801 21131
rect 49835 21128 49847 21131
rect 50893 21131 50951 21137
rect 49835 21100 50845 21128
rect 49835 21097 49847 21100
rect 49789 21091 49847 21097
rect 49510 21020 49516 21072
rect 49568 21060 49574 21072
rect 50157 21063 50215 21069
rect 50157 21060 50169 21063
rect 49568 21032 50169 21060
rect 49568 21020 49574 21032
rect 50157 21029 50169 21032
rect 50203 21029 50215 21063
rect 50817 21060 50845 21100
rect 50893 21097 50905 21131
rect 50939 21128 50951 21131
rect 50982 21128 50988 21140
rect 50939 21100 50988 21128
rect 50939 21097 50951 21100
rect 50893 21091 50951 21097
rect 50982 21088 50988 21100
rect 51040 21088 51046 21140
rect 51258 21088 51264 21140
rect 51316 21128 51322 21140
rect 52178 21128 52184 21140
rect 51316 21100 52184 21128
rect 51316 21088 51322 21100
rect 52178 21088 52184 21100
rect 52236 21088 52242 21140
rect 52454 21088 52460 21140
rect 52512 21088 52518 21140
rect 50817 21032 51120 21060
rect 50157 21023 50215 21029
rect 49528 20964 50696 20992
rect 49528 20933 49556 20964
rect 49421 20927 49479 20933
rect 49421 20893 49433 20927
rect 49467 20893 49479 20927
rect 49421 20887 49479 20893
rect 49513 20927 49571 20933
rect 49513 20893 49525 20927
rect 49559 20893 49571 20927
rect 49513 20887 49571 20893
rect 49651 20927 49709 20933
rect 49651 20893 49663 20927
rect 49697 20924 49709 20927
rect 49786 20924 49792 20936
rect 49697 20896 49792 20924
rect 49697 20893 49709 20896
rect 49651 20887 49709 20893
rect 49786 20884 49792 20896
rect 49844 20884 49850 20936
rect 49970 20884 49976 20936
rect 50028 20924 50034 20936
rect 50295 20927 50353 20933
rect 50295 20924 50307 20927
rect 50028 20896 50307 20924
rect 50028 20884 50034 20896
rect 50295 20893 50307 20896
rect 50341 20893 50353 20927
rect 50295 20887 50353 20893
rect 50522 20884 50528 20936
rect 50580 20884 50586 20936
rect 50668 20933 50696 20964
rect 50653 20927 50711 20933
rect 50653 20893 50665 20927
rect 50699 20893 50711 20927
rect 50653 20887 50711 20893
rect 44968 20828 46979 20856
rect 47029 20859 47087 20865
rect 44968 20816 44974 20828
rect 47029 20825 47041 20859
rect 47075 20856 47087 20859
rect 47302 20856 47308 20868
rect 47075 20828 47308 20856
rect 47075 20825 47087 20828
rect 47029 20819 47087 20825
rect 45925 20791 45983 20797
rect 45925 20788 45937 20791
rect 44836 20760 45937 20788
rect 45925 20757 45937 20760
rect 45971 20788 45983 20791
rect 46290 20788 46296 20800
rect 45971 20760 46296 20788
rect 45971 20757 45983 20760
rect 45925 20751 45983 20757
rect 46290 20748 46296 20760
rect 46348 20748 46354 20800
rect 46569 20791 46627 20797
rect 46569 20757 46581 20791
rect 46615 20788 46627 20791
rect 47044 20788 47072 20819
rect 47302 20816 47308 20828
rect 47360 20816 47366 20868
rect 50154 20856 50160 20868
rect 47412 20828 50160 20856
rect 47412 20797 47440 20828
rect 50154 20816 50160 20828
rect 50212 20816 50218 20868
rect 50433 20859 50491 20865
rect 50433 20825 50445 20859
rect 50479 20825 50491 20859
rect 50668 20856 50696 20887
rect 50798 20884 50804 20936
rect 50856 20884 50862 20936
rect 51092 20933 51120 21032
rect 51350 20952 51356 21004
rect 51408 20952 51414 21004
rect 54478 20992 54484 21004
rect 51736 20964 54484 20992
rect 51077 20927 51135 20933
rect 51077 20893 51089 20927
rect 51123 20893 51135 20927
rect 51736 20924 51764 20964
rect 54478 20952 54484 20964
rect 54536 20952 54542 21004
rect 54938 20952 54944 21004
rect 54996 20992 55002 21004
rect 54996 20964 56088 20992
rect 54996 20952 55002 20964
rect 51077 20887 51135 20893
rect 51189 20896 51764 20924
rect 51813 20927 51871 20933
rect 51189 20856 51217 20896
rect 51813 20893 51825 20927
rect 51859 20893 51871 20927
rect 51813 20887 51871 20893
rect 50668 20828 51217 20856
rect 50433 20819 50491 20825
rect 46615 20760 47072 20788
rect 47397 20791 47455 20797
rect 46615 20757 46627 20760
rect 46569 20751 46627 20757
rect 47397 20757 47409 20791
rect 47443 20757 47455 20791
rect 47397 20751 47455 20757
rect 47486 20748 47492 20800
rect 47544 20788 47550 20800
rect 48133 20791 48191 20797
rect 48133 20788 48145 20791
rect 47544 20760 48145 20788
rect 47544 20748 47550 20760
rect 48133 20757 48145 20760
rect 48179 20757 48191 20791
rect 48133 20751 48191 20757
rect 48409 20791 48467 20797
rect 48409 20757 48421 20791
rect 48455 20788 48467 20791
rect 48866 20788 48872 20800
rect 48455 20760 48872 20788
rect 48455 20757 48467 20760
rect 48409 20751 48467 20757
rect 48866 20748 48872 20760
rect 48924 20748 48930 20800
rect 49234 20748 49240 20800
rect 49292 20788 49298 20800
rect 49786 20788 49792 20800
rect 49292 20760 49792 20788
rect 49292 20748 49298 20760
rect 49786 20748 49792 20760
rect 49844 20788 49850 20800
rect 49881 20791 49939 20797
rect 49881 20788 49893 20791
rect 49844 20760 49893 20788
rect 49844 20748 49850 20760
rect 49881 20757 49893 20760
rect 49927 20757 49939 20791
rect 49881 20751 49939 20757
rect 50246 20748 50252 20800
rect 50304 20788 50310 20800
rect 50448 20788 50476 20819
rect 51258 20816 51264 20868
rect 51316 20856 51322 20868
rect 51828 20856 51856 20887
rect 51902 20884 51908 20936
rect 51960 20924 51966 20936
rect 51960 20896 52005 20924
rect 51960 20884 51966 20896
rect 52086 20884 52092 20936
rect 52144 20884 52150 20936
rect 52178 20884 52184 20936
rect 52236 20884 52242 20936
rect 52319 20927 52377 20933
rect 52319 20893 52331 20927
rect 52365 20924 52377 20927
rect 52454 20924 52460 20936
rect 52365 20896 52460 20924
rect 52365 20893 52377 20896
rect 52319 20887 52377 20893
rect 52454 20884 52460 20896
rect 52512 20924 52518 20936
rect 52638 20924 52644 20936
rect 52512 20896 52644 20924
rect 52512 20884 52518 20896
rect 52638 20884 52644 20896
rect 52696 20884 52702 20936
rect 56060 20933 56088 20964
rect 56134 20952 56140 21004
rect 56192 20992 56198 21004
rect 58069 20995 58127 21001
rect 58069 20992 58081 20995
rect 56192 20964 58081 20992
rect 56192 20952 56198 20964
rect 58069 20961 58081 20964
rect 58115 20961 58127 20995
rect 58069 20955 58127 20961
rect 55677 20927 55735 20933
rect 55677 20924 55689 20927
rect 54404 20896 55689 20924
rect 52196 20856 52224 20884
rect 54404 20868 54432 20896
rect 55677 20893 55689 20896
rect 55723 20893 55735 20927
rect 55677 20887 55735 20893
rect 56045 20927 56103 20933
rect 56045 20893 56057 20927
rect 56091 20893 56103 20927
rect 56045 20887 56103 20893
rect 56686 20884 56692 20936
rect 56744 20884 56750 20936
rect 54386 20856 54392 20868
rect 51316 20828 51948 20856
rect 52196 20828 54392 20856
rect 51316 20816 51322 20828
rect 51810 20788 51816 20800
rect 50304 20760 51816 20788
rect 50304 20748 50310 20760
rect 51810 20748 51816 20760
rect 51868 20748 51874 20800
rect 51920 20788 51948 20828
rect 54386 20816 54392 20828
rect 54444 20816 54450 20868
rect 55122 20816 55128 20868
rect 55180 20856 55186 20868
rect 55861 20859 55919 20865
rect 55861 20856 55873 20859
rect 55180 20828 55873 20856
rect 55180 20816 55186 20828
rect 55861 20825 55873 20828
rect 55907 20825 55919 20859
rect 55861 20819 55919 20825
rect 55950 20816 55956 20868
rect 56008 20816 56014 20868
rect 57790 20816 57796 20868
rect 57848 20816 57854 20868
rect 53466 20788 53472 20800
rect 51920 20760 53472 20788
rect 53466 20748 53472 20760
rect 53524 20788 53530 20800
rect 54478 20788 54484 20800
rect 53524 20760 54484 20788
rect 53524 20748 53530 20760
rect 54478 20748 54484 20760
rect 54536 20748 54542 20800
rect 54754 20748 54760 20800
rect 54812 20788 54818 20800
rect 55033 20791 55091 20797
rect 55033 20788 55045 20791
rect 54812 20760 55045 20788
rect 54812 20748 54818 20760
rect 55033 20757 55045 20760
rect 55079 20788 55091 20791
rect 55582 20788 55588 20800
rect 55079 20760 55588 20788
rect 55079 20757 55091 20760
rect 55033 20751 55091 20757
rect 55582 20748 55588 20760
rect 55640 20788 55646 20800
rect 56042 20788 56048 20800
rect 55640 20760 56048 20788
rect 55640 20748 55646 20760
rect 56042 20748 56048 20760
rect 56100 20748 56106 20800
rect 56226 20748 56232 20800
rect 56284 20748 56290 20800
rect 56318 20748 56324 20800
rect 56376 20748 56382 20800
rect 1104 20698 58880 20720
rect 1104 20646 4874 20698
rect 4926 20646 4938 20698
rect 4990 20646 5002 20698
rect 5054 20646 5066 20698
rect 5118 20646 5130 20698
rect 5182 20646 35594 20698
rect 35646 20646 35658 20698
rect 35710 20646 35722 20698
rect 35774 20646 35786 20698
rect 35838 20646 35850 20698
rect 35902 20646 58880 20698
rect 1104 20624 58880 20646
rect 19150 20544 19156 20596
rect 19208 20544 19214 20596
rect 20441 20587 20499 20593
rect 20441 20584 20453 20587
rect 19904 20556 20453 20584
rect 19168 20516 19196 20544
rect 18524 20488 19196 20516
rect 18524 20457 18552 20488
rect 18509 20451 18567 20457
rect 18509 20417 18521 20451
rect 18555 20417 18567 20451
rect 18509 20411 18567 20417
rect 19794 20408 19800 20460
rect 19852 20448 19858 20460
rect 19904 20448 19932 20556
rect 20441 20553 20453 20556
rect 20487 20553 20499 20587
rect 20441 20547 20499 20553
rect 20530 20544 20536 20596
rect 20588 20584 20594 20596
rect 20588 20556 23612 20584
rect 20588 20544 20594 20556
rect 20346 20476 20352 20528
rect 20404 20516 20410 20528
rect 20717 20519 20775 20525
rect 20717 20516 20729 20519
rect 20404 20488 20729 20516
rect 20404 20476 20410 20488
rect 20717 20485 20729 20488
rect 20763 20516 20775 20519
rect 20901 20519 20959 20525
rect 20901 20516 20913 20519
rect 20763 20488 20913 20516
rect 20763 20485 20775 20488
rect 20717 20479 20775 20485
rect 20901 20485 20913 20488
rect 20947 20485 20959 20519
rect 22094 20516 22100 20528
rect 20901 20479 20959 20485
rect 21836 20488 22100 20516
rect 21836 20457 21864 20488
rect 22094 20476 22100 20488
rect 22152 20476 22158 20528
rect 22554 20476 22560 20528
rect 22612 20476 22618 20528
rect 23584 20516 23612 20556
rect 23658 20544 23664 20596
rect 23716 20544 23722 20596
rect 25133 20587 25191 20593
rect 25133 20553 25145 20587
rect 25179 20584 25191 20587
rect 25406 20584 25412 20596
rect 25179 20556 25412 20584
rect 25179 20553 25191 20556
rect 25133 20547 25191 20553
rect 24489 20519 24547 20525
rect 24489 20516 24501 20519
rect 23584 20488 24501 20516
rect 24489 20485 24501 20488
rect 24535 20485 24547 20519
rect 24489 20479 24547 20485
rect 19852 20434 19932 20448
rect 21821 20451 21879 20457
rect 19852 20420 19918 20434
rect 19852 20408 19858 20420
rect 21821 20417 21833 20451
rect 21867 20417 21879 20451
rect 21821 20411 21879 20417
rect 23842 20408 23848 20460
rect 23900 20408 23906 20460
rect 24026 20408 24032 20460
rect 24084 20408 24090 20460
rect 24118 20408 24124 20460
rect 24176 20408 24182 20460
rect 24213 20451 24271 20457
rect 24213 20417 24225 20451
rect 24259 20417 24271 20451
rect 24213 20411 24271 20417
rect 24397 20451 24455 20457
rect 24397 20417 24409 20451
rect 24443 20417 24455 20451
rect 24397 20411 24455 20417
rect 24581 20451 24639 20457
rect 24581 20417 24593 20451
rect 24627 20448 24639 20451
rect 25222 20448 25228 20460
rect 24627 20420 25228 20448
rect 24627 20417 24639 20420
rect 24581 20411 24639 20417
rect 18782 20340 18788 20392
rect 18840 20340 18846 20392
rect 20257 20383 20315 20389
rect 20257 20349 20269 20383
rect 20303 20380 20315 20383
rect 20438 20380 20444 20392
rect 20303 20352 20444 20380
rect 20303 20349 20315 20352
rect 20257 20343 20315 20349
rect 20438 20340 20444 20352
rect 20496 20340 20502 20392
rect 22097 20383 22155 20389
rect 22097 20349 22109 20383
rect 22143 20380 22155 20383
rect 22186 20380 22192 20392
rect 22143 20352 22192 20380
rect 22143 20349 22155 20352
rect 22097 20343 22155 20349
rect 22186 20340 22192 20352
rect 22244 20340 22250 20392
rect 23566 20340 23572 20392
rect 23624 20380 23630 20392
rect 24228 20380 24256 20411
rect 23624 20352 24256 20380
rect 24412 20380 24440 20411
rect 25222 20408 25228 20420
rect 25280 20408 25286 20460
rect 25130 20380 25136 20392
rect 24412 20352 25136 20380
rect 23624 20340 23630 20352
rect 25130 20340 25136 20352
rect 25188 20380 25194 20392
rect 25332 20380 25360 20556
rect 25406 20544 25412 20556
rect 25464 20544 25470 20596
rect 26421 20587 26479 20593
rect 26421 20584 26433 20587
rect 25700 20556 26433 20584
rect 25700 20525 25728 20556
rect 26421 20553 26433 20556
rect 26467 20584 26479 20587
rect 26694 20584 26700 20596
rect 26467 20556 26700 20584
rect 26467 20553 26479 20556
rect 26421 20547 26479 20553
rect 26694 20544 26700 20556
rect 26752 20584 26758 20596
rect 27338 20584 27344 20596
rect 26752 20556 27344 20584
rect 26752 20544 26758 20556
rect 27338 20544 27344 20556
rect 27396 20544 27402 20596
rect 28813 20587 28871 20593
rect 28460 20556 28672 20584
rect 25685 20519 25743 20525
rect 25685 20485 25697 20519
rect 25731 20485 25743 20519
rect 25685 20479 25743 20485
rect 26326 20476 26332 20528
rect 26384 20516 26390 20528
rect 26970 20516 26976 20528
rect 26384 20488 26976 20516
rect 26384 20476 26390 20488
rect 26970 20476 26976 20488
rect 27028 20516 27034 20528
rect 28460 20525 28488 20556
rect 28445 20519 28503 20525
rect 28445 20516 28457 20519
rect 27028 20488 28457 20516
rect 27028 20476 27034 20488
rect 28445 20485 28457 20488
rect 28491 20485 28503 20519
rect 28445 20479 28503 20485
rect 28534 20476 28540 20528
rect 28592 20476 28598 20528
rect 28644 20516 28672 20556
rect 28813 20553 28825 20587
rect 28859 20584 28871 20587
rect 29822 20584 29828 20596
rect 28859 20556 29828 20584
rect 28859 20553 28871 20556
rect 28813 20547 28871 20553
rect 29822 20544 29828 20556
rect 29880 20544 29886 20596
rect 30926 20544 30932 20596
rect 30984 20584 30990 20596
rect 30984 20556 34284 20584
rect 30984 20544 30990 20556
rect 28644 20488 29224 20516
rect 25406 20408 25412 20460
rect 25464 20408 25470 20460
rect 25498 20408 25504 20460
rect 25556 20448 25562 20460
rect 25777 20451 25835 20457
rect 25556 20420 25601 20448
rect 25556 20408 25562 20420
rect 25777 20417 25789 20451
rect 25823 20417 25835 20451
rect 25777 20411 25835 20417
rect 25915 20451 25973 20457
rect 25915 20417 25927 20451
rect 25961 20448 25973 20451
rect 26142 20448 26148 20460
rect 25961 20420 26148 20448
rect 25961 20417 25973 20420
rect 25915 20411 25973 20417
rect 25188 20352 25360 20380
rect 25188 20340 25194 20352
rect 25792 20312 25820 20411
rect 26142 20408 26148 20420
rect 26200 20408 26206 20460
rect 27706 20408 27712 20460
rect 27764 20448 27770 20460
rect 28261 20451 28319 20457
rect 28261 20448 28273 20451
rect 27764 20420 28273 20448
rect 27764 20408 27770 20420
rect 28261 20417 28273 20420
rect 28307 20417 28319 20451
rect 28261 20411 28319 20417
rect 28629 20451 28687 20457
rect 28629 20417 28641 20451
rect 28675 20448 28687 20451
rect 28718 20448 28724 20460
rect 28675 20420 28724 20448
rect 28675 20417 28687 20420
rect 28629 20411 28687 20417
rect 28718 20408 28724 20420
rect 28776 20408 28782 20460
rect 29086 20408 29092 20460
rect 29144 20408 29150 20460
rect 29196 20448 29224 20488
rect 29270 20476 29276 20528
rect 29328 20476 29334 20528
rect 29914 20476 29920 20528
rect 29972 20476 29978 20528
rect 31294 20516 31300 20528
rect 31142 20488 31300 20516
rect 31294 20476 31300 20488
rect 31352 20476 31358 20528
rect 34256 20516 34284 20556
rect 34790 20544 34796 20596
rect 34848 20584 34854 20596
rect 34848 20556 35848 20584
rect 34848 20544 34854 20556
rect 34256 20488 34362 20516
rect 35268 20488 35664 20516
rect 29362 20448 29368 20460
rect 29196 20420 29368 20448
rect 29362 20408 29368 20420
rect 29420 20408 29426 20460
rect 34790 20408 34796 20460
rect 34848 20448 34854 20460
rect 35268 20448 35296 20488
rect 34848 20420 35296 20448
rect 34848 20408 34854 20420
rect 27798 20340 27804 20392
rect 27856 20380 27862 20392
rect 28810 20380 28816 20392
rect 27856 20352 28816 20380
rect 27856 20340 27862 20352
rect 28810 20340 28816 20352
rect 28868 20380 28874 20392
rect 28905 20383 28963 20389
rect 28905 20380 28917 20383
rect 28868 20352 28917 20380
rect 28868 20340 28874 20352
rect 28905 20349 28917 20352
rect 28951 20349 28963 20383
rect 28905 20343 28963 20349
rect 29638 20340 29644 20392
rect 29696 20340 29702 20392
rect 30926 20380 30932 20392
rect 29748 20352 30932 20380
rect 26510 20312 26516 20324
rect 23492 20284 25820 20312
rect 25884 20284 26516 20312
rect 19518 20204 19524 20256
rect 19576 20244 19582 20256
rect 23492 20244 23520 20284
rect 19576 20216 23520 20244
rect 19576 20204 19582 20216
rect 24762 20204 24768 20256
rect 24820 20204 24826 20256
rect 24949 20247 25007 20253
rect 24949 20213 24961 20247
rect 24995 20244 25007 20247
rect 25222 20244 25228 20256
rect 24995 20216 25228 20244
rect 24995 20213 25007 20216
rect 24949 20207 25007 20213
rect 25222 20204 25228 20216
rect 25280 20244 25286 20256
rect 25590 20244 25596 20256
rect 25280 20216 25596 20244
rect 25280 20204 25286 20216
rect 25590 20204 25596 20216
rect 25648 20244 25654 20256
rect 25884 20244 25912 20284
rect 26510 20272 26516 20284
rect 26568 20272 26574 20324
rect 28626 20272 28632 20324
rect 28684 20312 28690 20324
rect 29748 20312 29776 20352
rect 30926 20340 30932 20352
rect 30984 20340 30990 20392
rect 31110 20340 31116 20392
rect 31168 20380 31174 20392
rect 31386 20380 31392 20392
rect 31168 20352 31392 20380
rect 31168 20340 31174 20352
rect 31386 20340 31392 20352
rect 31444 20340 31450 20392
rect 33594 20340 33600 20392
rect 33652 20340 33658 20392
rect 33965 20383 34023 20389
rect 33965 20349 33977 20383
rect 34011 20380 34023 20383
rect 34698 20380 34704 20392
rect 34011 20352 34704 20380
rect 34011 20349 34023 20352
rect 33965 20343 34023 20349
rect 34698 20340 34704 20352
rect 34756 20340 34762 20392
rect 35158 20340 35164 20392
rect 35216 20380 35222 20392
rect 35342 20380 35348 20392
rect 35216 20352 35348 20380
rect 35216 20340 35222 20352
rect 35342 20340 35348 20352
rect 35400 20389 35406 20392
rect 35400 20383 35449 20389
rect 35400 20349 35403 20383
rect 35437 20349 35449 20383
rect 35400 20343 35449 20349
rect 35529 20383 35587 20389
rect 35529 20349 35541 20383
rect 35575 20349 35587 20383
rect 35636 20380 35664 20488
rect 35710 20408 35716 20460
rect 35768 20448 35774 20460
rect 35820 20457 35848 20556
rect 36446 20544 36452 20596
rect 36504 20584 36510 20596
rect 36633 20587 36691 20593
rect 36633 20584 36645 20587
rect 36504 20556 36645 20584
rect 36504 20544 36510 20556
rect 36633 20553 36645 20556
rect 36679 20553 36691 20587
rect 36633 20547 36691 20553
rect 38194 20544 38200 20596
rect 38252 20584 38258 20596
rect 38473 20587 38531 20593
rect 38473 20584 38485 20587
rect 38252 20556 38485 20584
rect 38252 20544 38258 20556
rect 38473 20553 38485 20556
rect 38519 20553 38531 20587
rect 39022 20584 39028 20596
rect 38473 20547 38531 20553
rect 38580 20556 39028 20584
rect 35805 20451 35863 20457
rect 35805 20448 35817 20451
rect 35768 20420 35817 20448
rect 35768 20408 35774 20420
rect 35805 20417 35817 20420
rect 35851 20417 35863 20451
rect 35805 20411 35863 20417
rect 36262 20408 36268 20460
rect 36320 20448 36326 20460
rect 36449 20451 36507 20457
rect 36449 20448 36461 20451
rect 36320 20420 36461 20448
rect 36320 20408 36326 20420
rect 36449 20417 36461 20420
rect 36495 20417 36507 20451
rect 36449 20411 36507 20417
rect 38580 20380 38608 20556
rect 39022 20544 39028 20556
rect 39080 20584 39086 20596
rect 40218 20584 40224 20596
rect 39080 20556 40224 20584
rect 39080 20544 39086 20556
rect 40218 20544 40224 20556
rect 40276 20544 40282 20596
rect 42610 20584 42616 20596
rect 40512 20556 42616 20584
rect 39117 20519 39175 20525
rect 39117 20516 39129 20519
rect 38764 20488 39129 20516
rect 38764 20457 38792 20488
rect 39117 20485 39129 20488
rect 39163 20485 39175 20519
rect 39850 20516 39856 20528
rect 39117 20479 39175 20485
rect 39224 20488 39856 20516
rect 38657 20451 38715 20457
rect 38657 20417 38669 20451
rect 38703 20417 38715 20451
rect 38657 20411 38715 20417
rect 38749 20451 38807 20457
rect 38749 20417 38761 20451
rect 38795 20417 38807 20451
rect 38749 20411 38807 20417
rect 39025 20451 39083 20457
rect 39025 20417 39037 20451
rect 39071 20448 39083 20451
rect 39224 20448 39252 20488
rect 39850 20476 39856 20488
rect 39908 20476 39914 20528
rect 39071 20420 39252 20448
rect 39071 20417 39083 20420
rect 39025 20411 39083 20417
rect 35636 20352 38608 20380
rect 38672 20380 38700 20411
rect 39298 20408 39304 20460
rect 39356 20448 39362 20460
rect 40512 20448 40540 20556
rect 42610 20544 42616 20556
rect 42668 20544 42674 20596
rect 42702 20544 42708 20596
rect 42760 20544 42766 20596
rect 43070 20544 43076 20596
rect 43128 20544 43134 20596
rect 43162 20544 43168 20596
rect 43220 20584 43226 20596
rect 44266 20584 44272 20596
rect 43220 20556 44272 20584
rect 43220 20544 43226 20556
rect 42720 20516 42748 20544
rect 41998 20488 42748 20516
rect 42794 20476 42800 20528
rect 42852 20476 42858 20528
rect 39356 20420 40540 20448
rect 39356 20408 39362 20420
rect 42610 20408 42616 20460
rect 42668 20408 42674 20460
rect 42705 20451 42763 20457
rect 42705 20417 42717 20451
rect 42751 20448 42763 20451
rect 42886 20448 42892 20460
rect 42751 20420 42892 20448
rect 42751 20417 42763 20420
rect 42705 20411 42763 20417
rect 42886 20408 42892 20420
rect 42944 20408 42950 20460
rect 42978 20408 42984 20460
rect 43036 20408 43042 20460
rect 43364 20457 43392 20556
rect 44266 20544 44272 20556
rect 44324 20544 44330 20596
rect 45094 20584 45100 20596
rect 45020 20556 45100 20584
rect 44910 20476 44916 20528
rect 44968 20476 44974 20528
rect 45020 20525 45048 20556
rect 45094 20544 45100 20556
rect 45152 20584 45158 20596
rect 45373 20587 45431 20593
rect 45373 20584 45385 20587
rect 45152 20556 45385 20584
rect 45152 20544 45158 20556
rect 45373 20553 45385 20556
rect 45419 20553 45431 20587
rect 45373 20547 45431 20553
rect 47118 20544 47124 20596
rect 47176 20544 47182 20596
rect 47305 20587 47363 20593
rect 47305 20553 47317 20587
rect 47351 20584 47363 20587
rect 47854 20584 47860 20596
rect 47351 20556 47860 20584
rect 47351 20553 47363 20556
rect 47305 20547 47363 20553
rect 47854 20544 47860 20556
rect 47912 20544 47918 20596
rect 48038 20544 48044 20596
rect 48096 20584 48102 20596
rect 48222 20584 48228 20596
rect 48096 20556 48228 20584
rect 48096 20544 48102 20556
rect 48222 20544 48228 20556
rect 48280 20544 48286 20596
rect 48866 20544 48872 20596
rect 48924 20584 48930 20596
rect 49326 20584 49332 20596
rect 48924 20556 49332 20584
rect 48924 20544 48930 20556
rect 49326 20544 49332 20556
rect 49384 20544 49390 20596
rect 49602 20544 49608 20596
rect 49660 20544 49666 20596
rect 56318 20584 56324 20596
rect 56244 20556 56324 20584
rect 45005 20519 45063 20525
rect 45005 20485 45017 20519
rect 45051 20485 45063 20519
rect 46750 20516 46756 20528
rect 45005 20479 45063 20485
rect 45204 20488 46756 20516
rect 43257 20451 43315 20457
rect 43257 20417 43269 20451
rect 43303 20417 43315 20451
rect 43257 20411 43315 20417
rect 43349 20451 43407 20457
rect 43349 20417 43361 20451
rect 43395 20417 43407 20451
rect 43349 20411 43407 20417
rect 43441 20451 43499 20457
rect 43441 20417 43453 20451
rect 43487 20448 43499 20451
rect 43530 20448 43536 20460
rect 43487 20420 43536 20448
rect 43487 20417 43499 20420
rect 43441 20411 43499 20417
rect 39114 20380 39120 20392
rect 38672 20352 39120 20380
rect 35529 20343 35587 20349
rect 35400 20340 35406 20343
rect 28684 20284 29776 20312
rect 28684 20272 28690 20284
rect 25648 20216 25912 20244
rect 25648 20204 25654 20216
rect 26050 20204 26056 20256
rect 26108 20204 26114 20256
rect 26602 20204 26608 20256
rect 26660 20244 26666 20256
rect 27062 20244 27068 20256
rect 26660 20216 27068 20244
rect 26660 20204 26666 20216
rect 27062 20204 27068 20216
rect 27120 20204 27126 20256
rect 29362 20204 29368 20256
rect 29420 20244 29426 20256
rect 35543 20244 35571 20343
rect 39114 20340 39120 20352
rect 39172 20340 39178 20392
rect 39482 20340 39488 20392
rect 39540 20340 39546 20392
rect 40494 20340 40500 20392
rect 40552 20340 40558 20392
rect 40773 20383 40831 20389
rect 40773 20349 40785 20383
rect 40819 20380 40831 20383
rect 41322 20380 41328 20392
rect 40819 20352 41328 20380
rect 40819 20349 40831 20352
rect 40773 20343 40831 20349
rect 41322 20340 41328 20352
rect 41380 20340 41386 20392
rect 42628 20380 42656 20408
rect 43272 20380 43300 20411
rect 43530 20408 43536 20420
rect 43588 20408 43594 20460
rect 43625 20451 43683 20457
rect 43625 20417 43637 20451
rect 43671 20448 43683 20451
rect 44358 20448 44364 20460
rect 43671 20420 44364 20448
rect 43671 20417 43683 20420
rect 43625 20411 43683 20417
rect 44358 20408 44364 20420
rect 44416 20408 44422 20460
rect 44818 20457 44824 20460
rect 44775 20451 44824 20457
rect 44775 20417 44787 20451
rect 44821 20417 44824 20451
rect 44775 20411 44824 20417
rect 44790 20408 44824 20411
rect 44876 20408 44882 20460
rect 45204 20457 45232 20488
rect 46750 20476 46756 20488
rect 46808 20516 46814 20528
rect 47949 20519 48007 20525
rect 47949 20516 47961 20519
rect 46808 20488 47961 20516
rect 46808 20476 46814 20488
rect 47949 20485 47961 20488
rect 47995 20516 48007 20519
rect 48593 20519 48651 20525
rect 47995 20488 48176 20516
rect 47995 20485 48007 20488
rect 47949 20479 48007 20485
rect 45188 20451 45246 20457
rect 45188 20417 45200 20451
rect 45234 20417 45246 20451
rect 45188 20411 45246 20417
rect 45281 20451 45339 20457
rect 45281 20417 45293 20451
rect 45327 20417 45339 20451
rect 45281 20411 45339 20417
rect 44790 20380 44818 20408
rect 42628 20352 44818 20380
rect 41874 20272 41880 20324
rect 41932 20312 41938 20324
rect 42245 20315 42303 20321
rect 42245 20312 42257 20315
rect 41932 20284 42257 20312
rect 41932 20272 41938 20284
rect 42245 20281 42257 20284
rect 42291 20312 42303 20315
rect 43162 20312 43168 20324
rect 42291 20284 43168 20312
rect 42291 20281 42303 20284
rect 42245 20275 42303 20281
rect 43162 20272 43168 20284
rect 43220 20272 43226 20324
rect 44545 20315 44603 20321
rect 44545 20281 44557 20315
rect 44591 20312 44603 20315
rect 45296 20312 45324 20411
rect 47578 20408 47584 20460
rect 47636 20408 47642 20460
rect 47762 20457 47768 20460
rect 47729 20451 47768 20457
rect 47729 20417 47741 20451
rect 47729 20411 47768 20417
rect 47762 20408 47768 20411
rect 47820 20408 47826 20460
rect 47854 20408 47860 20460
rect 47912 20408 47918 20460
rect 48046 20451 48104 20457
rect 48046 20448 48058 20451
rect 47964 20420 48058 20448
rect 47118 20340 47124 20392
rect 47176 20380 47182 20392
rect 47964 20380 47992 20420
rect 48046 20417 48058 20420
rect 48092 20417 48104 20451
rect 48046 20411 48104 20417
rect 48148 20392 48176 20488
rect 48240 20488 48544 20516
rect 47176 20352 47992 20380
rect 47176 20340 47182 20352
rect 47688 20324 47716 20352
rect 48130 20340 48136 20392
rect 48188 20340 48194 20392
rect 45646 20312 45652 20324
rect 44591 20284 45652 20312
rect 44591 20281 44603 20284
rect 44545 20275 44603 20281
rect 45646 20272 45652 20284
rect 45704 20312 45710 20324
rect 47026 20312 47032 20324
rect 45704 20284 47032 20312
rect 45704 20272 45710 20284
rect 47026 20272 47032 20284
rect 47084 20272 47090 20324
rect 47670 20272 47676 20324
rect 47728 20272 47734 20324
rect 48240 20321 48268 20488
rect 48317 20451 48375 20457
rect 48317 20417 48329 20451
rect 48363 20417 48375 20451
rect 48317 20411 48375 20417
rect 48410 20451 48468 20457
rect 48410 20417 48422 20451
rect 48456 20417 48468 20451
rect 48516 20448 48544 20488
rect 48593 20485 48605 20519
rect 48639 20516 48651 20519
rect 49620 20516 49648 20544
rect 48639 20488 49648 20516
rect 48639 20485 48651 20488
rect 48593 20479 48651 20485
rect 49878 20476 49884 20528
rect 49936 20476 49942 20528
rect 49970 20476 49976 20528
rect 50028 20516 50034 20528
rect 50157 20519 50215 20525
rect 50157 20516 50169 20519
rect 50028 20488 50169 20516
rect 50028 20476 50034 20488
rect 50157 20485 50169 20488
rect 50203 20485 50215 20519
rect 50157 20479 50215 20485
rect 52454 20476 52460 20528
rect 52512 20516 52518 20528
rect 52512 20488 53972 20516
rect 52512 20476 52518 20488
rect 48516 20420 48636 20448
rect 48410 20411 48468 20417
rect 48332 20324 48360 20411
rect 48225 20315 48283 20321
rect 48225 20281 48237 20315
rect 48271 20281 48283 20315
rect 48225 20275 48283 20281
rect 48314 20272 48320 20324
rect 48372 20272 48378 20324
rect 48424 20312 48452 20411
rect 48608 20380 48636 20420
rect 48682 20408 48688 20460
rect 48740 20408 48746 20460
rect 48774 20408 48780 20460
rect 48832 20457 48838 20460
rect 48832 20451 48859 20457
rect 48847 20417 48859 20451
rect 48832 20411 48859 20417
rect 49053 20451 49111 20457
rect 49053 20417 49065 20451
rect 49099 20417 49111 20451
rect 49053 20411 49111 20417
rect 48832 20408 48838 20411
rect 49068 20380 49096 20411
rect 49326 20408 49332 20460
rect 49384 20408 49390 20460
rect 50062 20408 50068 20460
rect 50120 20448 50126 20460
rect 50522 20448 50528 20460
rect 50120 20420 50528 20448
rect 50120 20408 50126 20420
rect 50522 20408 50528 20420
rect 50580 20408 50586 20460
rect 53653 20451 53711 20457
rect 53653 20417 53665 20451
rect 53699 20448 53711 20451
rect 53834 20448 53840 20460
rect 53699 20420 53840 20448
rect 53699 20417 53711 20420
rect 53653 20411 53711 20417
rect 53834 20408 53840 20420
rect 53892 20408 53898 20460
rect 53944 20448 53972 20488
rect 54570 20476 54576 20528
rect 54628 20516 54634 20528
rect 56244 20516 56272 20556
rect 56318 20544 56324 20556
rect 56376 20544 56382 20596
rect 56781 20587 56839 20593
rect 56781 20553 56793 20587
rect 56827 20584 56839 20587
rect 57790 20584 57796 20596
rect 56827 20556 57796 20584
rect 56827 20553 56839 20556
rect 56781 20547 56839 20553
rect 57790 20544 57796 20556
rect 57848 20544 57854 20596
rect 54628 20488 56272 20516
rect 54628 20476 54634 20488
rect 54938 20448 54944 20460
rect 53944 20420 54944 20448
rect 54938 20408 54944 20420
rect 54996 20408 55002 20460
rect 55398 20408 55404 20460
rect 55456 20408 55462 20460
rect 56244 20457 56272 20488
rect 56229 20451 56287 20457
rect 56229 20417 56241 20451
rect 56275 20417 56287 20451
rect 56229 20411 56287 20417
rect 56318 20408 56324 20460
rect 56376 20448 56382 20460
rect 56505 20451 56563 20457
rect 56505 20448 56517 20451
rect 56376 20420 56517 20448
rect 56376 20408 56382 20420
rect 56505 20417 56517 20420
rect 56551 20417 56563 20451
rect 56505 20411 56563 20417
rect 56597 20451 56655 20457
rect 56597 20417 56609 20451
rect 56643 20417 56655 20451
rect 56597 20411 56655 20417
rect 48608 20352 49096 20380
rect 49237 20383 49295 20389
rect 49237 20349 49249 20383
rect 49283 20380 49295 20383
rect 49418 20380 49424 20392
rect 49283 20352 49424 20380
rect 49283 20349 49295 20352
rect 49237 20343 49295 20349
rect 49418 20340 49424 20352
rect 49476 20340 49482 20392
rect 50890 20340 50896 20392
rect 50948 20380 50954 20392
rect 53929 20383 53987 20389
rect 53929 20380 53941 20383
rect 50948 20352 53941 20380
rect 50948 20340 50954 20352
rect 53929 20349 53941 20352
rect 53975 20380 53987 20383
rect 54846 20380 54852 20392
rect 53975 20352 54852 20380
rect 53975 20349 53987 20352
rect 53929 20343 53987 20349
rect 54846 20340 54852 20352
rect 54904 20340 54910 20392
rect 55125 20383 55183 20389
rect 55125 20349 55137 20383
rect 55171 20380 55183 20383
rect 55950 20380 55956 20392
rect 55171 20352 55956 20380
rect 55171 20349 55183 20352
rect 55125 20343 55183 20349
rect 48590 20312 48596 20324
rect 48424 20284 48596 20312
rect 48590 20272 48596 20284
rect 48648 20272 48654 20324
rect 48866 20312 48872 20324
rect 48797 20284 48872 20312
rect 36817 20247 36875 20253
rect 36817 20244 36829 20247
rect 29420 20216 36829 20244
rect 29420 20204 29426 20216
rect 36817 20213 36829 20216
rect 36863 20244 36875 20247
rect 37182 20244 37188 20256
rect 36863 20216 37188 20244
rect 36863 20213 36875 20216
rect 36817 20207 36875 20213
rect 37182 20204 37188 20216
rect 37240 20204 37246 20256
rect 38933 20247 38991 20253
rect 38933 20213 38945 20247
rect 38979 20244 38991 20247
rect 39669 20247 39727 20253
rect 39669 20244 39681 20247
rect 38979 20216 39681 20244
rect 38979 20213 38991 20216
rect 38933 20207 38991 20213
rect 39669 20213 39681 20216
rect 39715 20244 39727 20247
rect 41230 20244 41236 20256
rect 39715 20216 41236 20244
rect 39715 20213 39727 20216
rect 39669 20207 39727 20213
rect 41230 20204 41236 20216
rect 41288 20204 41294 20256
rect 42426 20204 42432 20256
rect 42484 20204 42490 20256
rect 42794 20204 42800 20256
rect 42852 20244 42858 20256
rect 43530 20244 43536 20256
rect 42852 20216 43536 20244
rect 42852 20204 42858 20216
rect 43530 20204 43536 20216
rect 43588 20204 43594 20256
rect 44637 20247 44695 20253
rect 44637 20213 44649 20247
rect 44683 20244 44695 20247
rect 45186 20244 45192 20256
rect 44683 20216 45192 20244
rect 44683 20213 44695 20216
rect 44637 20207 44695 20213
rect 45186 20204 45192 20216
rect 45244 20204 45250 20256
rect 45554 20204 45560 20256
rect 45612 20204 45618 20256
rect 47762 20204 47768 20256
rect 47820 20244 47826 20256
rect 48797 20244 48825 20284
rect 48866 20272 48872 20284
rect 48924 20272 48930 20324
rect 49510 20272 49516 20324
rect 49568 20272 49574 20324
rect 53374 20272 53380 20324
rect 53432 20312 53438 20324
rect 55140 20312 55168 20343
rect 55950 20340 55956 20352
rect 56008 20340 56014 20392
rect 53432 20284 55168 20312
rect 53432 20272 53438 20284
rect 55306 20272 55312 20324
rect 55364 20312 55370 20324
rect 56321 20315 56379 20321
rect 56321 20312 56333 20315
rect 55364 20284 56333 20312
rect 55364 20272 55370 20284
rect 56321 20281 56333 20284
rect 56367 20281 56379 20315
rect 56321 20275 56379 20281
rect 47820 20216 48825 20244
rect 48961 20247 49019 20253
rect 47820 20204 47826 20216
rect 48961 20213 48973 20247
rect 49007 20244 49019 20247
rect 49053 20247 49111 20253
rect 49053 20244 49065 20247
rect 49007 20216 49065 20244
rect 49007 20213 49019 20216
rect 48961 20207 49019 20213
rect 49053 20213 49065 20216
rect 49099 20213 49111 20247
rect 49053 20207 49111 20213
rect 50430 20204 50436 20256
rect 50488 20244 50494 20256
rect 53101 20247 53159 20253
rect 53101 20244 53113 20247
rect 50488 20216 53113 20244
rect 50488 20204 50494 20216
rect 53101 20213 53113 20216
rect 53147 20244 53159 20247
rect 53282 20244 53288 20256
rect 53147 20216 53288 20244
rect 53147 20213 53159 20216
rect 53101 20207 53159 20213
rect 53282 20204 53288 20216
rect 53340 20204 53346 20256
rect 53469 20247 53527 20253
rect 53469 20213 53481 20247
rect 53515 20244 53527 20247
rect 53650 20244 53656 20256
rect 53515 20216 53656 20244
rect 53515 20213 53527 20216
rect 53469 20207 53527 20213
rect 53650 20204 53656 20216
rect 53708 20204 53714 20256
rect 53837 20247 53895 20253
rect 53837 20213 53849 20247
rect 53883 20244 53895 20247
rect 53926 20244 53932 20256
rect 53883 20216 53932 20244
rect 53883 20213 53895 20216
rect 53837 20207 53895 20213
rect 53926 20204 53932 20216
rect 53984 20204 53990 20256
rect 55214 20204 55220 20256
rect 55272 20204 55278 20256
rect 55582 20204 55588 20256
rect 55640 20204 55646 20256
rect 56042 20204 56048 20256
rect 56100 20244 56106 20256
rect 56612 20244 56640 20411
rect 56100 20216 56640 20244
rect 56100 20204 56106 20216
rect 1104 20154 58880 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 58880 20154
rect 1104 20080 58880 20102
rect 25406 20000 25412 20052
rect 25464 20000 25470 20052
rect 25593 20043 25651 20049
rect 25593 20009 25605 20043
rect 25639 20040 25651 20043
rect 25682 20040 25688 20052
rect 25639 20012 25688 20040
rect 25639 20009 25651 20012
rect 25593 20003 25651 20009
rect 25682 20000 25688 20012
rect 25740 20000 25746 20052
rect 26050 20000 26056 20052
rect 26108 20040 26114 20052
rect 26605 20043 26663 20049
rect 26605 20040 26617 20043
rect 26108 20012 26617 20040
rect 26108 20000 26114 20012
rect 26605 20009 26617 20012
rect 26651 20009 26663 20043
rect 26605 20003 26663 20009
rect 27062 20000 27068 20052
rect 27120 20040 27126 20052
rect 27341 20043 27399 20049
rect 27341 20040 27353 20043
rect 27120 20012 27353 20040
rect 27120 20000 27126 20012
rect 27341 20009 27353 20012
rect 27387 20040 27399 20043
rect 29178 20040 29184 20052
rect 27387 20012 29184 20040
rect 27387 20009 27399 20012
rect 27341 20003 27399 20009
rect 29178 20000 29184 20012
rect 29236 20000 29242 20052
rect 33965 20043 34023 20049
rect 30760 20012 31754 20040
rect 22646 19932 22652 19984
rect 22704 19972 22710 19984
rect 26418 19972 26424 19984
rect 22704 19944 26424 19972
rect 22704 19932 22710 19944
rect 26418 19932 26424 19944
rect 26476 19932 26482 19984
rect 26513 19975 26571 19981
rect 26513 19941 26525 19975
rect 26559 19972 26571 19975
rect 26559 19944 26740 19972
rect 26559 19941 26571 19944
rect 26513 19935 26571 19941
rect 25498 19904 25504 19916
rect 25056 19876 25504 19904
rect 25056 19848 25084 19876
rect 25498 19864 25504 19876
rect 25556 19904 25562 19916
rect 25685 19907 25743 19913
rect 25685 19904 25697 19907
rect 25556 19876 25697 19904
rect 25556 19864 25562 19876
rect 25685 19873 25697 19876
rect 25731 19873 25743 19907
rect 26602 19904 26608 19916
rect 25685 19867 25743 19873
rect 26160 19876 26608 19904
rect 1673 19839 1731 19845
rect 1673 19805 1685 19839
rect 1719 19836 1731 19839
rect 15194 19836 15200 19848
rect 1719 19808 15200 19836
rect 1719 19805 1731 19808
rect 1673 19799 1731 19805
rect 15194 19796 15200 19808
rect 15252 19796 15258 19848
rect 24854 19796 24860 19848
rect 24912 19796 24918 19848
rect 25038 19796 25044 19848
rect 25096 19796 25102 19848
rect 25225 19839 25283 19845
rect 25225 19805 25237 19839
rect 25271 19805 25283 19839
rect 25225 19799 25283 19805
rect 25130 19728 25136 19780
rect 25188 19728 25194 19780
rect 25240 19768 25268 19799
rect 25314 19796 25320 19848
rect 25372 19836 25378 19848
rect 26160 19845 26188 19876
rect 26602 19864 26608 19876
rect 26660 19864 26666 19916
rect 26712 19913 26740 19944
rect 28718 19932 28724 19984
rect 28776 19972 28782 19984
rect 30760 19972 30788 20012
rect 31202 19972 31208 19984
rect 28776 19944 30788 19972
rect 30852 19944 31208 19972
rect 28776 19932 28782 19944
rect 26697 19907 26755 19913
rect 26697 19873 26709 19907
rect 26743 19873 26755 19907
rect 27706 19904 27712 19916
rect 26697 19867 26755 19873
rect 26804 19876 27712 19904
rect 25869 19839 25927 19845
rect 25869 19836 25881 19839
rect 25372 19808 25881 19836
rect 25372 19796 25378 19808
rect 25869 19805 25881 19808
rect 25915 19805 25927 19839
rect 25869 19799 25927 19805
rect 26017 19839 26075 19845
rect 26017 19805 26029 19839
rect 26063 19836 26075 19839
rect 26145 19839 26203 19845
rect 26063 19805 26096 19836
rect 26017 19799 26096 19805
rect 26145 19805 26157 19839
rect 26191 19805 26203 19839
rect 26145 19799 26203 19805
rect 25682 19768 25688 19780
rect 25240 19740 25688 19768
rect 25682 19728 25688 19740
rect 25740 19728 25746 19780
rect 842 19660 848 19712
rect 900 19700 906 19712
rect 1489 19703 1547 19709
rect 1489 19700 1501 19703
rect 900 19672 1501 19700
rect 900 19660 906 19672
rect 1489 19669 1501 19672
rect 1535 19669 1547 19703
rect 26068 19700 26096 19799
rect 26326 19796 26332 19848
rect 26384 19845 26390 19848
rect 26384 19836 26392 19845
rect 26804 19836 26832 19876
rect 27706 19864 27712 19876
rect 27764 19864 27770 19916
rect 29638 19864 29644 19916
rect 29696 19904 29702 19916
rect 30852 19913 30880 19944
rect 31202 19932 31208 19944
rect 31260 19972 31266 19984
rect 31570 19972 31576 19984
rect 31260 19944 31576 19972
rect 31260 19932 31266 19944
rect 31570 19932 31576 19944
rect 31628 19932 31634 19984
rect 31726 19972 31754 20012
rect 33965 20009 33977 20043
rect 34011 20040 34023 20043
rect 34054 20040 34060 20052
rect 34011 20012 34060 20040
rect 34011 20009 34023 20012
rect 33965 20003 34023 20009
rect 34054 20000 34060 20012
rect 34112 20000 34118 20052
rect 34698 20000 34704 20052
rect 34756 20000 34762 20052
rect 34790 20000 34796 20052
rect 34848 20000 34854 20052
rect 35161 20043 35219 20049
rect 35161 20009 35173 20043
rect 35207 20040 35219 20043
rect 36446 20040 36452 20052
rect 35207 20012 36452 20040
rect 35207 20009 35219 20012
rect 35161 20003 35219 20009
rect 36446 20000 36452 20012
rect 36504 20000 36510 20052
rect 36630 20000 36636 20052
rect 36688 20040 36694 20052
rect 36725 20043 36783 20049
rect 36725 20040 36737 20043
rect 36688 20012 36737 20040
rect 36688 20000 36694 20012
rect 36725 20009 36737 20012
rect 36771 20009 36783 20043
rect 36725 20003 36783 20009
rect 41230 20000 41236 20052
rect 41288 20000 41294 20052
rect 41322 20000 41328 20052
rect 41380 20000 41386 20052
rect 47949 20043 48007 20049
rect 47949 20009 47961 20043
rect 47995 20040 48007 20043
rect 48314 20040 48320 20052
rect 47995 20012 48320 20040
rect 47995 20009 48007 20012
rect 47949 20003 48007 20009
rect 48314 20000 48320 20012
rect 48372 20000 48378 20052
rect 48869 20043 48927 20049
rect 48869 20009 48881 20043
rect 48915 20040 48927 20043
rect 49050 20040 49056 20052
rect 48915 20012 49056 20040
rect 48915 20009 48927 20012
rect 48869 20003 48927 20009
rect 49050 20000 49056 20012
rect 49108 20000 49114 20052
rect 49234 20000 49240 20052
rect 49292 20040 49298 20052
rect 49878 20040 49884 20052
rect 49292 20012 49884 20040
rect 49292 20000 49298 20012
rect 49878 20000 49884 20012
rect 49936 20000 49942 20052
rect 50430 20000 50436 20052
rect 50488 20040 50494 20052
rect 50525 20043 50583 20049
rect 50525 20040 50537 20043
rect 50488 20012 50537 20040
rect 50488 20000 50494 20012
rect 50525 20009 50537 20012
rect 50571 20009 50583 20043
rect 51258 20040 51264 20052
rect 50525 20003 50583 20009
rect 51046 20012 51264 20040
rect 33781 19975 33839 19981
rect 33781 19972 33793 19975
rect 31726 19944 33793 19972
rect 33781 19941 33793 19944
rect 33827 19972 33839 19975
rect 34808 19972 34836 20000
rect 35345 19975 35403 19981
rect 35345 19972 35357 19975
rect 33827 19944 34836 19972
rect 34992 19944 35357 19972
rect 33827 19941 33839 19944
rect 33781 19935 33839 19941
rect 30837 19907 30895 19913
rect 30837 19904 30849 19907
rect 29696 19876 30849 19904
rect 29696 19864 29702 19876
rect 30837 19873 30849 19876
rect 30883 19873 30895 19907
rect 31849 19907 31907 19913
rect 31849 19904 31861 19907
rect 30837 19867 30895 19873
rect 31266 19876 31861 19904
rect 26384 19808 26429 19836
rect 26528 19808 26832 19836
rect 26881 19839 26939 19845
rect 26384 19799 26392 19808
rect 26384 19796 26390 19799
rect 26237 19771 26295 19777
rect 26237 19737 26249 19771
rect 26283 19768 26295 19771
rect 26528 19768 26556 19808
rect 26881 19805 26893 19839
rect 26927 19836 26939 19839
rect 28810 19836 28816 19848
rect 26927 19808 28816 19836
rect 26927 19805 26939 19808
rect 26881 19799 26939 19805
rect 28810 19796 28816 19808
rect 28868 19796 28874 19848
rect 30650 19796 30656 19848
rect 30708 19836 30714 19848
rect 31266 19845 31294 19876
rect 31849 19873 31861 19876
rect 31895 19904 31907 19907
rect 32030 19904 32036 19916
rect 31895 19876 32036 19904
rect 31895 19873 31907 19876
rect 31849 19867 31907 19873
rect 32030 19864 32036 19876
rect 32088 19864 32094 19916
rect 31253 19839 31311 19845
rect 31253 19836 31265 19839
rect 30708 19808 31265 19836
rect 30708 19796 30714 19808
rect 31253 19805 31265 19808
rect 31299 19805 31311 19839
rect 31253 19799 31311 19805
rect 31386 19796 31392 19848
rect 31444 19796 31450 19848
rect 31570 19796 31576 19848
rect 31628 19845 31634 19848
rect 31628 19839 31667 19845
rect 31655 19805 31667 19839
rect 31628 19799 31667 19805
rect 31628 19796 31634 19799
rect 31754 19796 31760 19848
rect 31812 19796 31818 19848
rect 33796 19836 33824 19935
rect 34790 19904 34796 19916
rect 34348 19876 34796 19904
rect 34348 19845 34376 19876
rect 34790 19864 34796 19876
rect 34848 19864 34854 19916
rect 34149 19839 34207 19845
rect 34149 19836 34161 19839
rect 33796 19808 34161 19836
rect 34149 19805 34161 19808
rect 34195 19805 34207 19839
rect 34149 19799 34207 19805
rect 34333 19839 34391 19845
rect 34333 19805 34345 19839
rect 34379 19805 34391 19839
rect 34333 19799 34391 19805
rect 26283 19740 26556 19768
rect 26283 19737 26295 19740
rect 26237 19731 26295 19737
rect 26602 19728 26608 19780
rect 26660 19728 26666 19780
rect 27890 19728 27896 19780
rect 27948 19768 27954 19780
rect 28718 19768 28724 19780
rect 27948 19740 28724 19768
rect 27948 19728 27954 19740
rect 28718 19728 28724 19740
rect 28776 19728 28782 19780
rect 29546 19728 29552 19780
rect 29604 19768 29610 19780
rect 30009 19771 30067 19777
rect 30009 19768 30021 19771
rect 29604 19740 30021 19768
rect 29604 19728 29610 19740
rect 29840 19712 29868 19740
rect 30009 19737 30021 19740
rect 30055 19737 30067 19771
rect 30009 19731 30067 19737
rect 30834 19728 30840 19780
rect 30892 19768 30898 19780
rect 31481 19771 31539 19777
rect 30892 19740 31340 19768
rect 30892 19728 30898 19740
rect 26326 19700 26332 19712
rect 26068 19672 26332 19700
rect 1489 19663 1547 19669
rect 26326 19660 26332 19672
rect 26384 19660 26390 19712
rect 26418 19660 26424 19712
rect 26476 19700 26482 19712
rect 27065 19703 27123 19709
rect 27065 19700 27077 19703
rect 26476 19672 27077 19700
rect 26476 19660 26482 19672
rect 27065 19669 27077 19672
rect 27111 19700 27123 19703
rect 27157 19703 27215 19709
rect 27157 19700 27169 19703
rect 27111 19672 27169 19700
rect 27111 19669 27123 19672
rect 27065 19663 27123 19669
rect 27157 19669 27169 19672
rect 27203 19669 27215 19703
rect 27157 19663 27215 19669
rect 28534 19660 28540 19712
rect 28592 19700 28598 19712
rect 28902 19700 28908 19712
rect 28592 19672 28908 19700
rect 28592 19660 28598 19672
rect 28902 19660 28908 19672
rect 28960 19660 28966 19712
rect 29822 19660 29828 19712
rect 29880 19660 29886 19712
rect 30374 19660 30380 19712
rect 30432 19700 30438 19712
rect 31113 19703 31171 19709
rect 31113 19700 31125 19703
rect 30432 19672 31125 19700
rect 30432 19660 30438 19672
rect 31113 19669 31125 19672
rect 31159 19669 31171 19703
rect 31312 19700 31340 19740
rect 31481 19737 31493 19771
rect 31527 19768 31539 19771
rect 31527 19740 32168 19768
rect 31527 19737 31539 19740
rect 31481 19731 31539 19737
rect 31496 19700 31524 19731
rect 32140 19709 32168 19740
rect 34238 19728 34244 19780
rect 34296 19728 34302 19780
rect 31312 19672 31524 19700
rect 32125 19703 32183 19709
rect 31113 19663 31171 19669
rect 32125 19669 32137 19703
rect 32171 19700 32183 19703
rect 32214 19700 32220 19712
rect 32171 19672 32220 19700
rect 32171 19669 32183 19672
rect 32125 19663 32183 19669
rect 32214 19660 32220 19672
rect 32272 19700 32278 19712
rect 34348 19700 34376 19799
rect 34514 19796 34520 19848
rect 34572 19796 34578 19848
rect 34606 19796 34612 19848
rect 34664 19796 34670 19848
rect 34698 19796 34704 19848
rect 34756 19836 34762 19848
rect 34992 19845 35020 19944
rect 35345 19941 35357 19944
rect 35391 19941 35403 19975
rect 35345 19935 35403 19941
rect 35434 19932 35440 19984
rect 35492 19972 35498 19984
rect 36648 19972 36676 20000
rect 35492 19944 36676 19972
rect 41248 19972 41276 20000
rect 51046 19984 51074 20012
rect 51258 20000 51264 20012
rect 51316 20040 51322 20052
rect 51316 20012 53236 20040
rect 51316 20000 51322 20012
rect 41785 19975 41843 19981
rect 41785 19972 41797 19975
rect 41248 19944 41797 19972
rect 35492 19932 35498 19944
rect 41785 19941 41797 19944
rect 41831 19972 41843 19975
rect 42058 19972 42064 19984
rect 41831 19944 42064 19972
rect 41831 19941 41843 19944
rect 41785 19935 41843 19941
rect 42058 19932 42064 19944
rect 42116 19932 42122 19984
rect 48222 19932 48228 19984
rect 48280 19972 48286 19984
rect 50982 19972 50988 19984
rect 48280 19944 50988 19972
rect 48280 19932 48286 19944
rect 50982 19932 50988 19944
rect 51040 19944 51074 19984
rect 51040 19932 51046 19944
rect 37093 19907 37151 19913
rect 35360 19876 36584 19904
rect 35360 19848 35388 19876
rect 34885 19839 34943 19845
rect 34885 19836 34897 19839
rect 34756 19808 34897 19836
rect 34756 19796 34762 19808
rect 34885 19805 34897 19808
rect 34931 19805 34943 19839
rect 34885 19799 34943 19805
rect 34977 19839 35035 19845
rect 34977 19805 34989 19839
rect 35023 19805 35035 19839
rect 34977 19799 35035 19805
rect 35253 19839 35311 19845
rect 35253 19805 35265 19839
rect 35299 19836 35311 19839
rect 35342 19836 35348 19848
rect 35299 19808 35348 19836
rect 35299 19805 35311 19808
rect 35253 19799 35311 19805
rect 35342 19796 35348 19808
rect 35400 19796 35406 19848
rect 35529 19839 35587 19845
rect 35529 19805 35541 19839
rect 35575 19805 35587 19839
rect 35529 19799 35587 19805
rect 34624 19768 34652 19796
rect 35544 19768 35572 19799
rect 35710 19796 35716 19848
rect 35768 19796 35774 19848
rect 35897 19839 35955 19845
rect 35897 19805 35909 19839
rect 35943 19836 35955 19839
rect 36078 19836 36084 19848
rect 35943 19808 36084 19836
rect 35943 19805 35955 19808
rect 35897 19799 35955 19805
rect 36078 19796 36084 19808
rect 36136 19796 36142 19848
rect 36556 19845 36584 19876
rect 37093 19873 37105 19907
rect 37139 19904 37151 19907
rect 37918 19904 37924 19916
rect 37139 19876 37924 19904
rect 37139 19873 37151 19876
rect 37093 19867 37151 19873
rect 37918 19864 37924 19876
rect 37976 19864 37982 19916
rect 44174 19864 44180 19916
rect 44232 19904 44238 19916
rect 44821 19907 44879 19913
rect 44821 19904 44833 19907
rect 44232 19876 44833 19904
rect 44232 19864 44238 19876
rect 44821 19873 44833 19876
rect 44867 19873 44879 19907
rect 44821 19867 44879 19873
rect 46382 19864 46388 19916
rect 46440 19904 46446 19916
rect 46842 19904 46848 19916
rect 46440 19876 46848 19904
rect 46440 19864 46446 19876
rect 46842 19864 46848 19876
rect 46900 19904 46906 19916
rect 48685 19907 48743 19913
rect 48685 19904 48697 19907
rect 46900 19876 48697 19904
rect 46900 19864 46906 19876
rect 48685 19873 48697 19876
rect 48731 19873 48743 19907
rect 51445 19907 51503 19913
rect 48685 19867 48743 19873
rect 48884 19876 51120 19904
rect 36173 19839 36231 19845
rect 36173 19805 36185 19839
rect 36219 19805 36231 19839
rect 36173 19799 36231 19805
rect 36541 19839 36599 19845
rect 36541 19805 36553 19839
rect 36587 19805 36599 19839
rect 36541 19799 36599 19805
rect 34624 19740 35572 19768
rect 35618 19728 35624 19780
rect 35676 19768 35682 19780
rect 35676 19740 36124 19768
rect 35676 19728 35682 19740
rect 36096 19712 36124 19740
rect 32272 19672 34376 19700
rect 32272 19660 32278 19672
rect 34606 19660 34612 19712
rect 34664 19700 34670 19712
rect 35989 19703 36047 19709
rect 35989 19700 36001 19703
rect 34664 19672 36001 19700
rect 34664 19660 34670 19672
rect 35989 19669 36001 19672
rect 36035 19669 36047 19703
rect 35989 19663 36047 19669
rect 36078 19660 36084 19712
rect 36136 19660 36142 19712
rect 36188 19700 36216 19799
rect 36906 19796 36912 19848
rect 36964 19796 36970 19848
rect 38470 19796 38476 19848
rect 38528 19796 38534 19848
rect 39482 19836 39488 19848
rect 38856 19808 39488 19836
rect 36262 19728 36268 19780
rect 36320 19728 36326 19780
rect 36357 19771 36415 19777
rect 36357 19737 36369 19771
rect 36403 19768 36415 19771
rect 36446 19768 36452 19780
rect 36403 19740 36452 19768
rect 36403 19737 36415 19740
rect 36357 19731 36415 19737
rect 36446 19728 36452 19740
rect 36504 19728 36510 19780
rect 37366 19728 37372 19780
rect 37424 19728 37430 19780
rect 38856 19712 38884 19808
rect 39482 19796 39488 19808
rect 39540 19796 39546 19848
rect 41506 19836 41512 19848
rect 41386 19808 41512 19836
rect 39114 19728 39120 19780
rect 39172 19768 39178 19780
rect 41046 19768 41052 19780
rect 39172 19740 41052 19768
rect 39172 19728 39178 19740
rect 41046 19728 41052 19740
rect 41104 19768 41110 19780
rect 41386 19768 41414 19808
rect 41506 19796 41512 19808
rect 41564 19796 41570 19848
rect 41601 19839 41659 19845
rect 41601 19805 41613 19839
rect 41647 19805 41659 19839
rect 41601 19799 41659 19805
rect 41104 19740 41414 19768
rect 41616 19768 41644 19799
rect 41690 19796 41696 19848
rect 41748 19836 41754 19848
rect 41874 19836 41880 19848
rect 41748 19808 41880 19836
rect 41748 19796 41754 19808
rect 41874 19796 41880 19808
rect 41932 19796 41938 19848
rect 45186 19796 45192 19848
rect 45244 19796 45250 19848
rect 45370 19796 45376 19848
rect 45428 19796 45434 19848
rect 45462 19796 45468 19848
rect 45520 19796 45526 19848
rect 46658 19796 46664 19848
rect 46716 19836 46722 19848
rect 47397 19839 47455 19845
rect 47397 19836 47409 19839
rect 46716 19808 47409 19836
rect 46716 19796 46722 19808
rect 47397 19805 47409 19808
rect 47443 19805 47455 19839
rect 47397 19799 47455 19805
rect 47762 19796 47768 19848
rect 47820 19796 47826 19848
rect 48041 19839 48099 19845
rect 48041 19805 48053 19839
rect 48087 19805 48099 19839
rect 48041 19799 48099 19805
rect 42426 19768 42432 19780
rect 41616 19740 42432 19768
rect 41104 19728 41110 19740
rect 42426 19728 42432 19740
rect 42484 19728 42490 19780
rect 42702 19728 42708 19780
rect 42760 19768 42766 19780
rect 44545 19771 44603 19777
rect 42760 19740 43378 19768
rect 42760 19728 42766 19740
rect 44545 19737 44557 19771
rect 44591 19768 44603 19771
rect 45005 19771 45063 19777
rect 45005 19768 45017 19771
rect 44591 19740 45017 19768
rect 44591 19737 44603 19740
rect 44545 19731 44603 19737
rect 45005 19737 45017 19740
rect 45051 19737 45063 19771
rect 45005 19731 45063 19737
rect 45554 19728 45560 19780
rect 45612 19728 45618 19780
rect 47486 19728 47492 19780
rect 47544 19768 47550 19780
rect 47581 19771 47639 19777
rect 47581 19768 47593 19771
rect 47544 19740 47593 19768
rect 47544 19728 47550 19740
rect 47581 19737 47593 19740
rect 47627 19737 47639 19771
rect 47581 19731 47639 19737
rect 47673 19771 47731 19777
rect 47673 19737 47685 19771
rect 47719 19768 47731 19771
rect 48056 19768 48084 19799
rect 48130 19796 48136 19848
rect 48188 19836 48194 19848
rect 48317 19839 48375 19845
rect 48317 19836 48329 19839
rect 48188 19808 48329 19836
rect 48188 19796 48194 19808
rect 48317 19805 48329 19808
rect 48363 19805 48375 19839
rect 48317 19799 48375 19805
rect 48406 19796 48412 19848
rect 48464 19796 48470 19848
rect 47719 19740 48084 19768
rect 47719 19737 47731 19740
rect 47673 19731 47731 19737
rect 36722 19700 36728 19712
rect 36188 19672 36728 19700
rect 36722 19660 36728 19672
rect 36780 19660 36786 19712
rect 38838 19660 38844 19712
rect 38896 19660 38902 19712
rect 38930 19660 38936 19712
rect 38988 19660 38994 19712
rect 43073 19703 43131 19709
rect 43073 19669 43085 19703
rect 43119 19700 43131 19703
rect 44358 19700 44364 19712
rect 43119 19672 44364 19700
rect 43119 19669 43131 19672
rect 43073 19663 43131 19669
rect 44358 19660 44364 19672
rect 44416 19700 44422 19712
rect 46658 19700 46664 19712
rect 44416 19672 46664 19700
rect 44416 19660 44422 19672
rect 46658 19660 46664 19672
rect 46716 19660 46722 19712
rect 46842 19660 46848 19712
rect 46900 19660 46906 19712
rect 47596 19700 47624 19731
rect 47946 19700 47952 19712
rect 47596 19672 47952 19700
rect 47946 19660 47952 19672
rect 48004 19660 48010 19712
rect 48056 19700 48084 19740
rect 48222 19728 48228 19780
rect 48280 19728 48286 19780
rect 48884 19768 48912 19876
rect 49050 19796 49056 19848
rect 49108 19796 49114 19848
rect 49145 19839 49203 19845
rect 49145 19805 49157 19839
rect 49191 19836 49203 19839
rect 49191 19808 49372 19836
rect 49191 19805 49203 19808
rect 49145 19799 49203 19805
rect 48424 19740 48912 19768
rect 49237 19771 49295 19777
rect 48424 19700 48452 19740
rect 49237 19737 49249 19771
rect 49283 19737 49295 19771
rect 49344 19768 49372 19808
rect 49418 19796 49424 19848
rect 49476 19796 49482 19848
rect 50430 19796 50436 19848
rect 50488 19836 50494 19848
rect 50706 19836 50712 19848
rect 50488 19808 50712 19836
rect 50488 19796 50494 19808
rect 50706 19796 50712 19808
rect 50764 19796 50770 19848
rect 50802 19839 50860 19845
rect 50802 19805 50814 19839
rect 50848 19836 50860 19839
rect 50890 19836 50896 19848
rect 50848 19808 50896 19836
rect 50848 19805 50860 19808
rect 50802 19799 50860 19805
rect 50816 19768 50844 19799
rect 50890 19796 50896 19808
rect 50948 19796 50954 19848
rect 50982 19796 50988 19848
rect 51040 19796 51046 19848
rect 51092 19780 51120 19876
rect 51445 19873 51457 19907
rect 51491 19904 51503 19907
rect 51718 19904 51724 19916
rect 51491 19876 51724 19904
rect 51491 19873 51503 19876
rect 51445 19867 51503 19873
rect 51718 19864 51724 19876
rect 51776 19864 51782 19916
rect 52914 19864 52920 19916
rect 52972 19864 52978 19916
rect 51174 19839 51232 19845
rect 51174 19805 51186 19839
rect 51220 19805 51232 19839
rect 52932 19836 52960 19864
rect 52854 19808 52960 19836
rect 51174 19799 51232 19805
rect 49344 19740 50844 19768
rect 49237 19731 49295 19737
rect 48056 19672 48452 19700
rect 48593 19703 48651 19709
rect 48593 19669 48605 19703
rect 48639 19700 48651 19703
rect 48774 19700 48780 19712
rect 48639 19672 48780 19700
rect 48639 19669 48651 19672
rect 48593 19663 48651 19669
rect 48774 19660 48780 19672
rect 48832 19660 48838 19712
rect 49252 19700 49280 19731
rect 51074 19728 51080 19780
rect 51132 19728 51138 19780
rect 49510 19700 49516 19712
rect 49252 19672 49516 19700
rect 49510 19660 49516 19672
rect 49568 19660 49574 19712
rect 49786 19660 49792 19712
rect 49844 19660 49850 19712
rect 50430 19660 50436 19712
rect 50488 19700 50494 19712
rect 51184 19700 51212 19799
rect 51718 19728 51724 19780
rect 51776 19728 51782 19780
rect 53208 19768 53236 20012
rect 53834 20000 53840 20052
rect 53892 20040 53898 20052
rect 53929 20043 53987 20049
rect 53929 20040 53941 20043
rect 53892 20012 53941 20040
rect 53892 20000 53898 20012
rect 53929 20009 53941 20012
rect 53975 20009 53987 20043
rect 53929 20003 53987 20009
rect 55125 20043 55183 20049
rect 55125 20009 55137 20043
rect 55171 20040 55183 20043
rect 55398 20040 55404 20052
rect 55171 20012 55404 20040
rect 55171 20009 55183 20012
rect 55125 20003 55183 20009
rect 55398 20000 55404 20012
rect 55456 20000 55462 20052
rect 55950 20000 55956 20052
rect 56008 20040 56014 20052
rect 57057 20043 57115 20049
rect 57057 20040 57069 20043
rect 56008 20012 57069 20040
rect 56008 20000 56014 20012
rect 57057 20009 57069 20012
rect 57103 20009 57115 20043
rect 57057 20003 57115 20009
rect 53466 19864 53472 19916
rect 53524 19904 53530 19916
rect 55309 19907 55367 19913
rect 53524 19876 53696 19904
rect 53524 19864 53530 19876
rect 53282 19796 53288 19848
rect 53340 19796 53346 19848
rect 53374 19796 53380 19848
rect 53432 19836 53438 19848
rect 53668 19845 53696 19876
rect 55309 19873 55321 19907
rect 55355 19904 55367 19907
rect 56134 19904 56140 19916
rect 55355 19876 56140 19904
rect 55355 19873 55367 19876
rect 55309 19867 55367 19873
rect 56134 19864 56140 19876
rect 56192 19864 56198 19916
rect 53653 19839 53711 19845
rect 53432 19808 53477 19836
rect 53432 19796 53438 19808
rect 53653 19805 53665 19839
rect 53699 19805 53711 19839
rect 53653 19799 53711 19805
rect 53742 19796 53748 19848
rect 53800 19845 53806 19848
rect 53800 19836 53808 19845
rect 53800 19808 53845 19836
rect 53800 19799 53808 19808
rect 53800 19796 53806 19799
rect 54478 19796 54484 19848
rect 54536 19796 54542 19848
rect 54570 19796 54576 19848
rect 54628 19836 54634 19848
rect 54628 19808 54673 19836
rect 54628 19796 54634 19808
rect 54938 19796 54944 19848
rect 54996 19845 55002 19848
rect 54996 19799 55004 19845
rect 54996 19796 55002 19799
rect 56686 19796 56692 19848
rect 56744 19796 56750 19848
rect 57885 19839 57943 19845
rect 57885 19805 57897 19839
rect 57931 19836 57943 19839
rect 58158 19836 58164 19848
rect 57931 19808 58164 19836
rect 57931 19805 57943 19808
rect 57885 19799 57943 19805
rect 58158 19796 58164 19808
rect 58216 19796 58222 19848
rect 58250 19796 58256 19848
rect 58308 19796 58314 19848
rect 53561 19771 53619 19777
rect 53561 19768 53573 19771
rect 53208 19740 53573 19768
rect 53561 19737 53573 19740
rect 53607 19737 53619 19771
rect 53561 19731 53619 19737
rect 54757 19771 54815 19777
rect 54757 19737 54769 19771
rect 54803 19737 54815 19771
rect 54757 19731 54815 19737
rect 50488 19672 51212 19700
rect 51353 19703 51411 19709
rect 50488 19660 50494 19672
rect 51353 19669 51365 19703
rect 51399 19700 51411 19703
rect 51810 19700 51816 19712
rect 51399 19672 51816 19700
rect 51399 19669 51411 19672
rect 51353 19663 51411 19669
rect 51810 19660 51816 19672
rect 51868 19660 51874 19712
rect 52086 19660 52092 19712
rect 52144 19700 52150 19712
rect 53193 19703 53251 19709
rect 53193 19700 53205 19703
rect 52144 19672 53205 19700
rect 52144 19660 52150 19672
rect 53193 19669 53205 19672
rect 53239 19700 53251 19703
rect 53466 19700 53472 19712
rect 53239 19672 53472 19700
rect 53239 19669 53251 19672
rect 53193 19663 53251 19669
rect 53466 19660 53472 19672
rect 53524 19660 53530 19712
rect 53576 19700 53604 19731
rect 54772 19700 54800 19731
rect 54846 19728 54852 19780
rect 54904 19728 54910 19780
rect 55582 19728 55588 19780
rect 55640 19728 55646 19780
rect 55950 19700 55956 19712
rect 53576 19672 55956 19700
rect 55950 19660 55956 19672
rect 56008 19660 56014 19712
rect 57882 19660 57888 19712
rect 57940 19700 57946 19712
rect 58069 19703 58127 19709
rect 58069 19700 58081 19703
rect 57940 19672 58081 19700
rect 57940 19660 57946 19672
rect 58069 19669 58081 19672
rect 58115 19669 58127 19703
rect 58069 19663 58127 19669
rect 58434 19660 58440 19712
rect 58492 19660 58498 19712
rect 1104 19610 58880 19632
rect 1104 19558 4874 19610
rect 4926 19558 4938 19610
rect 4990 19558 5002 19610
rect 5054 19558 5066 19610
rect 5118 19558 5130 19610
rect 5182 19558 35594 19610
rect 35646 19558 35658 19610
rect 35710 19558 35722 19610
rect 35774 19558 35786 19610
rect 35838 19558 35850 19610
rect 35902 19558 58880 19610
rect 1104 19536 58880 19558
rect 15013 19499 15071 19505
rect 15013 19465 15025 19499
rect 15059 19496 15071 19499
rect 15194 19496 15200 19508
rect 15059 19468 15200 19496
rect 15059 19465 15071 19468
rect 15013 19459 15071 19465
rect 15194 19456 15200 19468
rect 15252 19456 15258 19508
rect 19334 19496 19340 19508
rect 18984 19468 19340 19496
rect 16114 19320 16120 19372
rect 16172 19369 16178 19372
rect 16172 19323 16184 19369
rect 16393 19363 16451 19369
rect 16393 19329 16405 19363
rect 16439 19360 16451 19363
rect 16666 19360 16672 19372
rect 16439 19332 16672 19360
rect 16439 19329 16451 19332
rect 16393 19323 16451 19329
rect 16172 19320 16178 19323
rect 16666 19320 16672 19332
rect 16724 19320 16730 19372
rect 18984 19369 19012 19468
rect 19334 19456 19340 19468
rect 19392 19456 19398 19508
rect 19429 19499 19487 19505
rect 19429 19465 19441 19499
rect 19475 19465 19487 19499
rect 19429 19459 19487 19465
rect 19444 19428 19472 19459
rect 20070 19456 20076 19508
rect 20128 19496 20134 19508
rect 22465 19499 22523 19505
rect 22465 19496 22477 19499
rect 20128 19468 22477 19496
rect 20128 19456 20134 19468
rect 19076 19400 19472 19428
rect 19705 19431 19763 19437
rect 19076 19369 19104 19400
rect 19705 19397 19717 19431
rect 19751 19428 19763 19431
rect 19886 19428 19892 19440
rect 19751 19400 19892 19428
rect 19751 19397 19763 19400
rect 19705 19391 19763 19397
rect 19886 19388 19892 19400
rect 19944 19388 19950 19440
rect 20438 19428 20444 19440
rect 19996 19400 20444 19428
rect 18969 19363 19027 19369
rect 18969 19329 18981 19363
rect 19015 19329 19027 19363
rect 18969 19323 19027 19329
rect 19061 19363 19119 19369
rect 19061 19329 19073 19363
rect 19107 19329 19119 19363
rect 19061 19323 19119 19329
rect 19337 19363 19395 19369
rect 19337 19329 19349 19363
rect 19383 19360 19395 19363
rect 19518 19360 19524 19372
rect 19383 19332 19524 19360
rect 19383 19329 19395 19332
rect 19337 19323 19395 19329
rect 19518 19320 19524 19332
rect 19576 19320 19582 19372
rect 19610 19320 19616 19372
rect 19668 19320 19674 19372
rect 19794 19320 19800 19372
rect 19852 19320 19858 19372
rect 19996 19369 20024 19400
rect 20438 19388 20444 19400
rect 20496 19388 20502 19440
rect 19981 19363 20039 19369
rect 19981 19329 19993 19363
rect 20027 19329 20039 19363
rect 21928 19360 21956 19468
rect 22465 19465 22477 19468
rect 22511 19465 22523 19499
rect 22465 19459 22523 19465
rect 22186 19369 22192 19372
rect 21988 19363 22046 19369
rect 21988 19360 22000 19363
rect 21928 19332 22000 19360
rect 19981 19323 20039 19329
rect 21988 19329 22000 19332
rect 22034 19329 22046 19363
rect 21988 19323 22046 19329
rect 22157 19363 22192 19369
rect 22157 19329 22169 19363
rect 22157 19323 22192 19329
rect 22186 19320 22192 19323
rect 22244 19320 22250 19372
rect 22370 19320 22376 19372
rect 22428 19320 22434 19372
rect 22480 19360 22508 19459
rect 25682 19456 25688 19508
rect 25740 19496 25746 19508
rect 26142 19496 26148 19508
rect 25740 19468 26148 19496
rect 25740 19456 25746 19468
rect 26142 19456 26148 19468
rect 26200 19456 26206 19508
rect 26234 19456 26240 19508
rect 26292 19496 26298 19508
rect 26605 19499 26663 19505
rect 26605 19496 26617 19499
rect 26292 19468 26617 19496
rect 26292 19456 26298 19468
rect 26605 19465 26617 19468
rect 26651 19496 26663 19499
rect 26878 19496 26884 19508
rect 26651 19468 26884 19496
rect 26651 19465 26663 19468
rect 26605 19459 26663 19465
rect 26878 19456 26884 19468
rect 26936 19496 26942 19508
rect 28166 19496 28172 19508
rect 26936 19468 28172 19496
rect 26936 19456 26942 19468
rect 28166 19456 28172 19468
rect 28224 19456 28230 19508
rect 28534 19496 28540 19508
rect 28276 19468 28540 19496
rect 24762 19388 24768 19440
rect 24820 19428 24826 19440
rect 28276 19437 28304 19468
rect 28534 19456 28540 19468
rect 28592 19456 28598 19508
rect 28629 19499 28687 19505
rect 28629 19465 28641 19499
rect 28675 19496 28687 19499
rect 28810 19496 28816 19508
rect 28675 19468 28816 19496
rect 28675 19465 28687 19468
rect 28629 19459 28687 19465
rect 28810 19456 28816 19468
rect 28868 19456 28874 19508
rect 28902 19456 28908 19508
rect 28960 19456 28966 19508
rect 31128 19468 31754 19496
rect 28261 19431 28319 19437
rect 24820 19400 28028 19428
rect 24820 19388 24826 19400
rect 23014 19360 23020 19372
rect 22480 19332 23020 19360
rect 23014 19320 23020 19332
rect 23072 19320 23078 19372
rect 23106 19320 23112 19372
rect 23164 19320 23170 19372
rect 23290 19320 23296 19372
rect 23348 19360 23354 19372
rect 23385 19363 23443 19369
rect 23385 19360 23397 19363
rect 23348 19332 23397 19360
rect 23348 19320 23354 19332
rect 23385 19329 23397 19332
rect 23431 19329 23443 19363
rect 26329 19363 26387 19369
rect 23385 19323 23443 19329
rect 25240 19332 26188 19360
rect 18138 19252 18144 19304
rect 18196 19292 18202 19304
rect 24578 19292 24584 19304
rect 18196 19264 24584 19292
rect 18196 19252 18202 19264
rect 24578 19252 24584 19264
rect 24636 19252 24642 19304
rect 25240 19292 25268 19332
rect 24688 19264 25268 19292
rect 19334 19184 19340 19236
rect 19392 19224 19398 19236
rect 20070 19224 20076 19236
rect 19392 19196 20076 19224
rect 19392 19184 19398 19196
rect 20070 19184 20076 19196
rect 20128 19184 20134 19236
rect 23293 19227 23351 19233
rect 23293 19224 23305 19227
rect 22296 19196 23305 19224
rect 17586 19116 17592 19168
rect 17644 19156 17650 19168
rect 18785 19159 18843 19165
rect 18785 19156 18797 19159
rect 17644 19128 18797 19156
rect 17644 19116 17650 19128
rect 18785 19125 18797 19128
rect 18831 19125 18843 19159
rect 18785 19119 18843 19125
rect 19242 19116 19248 19168
rect 19300 19116 19306 19168
rect 21821 19159 21879 19165
rect 21821 19125 21833 19159
rect 21867 19156 21879 19159
rect 21910 19156 21916 19168
rect 21867 19128 21916 19156
rect 21867 19125 21879 19128
rect 21821 19119 21879 19125
rect 21910 19116 21916 19128
rect 21968 19116 21974 19168
rect 22094 19116 22100 19168
rect 22152 19156 22158 19168
rect 22296 19165 22324 19196
rect 23293 19193 23305 19196
rect 23339 19193 23351 19227
rect 23293 19187 23351 19193
rect 23569 19227 23627 19233
rect 23569 19193 23581 19227
rect 23615 19224 23627 19227
rect 24688 19224 24716 19264
rect 23615 19196 24716 19224
rect 23615 19193 23627 19196
rect 23569 19187 23627 19193
rect 22281 19159 22339 19165
rect 22281 19156 22293 19159
rect 22152 19128 22293 19156
rect 22152 19116 22158 19128
rect 22281 19125 22293 19128
rect 22327 19125 22339 19159
rect 22281 19119 22339 19125
rect 22554 19116 22560 19168
rect 22612 19156 22618 19168
rect 22833 19159 22891 19165
rect 22833 19156 22845 19159
rect 22612 19128 22845 19156
rect 22612 19116 22618 19128
rect 22833 19125 22845 19128
rect 22879 19125 22891 19159
rect 22833 19119 22891 19125
rect 23014 19116 23020 19168
rect 23072 19156 23078 19168
rect 23584 19156 23612 19187
rect 25866 19184 25872 19236
rect 25924 19224 25930 19236
rect 26160 19224 26188 19332
rect 26329 19329 26341 19363
rect 26375 19360 26387 19363
rect 26510 19360 26516 19372
rect 26375 19332 26516 19360
rect 26375 19329 26387 19332
rect 26329 19323 26387 19329
rect 26510 19320 26516 19332
rect 26568 19320 26574 19372
rect 28000 19369 28028 19400
rect 28261 19397 28273 19431
rect 28307 19397 28319 19431
rect 28261 19391 28319 19397
rect 28353 19431 28411 19437
rect 28353 19397 28365 19431
rect 28399 19428 28411 19431
rect 30282 19428 30288 19440
rect 28399 19400 30288 19428
rect 28399 19397 28411 19400
rect 28353 19391 28411 19397
rect 30282 19388 30288 19400
rect 30340 19388 30346 19440
rect 27985 19363 28043 19369
rect 27985 19329 27997 19363
rect 28031 19329 28043 19363
rect 27985 19323 28043 19329
rect 28133 19363 28191 19369
rect 28133 19329 28145 19363
rect 28179 19360 28191 19363
rect 28491 19363 28549 19369
rect 28179 19329 28212 19360
rect 28133 19323 28212 19329
rect 28491 19329 28503 19363
rect 28537 19360 28549 19363
rect 28718 19360 28724 19372
rect 28537 19332 28724 19360
rect 28537 19329 28549 19332
rect 28491 19323 28549 19329
rect 26602 19252 26608 19304
rect 26660 19292 26666 19304
rect 27246 19292 27252 19304
rect 26660 19264 27252 19292
rect 26660 19252 26666 19264
rect 27246 19252 27252 19264
rect 27304 19252 27310 19304
rect 28184 19292 28212 19323
rect 28718 19320 28724 19332
rect 28776 19320 28782 19372
rect 29730 19320 29736 19372
rect 29788 19360 29794 19372
rect 30190 19360 30196 19372
rect 29788 19332 30196 19360
rect 29788 19320 29794 19332
rect 30190 19320 30196 19332
rect 30248 19360 30254 19372
rect 31128 19369 31156 19468
rect 31726 19428 31754 19468
rect 34238 19456 34244 19508
rect 34296 19496 34302 19508
rect 36262 19496 36268 19508
rect 34296 19468 36268 19496
rect 34296 19456 34302 19468
rect 36262 19456 36268 19468
rect 36320 19456 36326 19508
rect 38933 19499 38991 19505
rect 38933 19496 38945 19499
rect 38212 19468 38945 19496
rect 31726 19400 34284 19428
rect 31113 19363 31171 19369
rect 31113 19360 31125 19363
rect 30248 19332 31125 19360
rect 30248 19320 30254 19332
rect 31113 19329 31125 19332
rect 31159 19329 31171 19363
rect 31113 19323 31171 19329
rect 31205 19363 31263 19369
rect 31205 19329 31217 19363
rect 31251 19329 31263 19363
rect 31205 19323 31263 19329
rect 28626 19292 28632 19304
rect 28184 19264 28632 19292
rect 28626 19252 28632 19264
rect 28684 19252 28690 19304
rect 30558 19252 30564 19304
rect 30616 19292 30622 19304
rect 31220 19292 31248 19323
rect 31478 19320 31484 19372
rect 31536 19320 31542 19372
rect 31662 19320 31668 19372
rect 31720 19360 31726 19372
rect 33594 19360 33600 19372
rect 31720 19332 33600 19360
rect 31720 19320 31726 19332
rect 33594 19320 33600 19332
rect 33652 19360 33658 19372
rect 34149 19363 34207 19369
rect 34149 19360 34161 19363
rect 33652 19332 34161 19360
rect 33652 19320 33658 19332
rect 34149 19329 34161 19332
rect 34195 19329 34207 19363
rect 34256 19360 34284 19400
rect 35342 19388 35348 19440
rect 35400 19388 35406 19440
rect 34422 19360 34428 19372
rect 34256 19332 34428 19360
rect 34149 19323 34207 19329
rect 34422 19320 34428 19332
rect 34480 19320 34486 19372
rect 35943 19363 36001 19369
rect 35943 19329 35955 19363
rect 35989 19360 36001 19363
rect 36078 19360 36084 19372
rect 35989 19332 36084 19360
rect 35989 19329 36001 19332
rect 35943 19323 36001 19329
rect 36078 19320 36084 19332
rect 36136 19360 36142 19372
rect 36354 19360 36360 19372
rect 36136 19332 36360 19360
rect 36136 19320 36142 19332
rect 36354 19320 36360 19332
rect 36412 19320 36418 19372
rect 38102 19320 38108 19372
rect 38160 19320 38166 19372
rect 38212 19369 38240 19468
rect 38933 19465 38945 19468
rect 38979 19465 38991 19499
rect 40494 19496 40500 19508
rect 38933 19459 38991 19465
rect 40420 19468 40500 19496
rect 40420 19428 40448 19468
rect 40494 19456 40500 19468
rect 40552 19496 40558 19508
rect 44913 19499 44971 19505
rect 40552 19468 40908 19496
rect 40552 19456 40558 19468
rect 38396 19400 40448 19428
rect 38197 19363 38255 19369
rect 38197 19329 38209 19363
rect 38243 19329 38255 19363
rect 38197 19323 38255 19329
rect 30616 19264 31248 19292
rect 30616 19252 30622 19264
rect 34514 19252 34520 19304
rect 34572 19252 34578 19304
rect 34698 19252 34704 19304
rect 34756 19292 34762 19304
rect 35434 19292 35440 19304
rect 34756 19264 35440 19292
rect 34756 19252 34762 19264
rect 35434 19252 35440 19264
rect 35492 19252 35498 19304
rect 37366 19252 37372 19304
rect 37424 19292 37430 19304
rect 37921 19295 37979 19301
rect 37921 19292 37933 19295
rect 37424 19264 37933 19292
rect 37424 19252 37430 19264
rect 37921 19261 37933 19264
rect 37967 19261 37979 19295
rect 37921 19255 37979 19261
rect 38010 19252 38016 19304
rect 38068 19292 38074 19304
rect 38396 19292 38424 19400
rect 38473 19363 38531 19369
rect 38473 19329 38485 19363
rect 38519 19360 38531 19363
rect 38930 19360 38936 19372
rect 38519 19332 38936 19360
rect 38519 19329 38531 19332
rect 38473 19323 38531 19329
rect 38930 19320 38936 19332
rect 38988 19320 38994 19372
rect 39114 19320 39120 19372
rect 39172 19320 39178 19372
rect 39206 19320 39212 19372
rect 39264 19320 39270 19372
rect 39301 19363 39359 19369
rect 39301 19329 39313 19363
rect 39347 19360 39359 19363
rect 39485 19363 39543 19369
rect 39347 19332 39436 19360
rect 39347 19329 39359 19332
rect 39301 19323 39359 19329
rect 38068 19264 38424 19292
rect 39408 19292 39436 19332
rect 39485 19329 39497 19363
rect 39531 19360 39543 19363
rect 40034 19360 40040 19372
rect 39531 19332 40040 19360
rect 39531 19329 39543 19332
rect 39485 19323 39543 19329
rect 40034 19320 40040 19332
rect 40092 19360 40098 19372
rect 40218 19360 40224 19372
rect 40092 19332 40224 19360
rect 40092 19320 40098 19332
rect 40218 19320 40224 19332
rect 40276 19320 40282 19372
rect 40420 19369 40448 19400
rect 40678 19388 40684 19440
rect 40736 19428 40742 19440
rect 40773 19431 40831 19437
rect 40773 19428 40785 19431
rect 40736 19400 40785 19428
rect 40736 19388 40742 19400
rect 40773 19397 40785 19400
rect 40819 19397 40831 19431
rect 40773 19391 40831 19397
rect 40405 19363 40463 19369
rect 40405 19329 40417 19363
rect 40451 19329 40463 19363
rect 40405 19323 40463 19329
rect 39408 19264 40724 19292
rect 38068 19252 38074 19264
rect 28258 19224 28264 19236
rect 25924 19196 26096 19224
rect 26160 19196 28264 19224
rect 25924 19184 25930 19196
rect 23072 19128 23612 19156
rect 23072 19116 23078 19128
rect 25038 19116 25044 19168
rect 25096 19156 25102 19168
rect 25958 19156 25964 19168
rect 25096 19128 25964 19156
rect 25096 19116 25102 19128
rect 25958 19116 25964 19128
rect 26016 19116 26022 19168
rect 26068 19156 26096 19196
rect 28258 19184 28264 19196
rect 28316 19184 28322 19236
rect 35526 19184 35532 19236
rect 35584 19224 35590 19236
rect 40402 19224 40408 19236
rect 35584 19196 40408 19224
rect 35584 19184 35590 19196
rect 40402 19184 40408 19196
rect 40460 19184 40466 19236
rect 26970 19156 26976 19168
rect 26068 19128 26976 19156
rect 26970 19116 26976 19128
rect 27028 19116 27034 19168
rect 30929 19159 30987 19165
rect 30929 19125 30941 19159
rect 30975 19156 30987 19159
rect 31018 19156 31024 19168
rect 30975 19128 31024 19156
rect 30975 19125 30987 19128
rect 30929 19119 30987 19125
rect 31018 19116 31024 19128
rect 31076 19116 31082 19168
rect 31389 19159 31447 19165
rect 31389 19125 31401 19159
rect 31435 19156 31447 19159
rect 32490 19156 32496 19168
rect 31435 19128 32496 19156
rect 31435 19125 31447 19128
rect 31389 19119 31447 19125
rect 32490 19116 32496 19128
rect 32548 19116 32554 19168
rect 34882 19116 34888 19168
rect 34940 19156 34946 19168
rect 35544 19156 35572 19184
rect 34940 19128 35572 19156
rect 38381 19159 38439 19165
rect 34940 19116 34946 19128
rect 38381 19125 38393 19159
rect 38427 19156 38439 19159
rect 39482 19156 39488 19168
rect 38427 19128 39488 19156
rect 38427 19125 38439 19128
rect 38381 19119 38439 19125
rect 39482 19116 39488 19128
rect 39540 19116 39546 19168
rect 40696 19156 40724 19264
rect 40788 19224 40816 19391
rect 40880 19292 40908 19468
rect 44913 19465 44925 19499
rect 44959 19496 44971 19499
rect 45462 19496 45468 19508
rect 44959 19468 45468 19496
rect 44959 19465 44971 19468
rect 44913 19459 44971 19465
rect 45462 19456 45468 19468
rect 45520 19456 45526 19508
rect 46385 19499 46443 19505
rect 46385 19496 46397 19499
rect 46032 19468 46397 19496
rect 41322 19388 41328 19440
rect 41380 19428 41386 19440
rect 46032 19428 46060 19468
rect 46385 19465 46397 19468
rect 46431 19465 46443 19499
rect 46385 19459 46443 19465
rect 46492 19468 46796 19496
rect 46492 19428 46520 19468
rect 41380 19400 45140 19428
rect 41380 19388 41386 19400
rect 40954 19320 40960 19372
rect 41012 19360 41018 19372
rect 42150 19360 42156 19372
rect 41012 19332 42156 19360
rect 41012 19320 41018 19332
rect 42150 19320 42156 19332
rect 42208 19320 42214 19372
rect 42886 19320 42892 19372
rect 42944 19360 42950 19372
rect 43714 19360 43720 19372
rect 42944 19332 43720 19360
rect 42944 19320 42950 19332
rect 43714 19320 43720 19332
rect 43772 19320 43778 19372
rect 41230 19292 41236 19304
rect 40880 19264 41236 19292
rect 41230 19252 41236 19264
rect 41288 19292 41294 19304
rect 41509 19295 41567 19301
rect 41509 19292 41521 19295
rect 41288 19264 41521 19292
rect 41288 19252 41294 19264
rect 41509 19261 41521 19264
rect 41555 19261 41567 19295
rect 41509 19255 41567 19261
rect 44358 19252 44364 19304
rect 44416 19252 44422 19304
rect 45112 19292 45140 19400
rect 45204 19400 46060 19428
rect 46400 19400 46520 19428
rect 45204 19369 45232 19400
rect 46400 19372 46428 19400
rect 46658 19388 46664 19440
rect 46716 19388 46722 19440
rect 46768 19437 46796 19468
rect 46934 19456 46940 19508
rect 46992 19456 46998 19508
rect 48038 19456 48044 19508
rect 48096 19496 48102 19508
rect 49326 19496 49332 19508
rect 48096 19468 49332 19496
rect 48096 19456 48102 19468
rect 49326 19456 49332 19468
rect 49384 19496 49390 19508
rect 49510 19496 49516 19508
rect 49384 19468 49516 19496
rect 49384 19456 49390 19468
rect 49510 19456 49516 19468
rect 49568 19456 49574 19508
rect 49878 19456 49884 19508
rect 49936 19496 49942 19508
rect 50062 19496 50068 19508
rect 49936 19468 50068 19496
rect 49936 19456 49942 19468
rect 50062 19456 50068 19468
rect 50120 19456 50126 19508
rect 52914 19456 52920 19508
rect 52972 19456 52978 19508
rect 54938 19456 54944 19508
rect 54996 19496 55002 19508
rect 55125 19499 55183 19505
rect 55125 19496 55137 19499
rect 54996 19468 55137 19496
rect 54996 19456 55002 19468
rect 55125 19465 55137 19468
rect 55171 19465 55183 19499
rect 55125 19459 55183 19465
rect 56689 19499 56747 19505
rect 56689 19465 56701 19499
rect 56735 19496 56747 19499
rect 56778 19496 56784 19508
rect 56735 19468 56784 19496
rect 56735 19465 56747 19468
rect 56689 19459 56747 19465
rect 56778 19456 56784 19468
rect 56836 19456 56842 19508
rect 46753 19431 46811 19437
rect 46753 19397 46765 19431
rect 46799 19397 46811 19431
rect 46952 19428 46980 19456
rect 50246 19428 50252 19440
rect 46753 19391 46811 19397
rect 46860 19400 46980 19428
rect 49068 19400 50252 19428
rect 45189 19363 45247 19369
rect 45189 19329 45201 19363
rect 45235 19329 45247 19363
rect 45373 19363 45431 19369
rect 45373 19360 45385 19363
rect 45189 19323 45247 19329
rect 45296 19332 45385 19360
rect 45296 19292 45324 19332
rect 45373 19329 45385 19332
rect 45419 19329 45431 19363
rect 45373 19323 45431 19329
rect 46201 19363 46259 19369
rect 46201 19329 46213 19363
rect 46247 19329 46259 19363
rect 46201 19323 46259 19329
rect 45112 19264 45324 19292
rect 45462 19252 45468 19304
rect 45520 19252 45526 19304
rect 46216 19292 46244 19323
rect 46382 19320 46388 19372
rect 46440 19320 46446 19372
rect 46564 19363 46622 19369
rect 46564 19329 46576 19363
rect 46610 19360 46622 19363
rect 46860 19360 46888 19400
rect 46610 19332 46888 19360
rect 46936 19363 46994 19369
rect 46610 19329 46622 19332
rect 46564 19323 46622 19329
rect 46936 19329 46948 19363
rect 46982 19329 46994 19363
rect 46936 19323 46994 19329
rect 46952 19292 46980 19323
rect 47026 19320 47032 19372
rect 47084 19320 47090 19372
rect 48593 19363 48651 19369
rect 48593 19329 48605 19363
rect 48639 19360 48651 19363
rect 48685 19363 48743 19369
rect 48685 19360 48697 19363
rect 48639 19332 48697 19360
rect 48639 19329 48651 19332
rect 48593 19323 48651 19329
rect 48685 19329 48697 19332
rect 48731 19329 48743 19363
rect 48685 19323 48743 19329
rect 48774 19320 48780 19372
rect 48832 19360 48838 19372
rect 49068 19369 49096 19400
rect 50246 19388 50252 19400
rect 50304 19388 50310 19440
rect 51350 19428 51356 19440
rect 51198 19400 51356 19428
rect 51350 19388 51356 19400
rect 51408 19388 51414 19440
rect 51442 19388 51448 19440
rect 51500 19428 51506 19440
rect 52825 19431 52883 19437
rect 52825 19428 52837 19431
rect 51500 19400 52837 19428
rect 51500 19388 51506 19400
rect 52825 19397 52837 19400
rect 52871 19397 52883 19431
rect 53926 19428 53932 19440
rect 52825 19391 52883 19397
rect 53392 19400 53932 19428
rect 53392 19369 53420 19400
rect 53926 19388 53932 19400
rect 53984 19388 53990 19440
rect 54110 19388 54116 19440
rect 54168 19388 54174 19440
rect 56796 19428 56824 19456
rect 56796 19400 57100 19428
rect 48961 19363 49019 19369
rect 48961 19360 48973 19363
rect 48832 19332 48973 19360
rect 48832 19320 48838 19332
rect 48961 19329 48973 19332
rect 49007 19329 49019 19363
rect 48961 19323 49019 19329
rect 49053 19363 49111 19369
rect 49053 19329 49065 19363
rect 49099 19329 49111 19363
rect 49053 19323 49111 19329
rect 53377 19363 53435 19369
rect 53377 19329 53389 19363
rect 53423 19329 53435 19363
rect 53377 19323 53435 19329
rect 56594 19320 56600 19372
rect 56652 19360 56658 19372
rect 57072 19369 57100 19400
rect 56781 19363 56839 19369
rect 56781 19360 56793 19363
rect 56652 19332 56793 19360
rect 56652 19320 56658 19332
rect 56781 19329 56793 19332
rect 56827 19329 56839 19363
rect 56781 19323 56839 19329
rect 56965 19363 57023 19369
rect 56965 19329 56977 19363
rect 57011 19329 57023 19363
rect 56965 19323 57023 19329
rect 57057 19363 57115 19369
rect 57057 19329 57069 19363
rect 57103 19329 57115 19363
rect 57057 19323 57115 19329
rect 57149 19363 57207 19369
rect 57149 19329 57161 19363
rect 57195 19360 57207 19363
rect 57885 19363 57943 19369
rect 57885 19360 57897 19363
rect 57195 19332 57897 19360
rect 57195 19329 57207 19332
rect 57149 19323 57207 19329
rect 57885 19329 57897 19332
rect 57931 19329 57943 19363
rect 57885 19323 57943 19329
rect 47118 19292 47124 19304
rect 46216 19264 46888 19292
rect 46952 19264 47124 19292
rect 41138 19224 41144 19236
rect 40788 19196 41144 19224
rect 41138 19184 41144 19196
rect 41196 19224 41202 19236
rect 41877 19227 41935 19233
rect 41877 19224 41889 19227
rect 41196 19196 41889 19224
rect 41196 19184 41202 19196
rect 41877 19193 41889 19196
rect 41923 19224 41935 19227
rect 46216 19224 46244 19264
rect 46860 19236 46888 19264
rect 47118 19252 47124 19264
rect 47176 19292 47182 19304
rect 48041 19295 48099 19301
rect 48041 19292 48053 19295
rect 47176 19264 48053 19292
rect 47176 19252 47182 19264
rect 48041 19261 48053 19264
rect 48087 19292 48099 19295
rect 49418 19292 49424 19304
rect 48087 19264 49424 19292
rect 48087 19261 48099 19264
rect 48041 19255 48099 19261
rect 49418 19252 49424 19264
rect 49476 19252 49482 19304
rect 49694 19252 49700 19304
rect 49752 19252 49758 19304
rect 49970 19252 49976 19304
rect 50028 19252 50034 19304
rect 51166 19252 51172 19304
rect 51224 19292 51230 19304
rect 51445 19295 51503 19301
rect 51445 19292 51457 19295
rect 51224 19264 51457 19292
rect 51224 19252 51230 19264
rect 51445 19261 51457 19264
rect 51491 19292 51503 19295
rect 52089 19295 52147 19301
rect 52089 19292 52101 19295
rect 51491 19264 52101 19292
rect 51491 19261 51503 19264
rect 51445 19255 51503 19261
rect 52089 19261 52101 19264
rect 52135 19261 52147 19295
rect 52089 19255 52147 19261
rect 53650 19252 53656 19304
rect 53708 19252 53714 19304
rect 56980 19292 57008 19323
rect 56980 19264 57100 19292
rect 57072 19236 57100 19264
rect 58250 19252 58256 19304
rect 58308 19292 58314 19304
rect 58437 19295 58495 19301
rect 58437 19292 58449 19295
rect 58308 19264 58449 19292
rect 58308 19252 58314 19264
rect 58437 19261 58449 19264
rect 58483 19261 58495 19295
rect 58437 19255 58495 19261
rect 41923 19196 46244 19224
rect 41923 19193 41935 19196
rect 41877 19187 41935 19193
rect 46842 19184 46848 19236
rect 46900 19224 46906 19236
rect 47305 19227 47363 19233
rect 47305 19224 47317 19227
rect 46900 19196 47317 19224
rect 46900 19184 46906 19196
rect 47305 19193 47317 19196
rect 47351 19193 47363 19227
rect 47305 19187 47363 19193
rect 47394 19184 47400 19236
rect 47452 19224 47458 19236
rect 47762 19224 47768 19236
rect 47452 19196 47768 19224
rect 47452 19184 47458 19196
rect 47762 19184 47768 19196
rect 47820 19184 47826 19236
rect 48777 19227 48835 19233
rect 48777 19193 48789 19227
rect 48823 19224 48835 19227
rect 49602 19224 49608 19236
rect 48823 19196 49608 19224
rect 48823 19193 48835 19196
rect 48777 19187 48835 19193
rect 49602 19184 49608 19196
rect 49660 19184 49666 19236
rect 57054 19184 57060 19236
rect 57112 19184 57118 19236
rect 40954 19156 40960 19168
rect 40696 19128 40960 19156
rect 40954 19116 40960 19128
rect 41012 19116 41018 19168
rect 45005 19159 45063 19165
rect 45005 19125 45017 19159
rect 45051 19156 45063 19159
rect 45278 19156 45284 19168
rect 45051 19128 45284 19156
rect 45051 19125 45063 19128
rect 45005 19119 45063 19125
rect 45278 19116 45284 19128
rect 45336 19116 45342 19168
rect 47026 19116 47032 19168
rect 47084 19156 47090 19168
rect 47121 19159 47179 19165
rect 47121 19156 47133 19159
rect 47084 19128 47133 19156
rect 47084 19116 47090 19128
rect 47121 19125 47133 19128
rect 47167 19125 47179 19159
rect 47121 19119 47179 19125
rect 47486 19116 47492 19168
rect 47544 19156 47550 19168
rect 47581 19159 47639 19165
rect 47581 19156 47593 19159
rect 47544 19128 47593 19156
rect 47544 19116 47550 19128
rect 47581 19125 47593 19128
rect 47627 19125 47639 19159
rect 47780 19156 47808 19184
rect 49142 19156 49148 19168
rect 47780 19128 49148 19156
rect 47581 19119 47639 19125
rect 49142 19116 49148 19128
rect 49200 19116 49206 19168
rect 49234 19116 49240 19168
rect 49292 19116 49298 19168
rect 51534 19116 51540 19168
rect 51592 19116 51598 19168
rect 57422 19116 57428 19168
rect 57480 19116 57486 19168
rect 1104 19066 58880 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 58880 19066
rect 1104 18992 58880 19014
rect 16114 18912 16120 18964
rect 16172 18912 16178 18964
rect 16850 18912 16856 18964
rect 16908 18912 16914 18964
rect 25041 18955 25099 18961
rect 25041 18921 25053 18955
rect 25087 18952 25099 18955
rect 25314 18952 25320 18964
rect 25087 18924 25320 18952
rect 25087 18921 25099 18924
rect 25041 18915 25099 18921
rect 25314 18912 25320 18924
rect 25372 18912 25378 18964
rect 25869 18955 25927 18961
rect 25869 18921 25881 18955
rect 25915 18952 25927 18955
rect 26970 18952 26976 18964
rect 25915 18924 26976 18952
rect 25915 18921 25927 18924
rect 25869 18915 25927 18921
rect 26970 18912 26976 18924
rect 27028 18912 27034 18964
rect 30374 18952 30380 18964
rect 27092 18924 30380 18952
rect 15194 18776 15200 18828
rect 15252 18816 15258 18828
rect 15381 18819 15439 18825
rect 15381 18816 15393 18819
rect 15252 18788 15393 18816
rect 15252 18776 15258 18788
rect 15381 18785 15393 18788
rect 15427 18785 15439 18819
rect 16868 18816 16896 18912
rect 19610 18844 19616 18896
rect 19668 18884 19674 18896
rect 20070 18884 20076 18896
rect 19668 18856 20076 18884
rect 19668 18844 19674 18856
rect 20070 18844 20076 18856
rect 20128 18844 20134 18896
rect 25130 18884 25136 18896
rect 24044 18856 25136 18884
rect 15381 18779 15439 18785
rect 16500 18788 16896 18816
rect 16500 18757 16528 18788
rect 17586 18776 17592 18828
rect 17644 18776 17650 18828
rect 19061 18819 19119 18825
rect 19061 18785 19073 18819
rect 19107 18816 19119 18819
rect 19518 18816 19524 18828
rect 19107 18788 19524 18816
rect 19107 18785 19119 18788
rect 19061 18779 19119 18785
rect 19518 18776 19524 18788
rect 19576 18816 19582 18828
rect 19576 18788 19748 18816
rect 19576 18776 19582 18788
rect 16025 18751 16083 18757
rect 16025 18717 16037 18751
rect 16071 18748 16083 18751
rect 16393 18751 16451 18757
rect 16393 18748 16405 18751
rect 16071 18720 16405 18748
rect 16071 18717 16083 18720
rect 16025 18711 16083 18717
rect 16393 18717 16405 18720
rect 16439 18717 16451 18751
rect 16393 18711 16451 18717
rect 16485 18751 16543 18757
rect 16485 18717 16497 18751
rect 16531 18717 16543 18751
rect 16485 18711 16543 18717
rect 16577 18751 16635 18757
rect 16577 18717 16589 18751
rect 16623 18717 16635 18751
rect 16577 18711 16635 18717
rect 16592 18680 16620 18711
rect 16758 18708 16764 18760
rect 16816 18708 16822 18760
rect 17310 18708 17316 18760
rect 17368 18708 17374 18760
rect 19720 18757 19748 18788
rect 20088 18757 20116 18844
rect 21910 18776 21916 18828
rect 21968 18776 21974 18828
rect 22554 18776 22560 18828
rect 22612 18776 22618 18828
rect 23014 18776 23020 18828
rect 23072 18816 23078 18828
rect 23290 18816 23296 18828
rect 23072 18788 23296 18816
rect 23072 18776 23078 18788
rect 23290 18776 23296 18788
rect 23348 18816 23354 18828
rect 24044 18825 24072 18856
rect 25130 18844 25136 18856
rect 25188 18844 25194 18896
rect 27092 18884 27120 18924
rect 30374 18912 30380 18924
rect 30432 18912 30438 18964
rect 30558 18912 30564 18964
rect 30616 18912 30622 18964
rect 34514 18912 34520 18964
rect 34572 18912 34578 18964
rect 34885 18955 34943 18961
rect 34885 18921 34897 18955
rect 34931 18952 34943 18955
rect 35526 18952 35532 18964
rect 34931 18924 35532 18952
rect 34931 18921 34943 18924
rect 34885 18915 34943 18921
rect 35526 18912 35532 18924
rect 35584 18912 35590 18964
rect 39206 18912 39212 18964
rect 39264 18952 39270 18964
rect 39669 18955 39727 18961
rect 39669 18952 39681 18955
rect 39264 18924 39681 18952
rect 39264 18912 39270 18924
rect 39669 18921 39681 18924
rect 39715 18952 39727 18955
rect 39758 18952 39764 18964
rect 39715 18924 39764 18952
rect 39715 18921 39727 18924
rect 39669 18915 39727 18921
rect 39758 18912 39764 18924
rect 39816 18912 39822 18964
rect 39850 18912 39856 18964
rect 39908 18952 39914 18964
rect 39908 18924 46704 18952
rect 39908 18912 39914 18924
rect 34330 18884 34336 18896
rect 25744 18856 27120 18884
rect 27264 18856 27752 18884
rect 24029 18819 24087 18825
rect 24029 18816 24041 18819
rect 23348 18788 24041 18816
rect 23348 18776 23354 18788
rect 24029 18785 24041 18788
rect 24075 18785 24087 18819
rect 24946 18816 24952 18828
rect 24029 18779 24087 18785
rect 24688 18788 24952 18816
rect 19613 18751 19671 18757
rect 19613 18748 19625 18751
rect 19536 18720 19625 18748
rect 19536 18692 19564 18720
rect 19613 18717 19625 18720
rect 19659 18717 19671 18751
rect 19613 18711 19671 18717
rect 19706 18751 19764 18757
rect 19706 18717 19718 18751
rect 19752 18717 19764 18751
rect 19706 18711 19764 18717
rect 20078 18751 20136 18757
rect 20078 18717 20090 18751
rect 20124 18717 20136 18751
rect 20078 18711 20136 18717
rect 22186 18708 22192 18760
rect 22244 18748 22250 18760
rect 22281 18751 22339 18757
rect 22281 18748 22293 18751
rect 22244 18720 22293 18748
rect 22244 18708 22250 18720
rect 22281 18717 22293 18720
rect 22327 18717 22339 18751
rect 22281 18711 22339 18717
rect 24394 18708 24400 18760
rect 24452 18748 24458 18760
rect 24688 18757 24716 18788
rect 24946 18776 24952 18788
rect 25004 18776 25010 18828
rect 25744 18816 25772 18856
rect 26602 18816 26608 18828
rect 25240 18788 25772 18816
rect 26252 18788 26608 18816
rect 24489 18751 24547 18757
rect 24489 18748 24501 18751
rect 24452 18720 24501 18748
rect 24452 18708 24458 18720
rect 24489 18717 24501 18720
rect 24535 18717 24547 18751
rect 24489 18711 24547 18717
rect 24673 18751 24731 18757
rect 24673 18717 24685 18751
rect 24719 18717 24731 18751
rect 24673 18711 24731 18717
rect 24857 18751 24915 18757
rect 24857 18717 24869 18751
rect 24903 18748 24915 18751
rect 25038 18748 25044 18760
rect 24903 18720 25044 18748
rect 24903 18717 24915 18720
rect 24857 18711 24915 18717
rect 16592 18652 18000 18680
rect 18814 18652 18920 18680
rect 17972 18624 18000 18652
rect 17954 18572 17960 18624
rect 18012 18572 18018 18624
rect 18892 18612 18920 18652
rect 19518 18640 19524 18692
rect 19576 18640 19582 18692
rect 19889 18683 19947 18689
rect 19889 18649 19901 18683
rect 19935 18649 19947 18683
rect 19889 18643 19947 18649
rect 19981 18683 20039 18689
rect 19981 18649 19993 18683
rect 20027 18680 20039 18683
rect 21910 18680 21916 18692
rect 20027 18652 20484 18680
rect 21482 18652 21916 18680
rect 20027 18649 20039 18652
rect 19981 18643 20039 18649
rect 19610 18612 19616 18624
rect 18892 18584 19616 18612
rect 19610 18572 19616 18584
rect 19668 18572 19674 18624
rect 19702 18572 19708 18624
rect 19760 18612 19766 18624
rect 19904 18612 19932 18643
rect 19760 18584 19932 18612
rect 19760 18572 19766 18584
rect 20254 18572 20260 18624
rect 20312 18572 20318 18624
rect 20456 18621 20484 18652
rect 21910 18640 21916 18652
rect 21968 18680 21974 18692
rect 21968 18652 23046 18680
rect 21968 18640 21974 18652
rect 24762 18640 24768 18692
rect 24820 18640 24826 18692
rect 20441 18615 20499 18621
rect 20441 18581 20453 18615
rect 20487 18612 20499 18615
rect 22370 18612 22376 18624
rect 20487 18584 22376 18612
rect 20487 18581 20499 18584
rect 20441 18575 20499 18581
rect 22370 18572 22376 18584
rect 22428 18612 22434 18624
rect 23842 18612 23848 18624
rect 22428 18584 23848 18612
rect 22428 18572 22434 18584
rect 23842 18572 23848 18584
rect 23900 18572 23906 18624
rect 24578 18572 24584 18624
rect 24636 18612 24642 18624
rect 24872 18612 24900 18711
rect 25038 18708 25044 18720
rect 25096 18708 25102 18760
rect 25240 18757 25268 18788
rect 25225 18751 25283 18757
rect 25225 18717 25237 18751
rect 25271 18717 25283 18751
rect 25225 18711 25283 18717
rect 25318 18751 25376 18757
rect 25318 18717 25330 18751
rect 25364 18717 25376 18751
rect 25318 18711 25376 18717
rect 25130 18640 25136 18692
rect 25188 18680 25194 18692
rect 25332 18680 25360 18711
rect 25406 18708 25412 18760
rect 25464 18748 25470 18760
rect 25501 18751 25559 18757
rect 25501 18748 25513 18751
rect 25464 18720 25513 18748
rect 25464 18708 25470 18720
rect 25501 18717 25513 18720
rect 25547 18717 25559 18751
rect 25501 18711 25559 18717
rect 25690 18751 25748 18757
rect 25690 18717 25702 18751
rect 25736 18717 25748 18751
rect 25690 18711 25748 18717
rect 25188 18652 25360 18680
rect 25593 18683 25651 18689
rect 25188 18640 25194 18652
rect 25593 18649 25605 18683
rect 25639 18649 25651 18683
rect 25593 18643 25651 18649
rect 24636 18584 24900 18612
rect 24636 18572 24642 18584
rect 25038 18572 25044 18624
rect 25096 18612 25102 18624
rect 25608 18612 25636 18643
rect 25096 18584 25636 18612
rect 25700 18612 25728 18711
rect 25866 18708 25872 18760
rect 25924 18748 25930 18760
rect 25961 18751 26019 18757
rect 25961 18748 25973 18751
rect 25924 18720 25973 18748
rect 25924 18708 25930 18720
rect 25961 18717 25973 18720
rect 26007 18717 26019 18751
rect 25961 18711 26019 18717
rect 26099 18751 26157 18757
rect 26099 18717 26111 18751
rect 26145 18748 26157 18751
rect 26252 18748 26280 18788
rect 26602 18776 26608 18788
rect 26660 18776 26666 18828
rect 26418 18748 26424 18760
rect 26476 18757 26482 18760
rect 27264 18757 27292 18856
rect 27614 18776 27620 18828
rect 27672 18776 27678 18828
rect 27724 18816 27752 18856
rect 34164 18856 34336 18884
rect 28626 18816 28632 18828
rect 27724 18788 28632 18816
rect 28626 18776 28632 18788
rect 28684 18816 28690 18828
rect 30558 18816 30564 18828
rect 28684 18788 30052 18816
rect 28684 18776 28690 18788
rect 26145 18720 26280 18748
rect 26384 18720 26424 18748
rect 26145 18717 26157 18720
rect 26099 18711 26157 18717
rect 26418 18708 26424 18720
rect 26476 18711 26484 18757
rect 26973 18751 27031 18757
rect 26973 18717 26985 18751
rect 27019 18717 27031 18751
rect 26973 18711 27031 18717
rect 27249 18751 27307 18757
rect 27249 18717 27261 18751
rect 27295 18717 27307 18751
rect 27249 18711 27307 18717
rect 26476 18708 26482 18711
rect 26237 18683 26295 18689
rect 26237 18649 26249 18683
rect 26283 18649 26295 18683
rect 26237 18643 26295 18649
rect 25958 18612 25964 18624
rect 25700 18584 25964 18612
rect 25096 18572 25102 18584
rect 25958 18572 25964 18584
rect 26016 18572 26022 18624
rect 26142 18572 26148 18624
rect 26200 18612 26206 18624
rect 26252 18612 26280 18643
rect 26326 18640 26332 18692
rect 26384 18640 26390 18692
rect 26988 18680 27016 18711
rect 27338 18708 27344 18760
rect 27396 18708 27402 18760
rect 30024 18757 30052 18788
rect 30208 18788 30564 18816
rect 30208 18757 30236 18788
rect 30558 18776 30564 18788
rect 30616 18776 30622 18828
rect 31662 18776 31668 18828
rect 31720 18816 31726 18828
rect 32401 18819 32459 18825
rect 32401 18816 32413 18819
rect 31720 18788 32413 18816
rect 31720 18776 31726 18788
rect 32401 18785 32413 18788
rect 32447 18785 32459 18819
rect 32401 18779 32459 18785
rect 34054 18776 34060 18828
rect 34112 18776 34118 18828
rect 30009 18751 30067 18757
rect 30009 18717 30021 18751
rect 30055 18717 30067 18751
rect 30009 18711 30067 18717
rect 30193 18751 30251 18757
rect 30193 18717 30205 18751
rect 30239 18717 30251 18751
rect 30193 18711 30251 18717
rect 26436 18652 27016 18680
rect 27157 18683 27215 18689
rect 26436 18624 26464 18652
rect 27157 18649 27169 18683
rect 27203 18649 27215 18683
rect 27157 18643 27215 18649
rect 27893 18683 27951 18689
rect 27893 18649 27905 18683
rect 27939 18680 27951 18683
rect 27982 18680 27988 18692
rect 27939 18652 27988 18680
rect 27939 18649 27951 18652
rect 27893 18643 27951 18649
rect 26200 18584 26280 18612
rect 26200 18572 26206 18584
rect 26418 18572 26424 18624
rect 26476 18572 26482 18624
rect 26602 18572 26608 18624
rect 26660 18572 26666 18624
rect 26786 18572 26792 18624
rect 26844 18572 26850 18624
rect 26970 18572 26976 18624
rect 27028 18612 27034 18624
rect 27172 18612 27200 18643
rect 27982 18640 27988 18652
rect 28040 18640 28046 18692
rect 28902 18640 28908 18692
rect 28960 18640 28966 18692
rect 27338 18612 27344 18624
rect 27028 18584 27344 18612
rect 27028 18572 27034 18584
rect 27338 18572 27344 18584
rect 27396 18572 27402 18624
rect 27525 18615 27583 18621
rect 27525 18581 27537 18615
rect 27571 18612 27583 18615
rect 28258 18612 28264 18624
rect 27571 18584 28264 18612
rect 27571 18581 27583 18584
rect 27525 18575 27583 18581
rect 28258 18572 28264 18584
rect 28316 18572 28322 18624
rect 29362 18572 29368 18624
rect 29420 18572 29426 18624
rect 30024 18612 30052 18711
rect 30282 18708 30288 18760
rect 30340 18708 30346 18760
rect 30377 18751 30435 18757
rect 30377 18717 30389 18751
rect 30423 18748 30435 18751
rect 30742 18748 30748 18760
rect 30423 18720 30748 18748
rect 30423 18717 30435 18720
rect 30377 18711 30435 18717
rect 30742 18708 30748 18720
rect 30800 18708 30806 18760
rect 33965 18751 34023 18757
rect 33965 18717 33977 18751
rect 34011 18748 34023 18751
rect 34164 18748 34192 18856
rect 34330 18844 34336 18856
rect 34388 18844 34394 18896
rect 39482 18844 39488 18896
rect 39540 18884 39546 18896
rect 41322 18884 41328 18896
rect 39540 18856 41328 18884
rect 39540 18844 39546 18856
rect 41322 18844 41328 18856
rect 41380 18844 41386 18896
rect 46676 18884 46704 18924
rect 46750 18912 46756 18964
rect 46808 18912 46814 18964
rect 47118 18912 47124 18964
rect 47176 18912 47182 18964
rect 48406 18912 48412 18964
rect 48464 18952 48470 18964
rect 49050 18952 49056 18964
rect 48464 18924 49056 18952
rect 48464 18912 48470 18924
rect 49050 18912 49056 18924
rect 49108 18912 49114 18964
rect 49694 18952 49700 18964
rect 49344 18924 49700 18952
rect 47394 18884 47400 18896
rect 46676 18856 47400 18884
rect 47394 18844 47400 18856
rect 47452 18844 47458 18896
rect 49234 18884 49240 18896
rect 48792 18856 49240 18884
rect 34606 18816 34612 18828
rect 34256 18788 34612 18816
rect 34256 18757 34284 18788
rect 34606 18776 34612 18788
rect 34664 18776 34670 18828
rect 37918 18776 37924 18828
rect 37976 18776 37982 18828
rect 45278 18776 45284 18828
rect 45336 18776 45342 18828
rect 48593 18819 48651 18825
rect 48593 18785 48605 18819
rect 48639 18816 48651 18819
rect 48792 18816 48820 18856
rect 49234 18844 49240 18856
rect 49292 18844 49298 18896
rect 48639 18788 48820 18816
rect 48869 18819 48927 18825
rect 48639 18785 48651 18788
rect 48593 18779 48651 18785
rect 48869 18785 48881 18819
rect 48915 18816 48927 18819
rect 49344 18816 49372 18924
rect 49694 18912 49700 18924
rect 49752 18912 49758 18964
rect 49970 18912 49976 18964
rect 50028 18952 50034 18964
rect 50157 18955 50215 18961
rect 50157 18952 50169 18955
rect 50028 18924 50169 18952
rect 50028 18912 50034 18924
rect 50157 18921 50169 18924
rect 50203 18921 50215 18955
rect 50157 18915 50215 18921
rect 51629 18955 51687 18961
rect 51629 18921 51641 18955
rect 51675 18952 51687 18955
rect 51718 18952 51724 18964
rect 51675 18924 51724 18952
rect 51675 18921 51687 18924
rect 51629 18915 51687 18921
rect 51718 18912 51724 18924
rect 51776 18912 51782 18964
rect 52546 18912 52552 18964
rect 52604 18952 52610 18964
rect 53193 18955 53251 18961
rect 53193 18952 53205 18955
rect 52604 18924 53205 18952
rect 52604 18912 52610 18924
rect 53193 18921 53205 18924
rect 53239 18952 53251 18955
rect 53282 18952 53288 18964
rect 53239 18924 53288 18952
rect 53239 18921 53251 18924
rect 53193 18915 53251 18921
rect 53282 18912 53288 18924
rect 53340 18952 53346 18964
rect 54110 18952 54116 18964
rect 53340 18924 54116 18952
rect 53340 18912 53346 18924
rect 54110 18912 54116 18924
rect 54168 18912 54174 18964
rect 58250 18912 58256 18964
rect 58308 18912 58314 18964
rect 49513 18887 49571 18893
rect 49513 18853 49525 18887
rect 49559 18853 49571 18887
rect 49513 18847 49571 18853
rect 48915 18788 49372 18816
rect 48915 18785 48927 18788
rect 48869 18779 48927 18785
rect 34011 18720 34192 18748
rect 34241 18751 34299 18757
rect 34011 18717 34023 18720
rect 33965 18711 34023 18717
rect 34241 18717 34253 18751
rect 34287 18717 34299 18751
rect 34241 18711 34299 18717
rect 34333 18751 34391 18757
rect 34333 18717 34345 18751
rect 34379 18748 34391 18751
rect 34698 18748 34704 18760
rect 34379 18720 34704 18748
rect 34379 18717 34391 18720
rect 34333 18711 34391 18717
rect 34698 18708 34704 18720
rect 34756 18708 34762 18760
rect 34790 18708 34796 18760
rect 34848 18748 34854 18760
rect 35161 18751 35219 18757
rect 35161 18748 35173 18751
rect 34848 18720 35173 18748
rect 34848 18708 34854 18720
rect 35161 18717 35173 18720
rect 35207 18748 35219 18751
rect 37090 18748 37096 18760
rect 35207 18720 37096 18748
rect 35207 18717 35219 18720
rect 35161 18711 35219 18717
rect 37090 18708 37096 18720
rect 37148 18708 37154 18760
rect 39758 18708 39764 18760
rect 39816 18748 39822 18760
rect 40405 18751 40463 18757
rect 40405 18748 40417 18751
rect 39816 18720 40417 18748
rect 39816 18708 39822 18720
rect 40405 18717 40417 18720
rect 40451 18748 40463 18751
rect 40494 18748 40500 18760
rect 40451 18720 40500 18748
rect 40451 18717 40463 18720
rect 40405 18711 40463 18717
rect 40494 18708 40500 18720
rect 40552 18708 40558 18760
rect 41230 18708 41236 18760
rect 41288 18748 41294 18760
rect 45002 18748 45008 18760
rect 41288 18720 45008 18748
rect 41288 18708 41294 18720
rect 45002 18708 45008 18720
rect 45060 18708 45066 18760
rect 48958 18708 48964 18760
rect 49016 18708 49022 18760
rect 49050 18708 49056 18760
rect 49108 18748 49114 18760
rect 49329 18751 49387 18757
rect 49329 18748 49341 18751
rect 49108 18720 49341 18748
rect 49108 18708 49114 18720
rect 49329 18717 49341 18720
rect 49375 18717 49387 18751
rect 49329 18711 49387 18717
rect 30300 18680 30328 18708
rect 30834 18680 30840 18692
rect 30300 18652 30840 18680
rect 30834 18640 30840 18652
rect 30892 18640 30898 18692
rect 31386 18640 31392 18692
rect 31444 18640 31450 18692
rect 32122 18640 32128 18692
rect 32180 18640 32186 18692
rect 36725 18683 36783 18689
rect 36725 18649 36737 18683
rect 36771 18680 36783 18683
rect 36771 18652 36860 18680
rect 36771 18649 36783 18652
rect 36725 18643 36783 18649
rect 36832 18624 36860 18652
rect 38194 18640 38200 18692
rect 38252 18640 38258 18692
rect 38286 18640 38292 18692
rect 38344 18680 38350 18692
rect 38344 18652 38686 18680
rect 38344 18640 38350 18652
rect 39574 18640 39580 18692
rect 39632 18680 39638 18692
rect 39853 18683 39911 18689
rect 39853 18680 39865 18683
rect 39632 18652 39865 18680
rect 39632 18640 39638 18652
rect 39853 18649 39865 18652
rect 39899 18649 39911 18683
rect 39853 18643 39911 18649
rect 44082 18640 44088 18692
rect 44140 18680 44146 18692
rect 44140 18652 45770 18680
rect 44140 18640 44146 18652
rect 47854 18640 47860 18692
rect 47912 18640 47918 18692
rect 48314 18640 48320 18692
rect 48372 18680 48378 18692
rect 49145 18683 49203 18689
rect 49145 18680 49157 18683
rect 48372 18652 49157 18680
rect 48372 18640 48378 18652
rect 49145 18649 49157 18652
rect 49191 18649 49203 18683
rect 49145 18643 49203 18649
rect 49237 18683 49295 18689
rect 49237 18649 49249 18683
rect 49283 18680 49295 18683
rect 49418 18680 49424 18692
rect 49283 18652 49424 18680
rect 49283 18649 49295 18652
rect 49237 18643 49295 18649
rect 49418 18640 49424 18652
rect 49476 18640 49482 18692
rect 49528 18680 49556 18847
rect 49602 18844 49608 18896
rect 49660 18884 49666 18896
rect 50617 18887 50675 18893
rect 50617 18884 50629 18887
rect 49660 18856 50629 18884
rect 49660 18844 49666 18856
rect 50617 18853 50629 18856
rect 50663 18853 50675 18887
rect 50617 18847 50675 18853
rect 50338 18708 50344 18760
rect 50396 18708 50402 18760
rect 50433 18751 50491 18757
rect 50433 18717 50445 18751
rect 50479 18717 50491 18751
rect 50433 18711 50491 18717
rect 50448 18680 50476 18711
rect 49528 18652 50476 18680
rect 50632 18680 50660 18847
rect 51997 18819 52055 18825
rect 51997 18785 52009 18819
rect 52043 18816 52055 18819
rect 53834 18816 53840 18828
rect 52043 18788 53840 18816
rect 52043 18785 52055 18788
rect 51997 18779 52055 18785
rect 53834 18776 53840 18788
rect 53892 18776 53898 18828
rect 50709 18751 50767 18757
rect 50709 18717 50721 18751
rect 50755 18748 50767 18751
rect 51534 18748 51540 18760
rect 50755 18720 51540 18748
rect 50755 18717 50767 18720
rect 50709 18711 50767 18717
rect 51534 18708 51540 18720
rect 51592 18708 51598 18760
rect 51810 18708 51816 18760
rect 51868 18708 51874 18760
rect 52086 18708 52092 18760
rect 52144 18708 52150 18760
rect 56870 18708 56876 18760
rect 56928 18708 56934 18760
rect 57140 18751 57198 18757
rect 57140 18717 57152 18751
rect 57186 18748 57198 18751
rect 57422 18748 57428 18760
rect 57186 18720 57428 18748
rect 57186 18717 57198 18720
rect 57140 18711 57198 18717
rect 57422 18708 57428 18720
rect 57480 18708 57486 18760
rect 51074 18680 51080 18692
rect 50632 18652 51080 18680
rect 51074 18640 51080 18652
rect 51132 18640 51138 18692
rect 30653 18615 30711 18621
rect 30653 18612 30665 18615
rect 30024 18584 30665 18612
rect 30653 18581 30665 18584
rect 30699 18612 30711 18615
rect 31110 18612 31116 18624
rect 30699 18584 31116 18612
rect 30699 18581 30711 18584
rect 30653 18575 30711 18581
rect 31110 18572 31116 18584
rect 31168 18572 31174 18624
rect 36814 18572 36820 18624
rect 36872 18572 36878 18624
rect 37090 18572 37096 18624
rect 37148 18612 37154 18624
rect 40862 18612 40868 18624
rect 37148 18584 40868 18612
rect 37148 18572 37154 18584
rect 40862 18572 40868 18584
rect 40920 18572 40926 18624
rect 48958 18572 48964 18624
rect 49016 18612 49022 18624
rect 52104 18612 52132 18708
rect 49016 18584 52132 18612
rect 49016 18572 49022 18584
rect 1104 18522 58880 18544
rect 1104 18470 4874 18522
rect 4926 18470 4938 18522
rect 4990 18470 5002 18522
rect 5054 18470 5066 18522
rect 5118 18470 5130 18522
rect 5182 18470 35594 18522
rect 35646 18470 35658 18522
rect 35710 18470 35722 18522
rect 35774 18470 35786 18522
rect 35838 18470 35850 18522
rect 35902 18470 58880 18522
rect 1104 18448 58880 18470
rect 19886 18368 19892 18420
rect 19944 18408 19950 18420
rect 19981 18411 20039 18417
rect 19981 18408 19993 18411
rect 19944 18380 19993 18408
rect 19944 18368 19950 18380
rect 19981 18377 19993 18380
rect 20027 18408 20039 18411
rect 20027 18380 20576 18408
rect 20027 18377 20039 18380
rect 19981 18371 20039 18377
rect 20548 18284 20576 18380
rect 21818 18368 21824 18420
rect 21876 18408 21882 18420
rect 21913 18411 21971 18417
rect 21913 18408 21925 18411
rect 21876 18380 21925 18408
rect 21876 18368 21882 18380
rect 21913 18377 21925 18380
rect 21959 18377 21971 18411
rect 23014 18408 23020 18420
rect 21913 18371 21971 18377
rect 22204 18380 23020 18408
rect 16574 18232 16580 18284
rect 16632 18272 16638 18284
rect 16669 18275 16727 18281
rect 16669 18272 16681 18275
rect 16632 18244 16681 18272
rect 16632 18232 16638 18244
rect 16669 18241 16681 18244
rect 16715 18272 16727 18275
rect 17681 18275 17739 18281
rect 17681 18272 17693 18275
rect 16715 18244 17693 18272
rect 16715 18241 16727 18244
rect 16669 18235 16727 18241
rect 17681 18241 17693 18244
rect 17727 18272 17739 18275
rect 18138 18272 18144 18284
rect 17727 18244 18144 18272
rect 17727 18241 17739 18244
rect 17681 18235 17739 18241
rect 18138 18232 18144 18244
rect 18196 18232 18202 18284
rect 19610 18232 19616 18284
rect 19668 18272 19674 18284
rect 19668 18244 20208 18272
rect 19668 18232 19674 18244
rect 17310 18204 17316 18216
rect 16684 18176 17316 18204
rect 16684 18148 16712 18176
rect 17310 18164 17316 18176
rect 17368 18204 17374 18216
rect 17405 18207 17463 18213
rect 17405 18204 17417 18207
rect 17368 18176 17417 18204
rect 17368 18164 17374 18176
rect 17405 18173 17417 18176
rect 17451 18204 17463 18207
rect 18233 18207 18291 18213
rect 18233 18204 18245 18207
rect 17451 18176 18245 18204
rect 17451 18173 17463 18176
rect 17405 18167 17463 18173
rect 18233 18173 18245 18176
rect 18279 18173 18291 18207
rect 18233 18167 18291 18173
rect 18509 18207 18567 18213
rect 18509 18173 18521 18207
rect 18555 18204 18567 18207
rect 20073 18207 20131 18213
rect 20073 18204 20085 18207
rect 18555 18176 20085 18204
rect 18555 18173 18567 18176
rect 18509 18167 18567 18173
rect 20073 18173 20085 18176
rect 20119 18173 20131 18207
rect 20180 18204 20208 18244
rect 20254 18232 20260 18284
rect 20312 18232 20318 18284
rect 20530 18232 20536 18284
rect 20588 18232 20594 18284
rect 22204 18281 22232 18380
rect 23014 18368 23020 18380
rect 23072 18368 23078 18420
rect 23106 18368 23112 18420
rect 23164 18408 23170 18420
rect 23201 18411 23259 18417
rect 23201 18408 23213 18411
rect 23164 18380 23213 18408
rect 23164 18368 23170 18380
rect 23201 18377 23213 18380
rect 23247 18377 23259 18411
rect 23201 18371 23259 18377
rect 24670 18368 24676 18420
rect 24728 18408 24734 18420
rect 24946 18408 24952 18420
rect 24728 18380 24952 18408
rect 24728 18368 24734 18380
rect 24946 18368 24952 18380
rect 25004 18368 25010 18420
rect 28902 18408 28908 18420
rect 26252 18380 28908 18408
rect 24762 18340 24768 18352
rect 22480 18312 24768 18340
rect 22480 18284 22508 18312
rect 24762 18300 24768 18312
rect 24820 18300 24826 18352
rect 26252 18340 26280 18380
rect 28902 18368 28908 18380
rect 28960 18368 28966 18420
rect 30929 18411 30987 18417
rect 30929 18377 30941 18411
rect 30975 18377 30987 18411
rect 30929 18371 30987 18377
rect 26082 18312 26280 18340
rect 26510 18300 26516 18352
rect 26568 18340 26574 18352
rect 29362 18340 29368 18352
rect 26568 18312 29368 18340
rect 26568 18300 26574 18312
rect 22073 18275 22131 18281
rect 22073 18241 22085 18275
rect 22119 18272 22131 18275
rect 22189 18275 22247 18281
rect 22119 18241 22140 18272
rect 22073 18235 22140 18241
rect 22189 18241 22201 18275
rect 22235 18241 22247 18275
rect 22189 18235 22247 18241
rect 22281 18275 22339 18281
rect 22281 18241 22293 18275
rect 22327 18272 22339 18275
rect 22370 18272 22376 18284
rect 22327 18244 22376 18272
rect 22327 18241 22339 18244
rect 22281 18235 22339 18241
rect 20622 18204 20628 18216
rect 20180 18176 20628 18204
rect 20073 18167 20131 18173
rect 20622 18164 20628 18176
rect 20680 18164 20686 18216
rect 22112 18204 22140 18235
rect 22370 18232 22376 18244
rect 22428 18232 22434 18284
rect 22462 18232 22468 18284
rect 22520 18232 22526 18284
rect 23385 18275 23443 18281
rect 23385 18241 23397 18275
rect 23431 18241 23443 18275
rect 23385 18235 23443 18241
rect 23477 18275 23535 18281
rect 23477 18241 23489 18275
rect 23523 18241 23535 18275
rect 23477 18235 23535 18241
rect 23290 18204 23296 18216
rect 22112 18176 23296 18204
rect 23290 18164 23296 18176
rect 23348 18204 23354 18216
rect 23400 18204 23428 18235
rect 23348 18176 23428 18204
rect 23492 18204 23520 18235
rect 23566 18232 23572 18284
rect 23624 18232 23630 18284
rect 23753 18275 23811 18281
rect 23753 18241 23765 18275
rect 23799 18272 23811 18275
rect 23842 18272 23848 18284
rect 23799 18244 23848 18272
rect 23799 18241 23811 18244
rect 23753 18235 23811 18241
rect 23842 18232 23848 18244
rect 23900 18272 23906 18284
rect 25130 18272 25136 18284
rect 23900 18244 25136 18272
rect 23900 18232 23906 18244
rect 25130 18232 25136 18244
rect 25188 18232 25194 18284
rect 27982 18232 27988 18284
rect 28040 18232 28046 18284
rect 28166 18232 28172 18284
rect 28224 18232 28230 18284
rect 28258 18232 28264 18284
rect 28316 18232 28322 18284
rect 28552 18281 28580 18312
rect 29362 18300 29368 18312
rect 29420 18340 29426 18352
rect 29420 18312 30420 18340
rect 29420 18300 29426 18312
rect 28537 18275 28595 18281
rect 28537 18241 28549 18275
rect 28583 18241 28595 18275
rect 28537 18235 28595 18241
rect 28813 18275 28871 18281
rect 28813 18241 28825 18275
rect 28859 18272 28871 18275
rect 30190 18272 30196 18284
rect 28859 18244 30196 18272
rect 28859 18241 28871 18244
rect 28813 18235 28871 18241
rect 30190 18232 30196 18244
rect 30248 18232 30254 18284
rect 30392 18281 30420 18312
rect 30285 18275 30343 18281
rect 30285 18241 30297 18275
rect 30331 18241 30343 18275
rect 30285 18235 30343 18241
rect 30378 18275 30436 18281
rect 30378 18241 30390 18275
rect 30424 18241 30436 18275
rect 30378 18235 30436 18241
rect 25038 18204 25044 18216
rect 23492 18176 25044 18204
rect 23348 18164 23354 18176
rect 25038 18164 25044 18176
rect 25096 18164 25102 18216
rect 26510 18164 26516 18216
rect 26568 18164 26574 18216
rect 26789 18207 26847 18213
rect 26789 18173 26801 18207
rect 26835 18204 26847 18207
rect 26970 18204 26976 18216
rect 26835 18176 26976 18204
rect 26835 18173 26847 18176
rect 26789 18167 26847 18173
rect 26970 18164 26976 18176
rect 27028 18164 27034 18216
rect 28184 18204 28212 18232
rect 28629 18207 28687 18213
rect 28629 18204 28641 18207
rect 28184 18176 28641 18204
rect 28629 18173 28641 18176
rect 28675 18204 28687 18207
rect 28997 18207 29055 18213
rect 28997 18204 29009 18207
rect 28675 18176 29009 18204
rect 28675 18173 28687 18176
rect 28629 18167 28687 18173
rect 28997 18173 29009 18176
rect 29043 18204 29055 18207
rect 29181 18207 29239 18213
rect 29181 18204 29193 18207
rect 29043 18176 29193 18204
rect 29043 18173 29055 18176
rect 28997 18167 29055 18173
rect 29181 18173 29193 18176
rect 29227 18173 29239 18207
rect 29181 18167 29239 18173
rect 30098 18164 30104 18216
rect 30156 18204 30162 18216
rect 30300 18204 30328 18235
rect 30558 18232 30564 18284
rect 30616 18232 30622 18284
rect 30653 18275 30711 18281
rect 30653 18241 30665 18275
rect 30699 18241 30711 18275
rect 30653 18235 30711 18241
rect 30156 18176 30328 18204
rect 30156 18164 30162 18176
rect 16666 18096 16672 18148
rect 16724 18096 16730 18148
rect 20441 18139 20499 18145
rect 20441 18105 20453 18139
rect 20487 18136 20499 18139
rect 22094 18136 22100 18148
rect 20487 18108 22100 18136
rect 20487 18105 20499 18108
rect 20441 18099 20499 18105
rect 22094 18096 22100 18108
rect 22152 18096 22158 18148
rect 24578 18096 24584 18148
rect 24636 18136 24642 18148
rect 24673 18139 24731 18145
rect 24673 18136 24685 18139
rect 24636 18108 24685 18136
rect 24636 18096 24642 18108
rect 24673 18105 24685 18108
rect 24719 18105 24731 18139
rect 24673 18099 24731 18105
rect 28445 18139 28503 18145
rect 28445 18105 28457 18139
rect 28491 18136 28503 18139
rect 29454 18136 29460 18148
rect 28491 18108 29460 18136
rect 28491 18105 28503 18108
rect 28445 18099 28503 18105
rect 29454 18096 29460 18108
rect 29512 18096 29518 18148
rect 22370 18028 22376 18080
rect 22428 18068 22434 18080
rect 23566 18068 23572 18080
rect 22428 18040 23572 18068
rect 22428 18028 22434 18040
rect 23566 18028 23572 18040
rect 23624 18028 23630 18080
rect 26050 18028 26056 18080
rect 26108 18068 26114 18080
rect 26973 18071 27031 18077
rect 26973 18068 26985 18071
rect 26108 18040 26985 18068
rect 26108 18028 26114 18040
rect 26973 18037 26985 18040
rect 27019 18037 27031 18071
rect 30300 18068 30328 18176
rect 30668 18136 30696 18235
rect 30742 18232 30748 18284
rect 30800 18281 30806 18284
rect 30800 18272 30808 18281
rect 30944 18272 30972 18371
rect 32122 18368 32128 18420
rect 32180 18368 32186 18420
rect 37090 18368 37096 18420
rect 37148 18368 37154 18420
rect 37734 18368 37740 18420
rect 37792 18368 37798 18420
rect 38010 18368 38016 18420
rect 38068 18368 38074 18420
rect 38289 18411 38347 18417
rect 38289 18377 38301 18411
rect 38335 18408 38347 18411
rect 40034 18408 40040 18420
rect 38335 18380 40040 18408
rect 38335 18377 38347 18380
rect 38289 18371 38347 18377
rect 40034 18368 40040 18380
rect 40092 18368 40098 18420
rect 40126 18368 40132 18420
rect 40184 18408 40190 18420
rect 40405 18411 40463 18417
rect 40405 18408 40417 18411
rect 40184 18380 40417 18408
rect 40184 18368 40190 18380
rect 40405 18377 40417 18380
rect 40451 18377 40463 18411
rect 40954 18408 40960 18420
rect 40405 18371 40463 18377
rect 40788 18380 40960 18408
rect 37366 18340 37372 18352
rect 36846 18312 37372 18340
rect 37366 18300 37372 18312
rect 37424 18300 37430 18352
rect 37752 18340 37780 18368
rect 37921 18343 37979 18349
rect 37921 18340 37933 18343
rect 37752 18312 37933 18340
rect 37921 18309 37933 18312
rect 37967 18309 37979 18343
rect 38028 18340 38056 18368
rect 38028 18312 38148 18340
rect 37921 18303 37979 18309
rect 32309 18275 32367 18281
rect 32309 18272 32321 18275
rect 30800 18244 30845 18272
rect 30944 18244 32321 18272
rect 30800 18235 30808 18244
rect 32309 18241 32321 18244
rect 32355 18241 32367 18275
rect 32309 18235 32367 18241
rect 30800 18232 30806 18235
rect 32490 18232 32496 18284
rect 32548 18272 32554 18284
rect 34054 18272 34060 18284
rect 32548 18244 34060 18272
rect 32548 18232 32554 18244
rect 34054 18232 34060 18244
rect 34112 18232 34118 18284
rect 37734 18232 37740 18284
rect 37792 18232 37798 18284
rect 31110 18164 31116 18216
rect 31168 18164 31174 18216
rect 31665 18207 31723 18213
rect 31665 18173 31677 18207
rect 31711 18204 31723 18207
rect 32585 18207 32643 18213
rect 32585 18204 32597 18207
rect 31711 18176 32597 18204
rect 31711 18173 31723 18176
rect 31665 18167 31723 18173
rect 32585 18173 32597 18176
rect 32631 18173 32643 18207
rect 32585 18167 32643 18173
rect 33502 18164 33508 18216
rect 33560 18204 33566 18216
rect 35345 18207 35403 18213
rect 35345 18204 35357 18207
rect 33560 18176 35357 18204
rect 33560 18164 33566 18176
rect 35345 18173 35357 18176
rect 35391 18173 35403 18207
rect 35345 18167 35403 18173
rect 35621 18207 35679 18213
rect 35621 18173 35633 18207
rect 35667 18204 35679 18207
rect 35986 18204 35992 18216
rect 35667 18176 35992 18204
rect 35667 18173 35679 18176
rect 35621 18167 35679 18173
rect 35986 18164 35992 18176
rect 36044 18164 36050 18216
rect 31478 18136 31484 18148
rect 30668 18108 31484 18136
rect 31478 18096 31484 18108
rect 31536 18136 31542 18148
rect 32306 18136 32312 18148
rect 31536 18108 32312 18136
rect 31536 18096 31542 18108
rect 32306 18096 32312 18108
rect 32364 18096 32370 18148
rect 37936 18136 37964 18303
rect 38120 18281 38148 18312
rect 38194 18300 38200 18352
rect 38252 18340 38258 18352
rect 39025 18343 39083 18349
rect 39025 18340 39037 18343
rect 38252 18312 39037 18340
rect 38252 18300 38258 18312
rect 39025 18309 39037 18312
rect 39071 18309 39083 18343
rect 39025 18303 39083 18309
rect 39945 18343 40003 18349
rect 39945 18309 39957 18343
rect 39991 18340 40003 18343
rect 40144 18340 40172 18368
rect 40788 18349 40816 18380
rect 40954 18368 40960 18380
rect 41012 18368 41018 18420
rect 41141 18411 41199 18417
rect 41141 18377 41153 18411
rect 41187 18377 41199 18411
rect 41141 18371 41199 18377
rect 42981 18411 43039 18417
rect 42981 18377 42993 18411
rect 43027 18408 43039 18411
rect 43346 18408 43352 18420
rect 43027 18380 43352 18408
rect 43027 18377 43039 18380
rect 42981 18371 43039 18377
rect 39991 18312 40172 18340
rect 40773 18343 40831 18349
rect 39991 18309 40003 18312
rect 39945 18303 40003 18309
rect 40773 18309 40785 18343
rect 40819 18309 40831 18343
rect 41156 18340 41184 18371
rect 43346 18368 43352 18380
rect 43404 18368 43410 18420
rect 45462 18368 45468 18420
rect 45520 18408 45526 18420
rect 45557 18411 45615 18417
rect 45557 18408 45569 18411
rect 45520 18380 45569 18408
rect 45520 18368 45526 18380
rect 45557 18377 45569 18380
rect 45603 18377 45615 18411
rect 45557 18371 45615 18377
rect 56689 18411 56747 18417
rect 56689 18377 56701 18411
rect 56735 18408 56747 18411
rect 56962 18408 56968 18420
rect 56735 18380 56968 18408
rect 56735 18377 56747 18380
rect 56689 18371 56747 18377
rect 56962 18368 56968 18380
rect 57020 18368 57026 18420
rect 50157 18343 50215 18349
rect 41156 18312 41552 18340
rect 40773 18303 40831 18309
rect 38013 18275 38071 18281
rect 38013 18241 38025 18275
rect 38059 18241 38071 18275
rect 38013 18235 38071 18241
rect 38105 18275 38163 18281
rect 38105 18241 38117 18275
rect 38151 18241 38163 18275
rect 38381 18275 38439 18281
rect 38381 18272 38393 18275
rect 38105 18235 38163 18241
rect 38304 18244 38393 18272
rect 38028 18204 38056 18235
rect 38304 18204 38332 18244
rect 38381 18241 38393 18244
rect 38427 18241 38439 18275
rect 38381 18235 38439 18241
rect 38562 18232 38568 18284
rect 38620 18232 38626 18284
rect 38654 18232 38660 18284
rect 38712 18232 38718 18284
rect 38749 18275 38807 18281
rect 38749 18241 38761 18275
rect 38795 18272 38807 18275
rect 38930 18272 38936 18284
rect 38795 18244 38936 18272
rect 38795 18241 38807 18244
rect 38749 18235 38807 18241
rect 38930 18232 38936 18244
rect 38988 18232 38994 18284
rect 39206 18232 39212 18284
rect 39264 18232 39270 18284
rect 39301 18275 39359 18281
rect 39301 18241 39313 18275
rect 39347 18241 39359 18275
rect 39301 18235 39359 18241
rect 38838 18204 38844 18216
rect 38028 18176 38844 18204
rect 38838 18164 38844 18176
rect 38896 18164 38902 18216
rect 39316 18204 39344 18235
rect 39574 18232 39580 18284
rect 39632 18232 39638 18284
rect 39666 18232 39672 18284
rect 39724 18232 39730 18284
rect 39758 18232 39764 18284
rect 39816 18272 39822 18284
rect 40037 18275 40095 18281
rect 39816 18244 39861 18272
rect 39816 18232 39822 18244
rect 40037 18241 40049 18275
rect 40083 18241 40095 18275
rect 40037 18235 40095 18241
rect 38948 18176 39344 18204
rect 38654 18136 38660 18148
rect 37936 18108 38660 18136
rect 38654 18096 38660 18108
rect 38712 18096 38718 18148
rect 38948 18145 38976 18176
rect 39482 18164 39488 18216
rect 39540 18164 39546 18216
rect 40052 18204 40080 18235
rect 40126 18232 40132 18284
rect 40184 18281 40190 18284
rect 40184 18272 40192 18281
rect 40310 18272 40316 18284
rect 40184 18244 40316 18272
rect 40184 18235 40192 18244
rect 40184 18232 40190 18235
rect 40310 18232 40316 18244
rect 40368 18232 40374 18284
rect 40494 18232 40500 18284
rect 40552 18272 40558 18284
rect 40589 18275 40647 18281
rect 40589 18272 40601 18275
rect 40552 18244 40601 18272
rect 40552 18232 40558 18244
rect 40589 18241 40601 18244
rect 40635 18241 40647 18275
rect 40589 18235 40647 18241
rect 40862 18232 40868 18284
rect 40920 18232 40926 18284
rect 40954 18232 40960 18284
rect 41012 18232 41018 18284
rect 41524 18281 41552 18312
rect 50157 18309 50169 18343
rect 50203 18340 50215 18343
rect 50522 18340 50528 18352
rect 50203 18312 50528 18340
rect 50203 18309 50215 18312
rect 50157 18303 50215 18309
rect 50522 18300 50528 18312
rect 50580 18340 50586 18352
rect 51258 18340 51264 18352
rect 50580 18312 51264 18340
rect 50580 18300 50586 18312
rect 51258 18300 51264 18312
rect 51316 18300 51322 18352
rect 56980 18340 57008 18368
rect 56980 18312 57100 18340
rect 41233 18275 41291 18281
rect 41233 18272 41245 18275
rect 41064 18244 41245 18272
rect 40218 18204 40224 18216
rect 40052 18176 40224 18204
rect 40218 18164 40224 18176
rect 40276 18164 40282 18216
rect 41064 18204 41092 18244
rect 41233 18241 41245 18244
rect 41279 18241 41291 18275
rect 41233 18235 41291 18241
rect 41509 18275 41567 18281
rect 41509 18241 41521 18275
rect 41555 18241 41567 18275
rect 41509 18235 41567 18241
rect 40880 18176 41092 18204
rect 41248 18204 41276 18235
rect 41598 18232 41604 18284
rect 41656 18232 41662 18284
rect 46201 18275 46259 18281
rect 46201 18241 46213 18275
rect 46247 18272 46259 18275
rect 46750 18272 46756 18284
rect 46247 18244 46756 18272
rect 46247 18241 46259 18244
rect 46201 18235 46259 18241
rect 46750 18232 46756 18244
rect 46808 18232 46814 18284
rect 49970 18232 49976 18284
rect 50028 18232 50034 18284
rect 50246 18232 50252 18284
rect 50304 18232 50310 18284
rect 50341 18275 50399 18281
rect 50341 18241 50353 18275
rect 50387 18272 50399 18275
rect 50430 18272 50436 18284
rect 50387 18244 50436 18272
rect 50387 18241 50399 18244
rect 50341 18235 50399 18241
rect 42978 18204 42984 18216
rect 41248 18176 42984 18204
rect 38933 18139 38991 18145
rect 38933 18105 38945 18139
rect 38979 18105 38991 18139
rect 38933 18099 38991 18105
rect 40313 18139 40371 18145
rect 40313 18105 40325 18139
rect 40359 18136 40371 18139
rect 40678 18136 40684 18148
rect 40359 18108 40684 18136
rect 40359 18105 40371 18108
rect 40313 18099 40371 18105
rect 40678 18096 40684 18108
rect 40736 18096 40742 18148
rect 31110 18068 31116 18080
rect 30300 18040 31116 18068
rect 26973 18031 27031 18037
rect 31110 18028 31116 18040
rect 31168 18068 31174 18080
rect 31757 18071 31815 18077
rect 31757 18068 31769 18071
rect 31168 18040 31769 18068
rect 31168 18028 31174 18040
rect 31757 18037 31769 18040
rect 31803 18068 31815 18071
rect 32490 18068 32496 18080
rect 31803 18040 32496 18068
rect 31803 18037 31815 18040
rect 31757 18031 31815 18037
rect 32490 18028 32496 18040
rect 32548 18028 32554 18080
rect 37366 18028 37372 18080
rect 37424 18068 37430 18080
rect 38286 18068 38292 18080
rect 37424 18040 38292 18068
rect 37424 18028 37430 18040
rect 38286 18028 38292 18040
rect 38344 18028 38350 18080
rect 38746 18028 38752 18080
rect 38804 18068 38810 18080
rect 40880 18068 40908 18176
rect 42978 18164 42984 18176
rect 43036 18164 43042 18216
rect 49050 18164 49056 18216
rect 49108 18204 49114 18216
rect 50356 18204 50384 18235
rect 50430 18232 50436 18244
rect 50488 18272 50494 18284
rect 50614 18272 50620 18284
rect 50488 18244 50620 18272
rect 50488 18232 50494 18244
rect 50614 18232 50620 18244
rect 50672 18232 50678 18284
rect 52917 18275 52975 18281
rect 52917 18241 52929 18275
rect 52963 18241 52975 18275
rect 52917 18235 52975 18241
rect 49108 18176 50384 18204
rect 49108 18164 49114 18176
rect 38804 18040 40908 18068
rect 38804 18028 38810 18040
rect 40954 18028 40960 18080
rect 41012 18068 41018 18080
rect 41322 18068 41328 18080
rect 41012 18040 41328 18068
rect 41012 18028 41018 18040
rect 41322 18028 41328 18040
rect 41380 18028 41386 18080
rect 41506 18028 41512 18080
rect 41564 18068 41570 18080
rect 41785 18071 41843 18077
rect 41785 18068 41797 18071
rect 41564 18040 41797 18068
rect 41564 18028 41570 18040
rect 41785 18037 41797 18040
rect 41831 18037 41843 18071
rect 41785 18031 41843 18037
rect 50525 18071 50583 18077
rect 50525 18037 50537 18071
rect 50571 18068 50583 18071
rect 50890 18068 50896 18080
rect 50571 18040 50896 18068
rect 50571 18037 50583 18040
rect 50525 18031 50583 18037
rect 50890 18028 50896 18040
rect 50948 18028 50954 18080
rect 52730 18028 52736 18080
rect 52788 18028 52794 18080
rect 52822 18028 52828 18080
rect 52880 18068 52886 18080
rect 52932 18068 52960 18235
rect 53006 18232 53012 18284
rect 53064 18232 53070 18284
rect 53285 18275 53343 18281
rect 53285 18241 53297 18275
rect 53331 18272 53343 18275
rect 53745 18275 53803 18281
rect 53745 18272 53757 18275
rect 53331 18244 53757 18272
rect 53331 18241 53343 18244
rect 53285 18235 53343 18241
rect 53745 18241 53757 18244
rect 53791 18241 53803 18275
rect 53745 18235 53803 18241
rect 56778 18232 56784 18284
rect 56836 18232 56842 18284
rect 56962 18232 56968 18284
rect 57020 18232 57026 18284
rect 57072 18281 57100 18312
rect 57057 18275 57115 18281
rect 57057 18241 57069 18275
rect 57103 18241 57115 18275
rect 57057 18235 57115 18241
rect 57149 18275 57207 18281
rect 57149 18241 57161 18275
rect 57195 18272 57207 18275
rect 57885 18275 57943 18281
rect 57885 18272 57897 18275
rect 57195 18244 57897 18272
rect 57195 18241 57207 18244
rect 57149 18235 57207 18241
rect 57885 18241 57897 18244
rect 57931 18241 57943 18275
rect 57885 18235 57943 18241
rect 58158 18232 58164 18284
rect 58216 18272 58222 18284
rect 58437 18275 58495 18281
rect 58437 18272 58449 18275
rect 58216 18244 58449 18272
rect 58216 18232 58222 18244
rect 58437 18241 58449 18244
rect 58483 18241 58495 18275
rect 58437 18235 58495 18241
rect 54202 18164 54208 18216
rect 54260 18204 54266 18216
rect 54297 18207 54355 18213
rect 54297 18204 54309 18207
rect 54260 18176 54309 18204
rect 54260 18164 54266 18176
rect 54297 18173 54309 18176
rect 54343 18173 54355 18207
rect 54297 18167 54355 18173
rect 53193 18139 53251 18145
rect 53193 18105 53205 18139
rect 53239 18136 53251 18139
rect 53834 18136 53840 18148
rect 53239 18108 53840 18136
rect 53239 18105 53251 18108
rect 53193 18099 53251 18105
rect 53834 18096 53840 18108
rect 53892 18136 53898 18148
rect 54754 18136 54760 18148
rect 53892 18108 54760 18136
rect 53892 18096 53898 18108
rect 54754 18096 54760 18108
rect 54812 18096 54818 18148
rect 53377 18071 53435 18077
rect 53377 18068 53389 18071
rect 52880 18040 53389 18068
rect 52880 18028 52886 18040
rect 53377 18037 53389 18040
rect 53423 18068 53435 18071
rect 54478 18068 54484 18080
rect 53423 18040 54484 18068
rect 53423 18037 53435 18040
rect 53377 18031 53435 18037
rect 54478 18028 54484 18040
rect 54536 18068 54542 18080
rect 56042 18068 56048 18080
rect 54536 18040 56048 18068
rect 54536 18028 54542 18040
rect 56042 18028 56048 18040
rect 56100 18068 56106 18080
rect 56410 18068 56416 18080
rect 56100 18040 56416 18068
rect 56100 18028 56106 18040
rect 56410 18028 56416 18040
rect 56468 18028 56474 18080
rect 57422 18028 57428 18080
rect 57480 18028 57486 18080
rect 1104 17978 58880 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 58880 17978
rect 1104 17904 58880 17926
rect 22094 17824 22100 17876
rect 22152 17864 22158 17876
rect 23106 17864 23112 17876
rect 22152 17836 23112 17864
rect 22152 17824 22158 17836
rect 23106 17824 23112 17836
rect 23164 17824 23170 17876
rect 24578 17824 24584 17876
rect 24636 17864 24642 17876
rect 24673 17867 24731 17873
rect 24673 17864 24685 17867
rect 24636 17836 24685 17864
rect 24636 17824 24642 17836
rect 24673 17833 24685 17836
rect 24719 17833 24731 17867
rect 24673 17827 24731 17833
rect 25774 17824 25780 17876
rect 25832 17824 25838 17876
rect 25961 17867 26019 17873
rect 25961 17833 25973 17867
rect 26007 17864 26019 17867
rect 26510 17864 26516 17876
rect 26007 17836 26516 17864
rect 26007 17833 26019 17836
rect 25961 17827 26019 17833
rect 26510 17824 26516 17836
rect 26568 17824 26574 17876
rect 34698 17824 34704 17876
rect 34756 17864 34762 17876
rect 35161 17867 35219 17873
rect 35161 17864 35173 17867
rect 34756 17836 35173 17864
rect 34756 17824 34762 17836
rect 35161 17833 35173 17836
rect 35207 17833 35219 17867
rect 35161 17827 35219 17833
rect 25792 17796 25820 17824
rect 26142 17796 26148 17808
rect 25792 17768 26148 17796
rect 26142 17756 26148 17768
rect 26200 17756 26206 17808
rect 35176 17796 35204 17827
rect 35986 17824 35992 17876
rect 36044 17824 36050 17876
rect 38010 17824 38016 17876
rect 38068 17864 38074 17876
rect 38381 17867 38439 17873
rect 38381 17864 38393 17867
rect 38068 17836 38393 17864
rect 38068 17824 38074 17836
rect 38381 17833 38393 17836
rect 38427 17864 38439 17867
rect 38470 17864 38476 17876
rect 38427 17836 38476 17864
rect 38427 17833 38439 17836
rect 38381 17827 38439 17833
rect 38470 17824 38476 17836
rect 38528 17824 38534 17876
rect 38654 17824 38660 17876
rect 38712 17824 38718 17876
rect 39942 17824 39948 17876
rect 40000 17824 40006 17876
rect 40678 17824 40684 17876
rect 40736 17824 40742 17876
rect 43717 17867 43775 17873
rect 43717 17864 43729 17867
rect 40972 17836 43729 17864
rect 36170 17796 36176 17808
rect 35176 17768 36176 17796
rect 36170 17756 36176 17768
rect 36228 17796 36234 17808
rect 36449 17799 36507 17805
rect 36449 17796 36461 17799
rect 36228 17768 36461 17796
rect 36228 17756 36234 17768
rect 36449 17765 36461 17768
rect 36495 17765 36507 17799
rect 36449 17759 36507 17765
rect 36633 17799 36691 17805
rect 36633 17765 36645 17799
rect 36679 17765 36691 17799
rect 37090 17796 37096 17808
rect 36633 17759 36691 17765
rect 36740 17768 37096 17796
rect 26602 17728 26608 17740
rect 26160 17700 26608 17728
rect 16666 17620 16672 17672
rect 16724 17620 16730 17672
rect 26160 17669 26188 17700
rect 26602 17688 26608 17700
rect 26660 17688 26666 17740
rect 30374 17688 30380 17740
rect 30432 17728 30438 17740
rect 30745 17731 30803 17737
rect 30745 17728 30757 17731
rect 30432 17700 30757 17728
rect 30432 17688 30438 17700
rect 30745 17697 30757 17700
rect 30791 17728 30803 17731
rect 31570 17728 31576 17740
rect 30791 17700 31576 17728
rect 30791 17697 30803 17700
rect 30745 17691 30803 17697
rect 31570 17688 31576 17700
rect 31628 17688 31634 17740
rect 36648 17728 36676 17759
rect 36464 17700 36676 17728
rect 26145 17663 26203 17669
rect 26145 17629 26157 17663
rect 26191 17629 26203 17663
rect 26145 17623 26203 17629
rect 26326 17620 26332 17672
rect 26384 17620 26390 17672
rect 26418 17620 26424 17672
rect 26476 17620 26482 17672
rect 30282 17620 30288 17672
rect 30340 17620 30346 17672
rect 34514 17620 34520 17672
rect 34572 17660 34578 17672
rect 34882 17660 34888 17672
rect 34572 17632 34888 17660
rect 34572 17620 34578 17632
rect 34882 17620 34888 17632
rect 34940 17620 34946 17672
rect 34977 17663 35035 17669
rect 34977 17629 34989 17663
rect 35023 17660 35035 17663
rect 35066 17660 35072 17672
rect 35023 17632 35072 17660
rect 35023 17629 35035 17632
rect 34977 17623 35035 17629
rect 35066 17620 35072 17632
rect 35124 17620 35130 17672
rect 35250 17669 35256 17672
rect 35235 17663 35256 17669
rect 35235 17629 35247 17663
rect 35235 17623 35256 17629
rect 35250 17620 35256 17623
rect 35308 17620 35314 17672
rect 36170 17620 36176 17672
rect 36228 17620 36234 17672
rect 36265 17663 36323 17669
rect 36265 17629 36277 17663
rect 36311 17660 36323 17663
rect 36464 17660 36492 17700
rect 36311 17632 36492 17660
rect 36311 17629 36323 17632
rect 36265 17623 36323 17629
rect 36538 17620 36544 17672
rect 36596 17660 36602 17672
rect 36740 17660 36768 17768
rect 37090 17756 37096 17768
rect 37148 17756 37154 17808
rect 38102 17756 38108 17808
rect 38160 17796 38166 17808
rect 39206 17796 39212 17808
rect 38160 17768 39212 17796
rect 38160 17756 38166 17768
rect 39206 17756 39212 17768
rect 39264 17756 39270 17808
rect 37734 17728 37740 17740
rect 36924 17700 37740 17728
rect 36596 17632 36768 17660
rect 36596 17620 36602 17632
rect 36814 17620 36820 17672
rect 36872 17620 36878 17672
rect 36924 17669 36952 17700
rect 37734 17688 37740 17700
rect 37792 17688 37798 17740
rect 40034 17688 40040 17740
rect 40092 17688 40098 17740
rect 36909 17663 36967 17669
rect 36909 17629 36921 17663
rect 36955 17629 36967 17663
rect 36909 17623 36967 17629
rect 37185 17663 37243 17669
rect 37185 17629 37197 17663
rect 37231 17660 37243 17663
rect 38746 17660 38752 17672
rect 37231 17632 38752 17660
rect 37231 17629 37243 17632
rect 37185 17623 37243 17629
rect 25038 17552 25044 17604
rect 25096 17592 25102 17604
rect 26436 17592 26464 17620
rect 25096 17564 26464 17592
rect 25096 17552 25102 17564
rect 31018 17552 31024 17604
rect 31076 17552 31082 17604
rect 31478 17552 31484 17604
rect 31536 17552 31542 17604
rect 35986 17592 35992 17604
rect 35360 17564 35992 17592
rect 30466 17484 30472 17536
rect 30524 17524 30530 17536
rect 30742 17524 30748 17536
rect 30524 17496 30748 17524
rect 30524 17484 30530 17496
rect 30742 17484 30748 17496
rect 30800 17524 30806 17536
rect 31662 17524 31668 17536
rect 30800 17496 31668 17524
rect 30800 17484 30806 17496
rect 31662 17484 31668 17496
rect 31720 17484 31726 17536
rect 32306 17484 32312 17536
rect 32364 17524 32370 17536
rect 32493 17527 32551 17533
rect 32493 17524 32505 17527
rect 32364 17496 32505 17524
rect 32364 17484 32370 17496
rect 32493 17493 32505 17496
rect 32539 17493 32551 17527
rect 32493 17487 32551 17493
rect 33778 17484 33784 17536
rect 33836 17524 33842 17536
rect 34701 17527 34759 17533
rect 34701 17524 34713 17527
rect 33836 17496 34713 17524
rect 33836 17484 33842 17496
rect 34701 17493 34713 17496
rect 34747 17493 34759 17527
rect 34701 17487 34759 17493
rect 35250 17484 35256 17536
rect 35308 17524 35314 17536
rect 35360 17524 35388 17564
rect 35986 17552 35992 17564
rect 36044 17592 36050 17604
rect 36924 17592 36952 17623
rect 38746 17620 38752 17632
rect 38804 17620 38810 17672
rect 40129 17663 40187 17669
rect 40129 17660 40141 17663
rect 38856 17632 40141 17660
rect 36044 17564 36952 17592
rect 36044 17552 36050 17564
rect 36998 17552 37004 17604
rect 37056 17552 37062 17604
rect 37090 17552 37096 17604
rect 37148 17592 37154 17604
rect 37550 17592 37556 17604
rect 37148 17564 37556 17592
rect 37148 17552 37154 17564
rect 37550 17552 37556 17564
rect 37608 17592 37614 17604
rect 38856 17592 38884 17632
rect 40129 17629 40141 17632
rect 40175 17660 40187 17663
rect 40405 17663 40463 17669
rect 40405 17660 40417 17663
rect 40175 17632 40417 17660
rect 40175 17629 40187 17632
rect 40129 17623 40187 17629
rect 40405 17629 40417 17632
rect 40451 17629 40463 17663
rect 40405 17623 40463 17629
rect 40586 17620 40592 17672
rect 40644 17660 40650 17672
rect 40972 17669 41000 17836
rect 43717 17833 43729 17836
rect 43763 17833 43775 17867
rect 43717 17827 43775 17833
rect 43806 17824 43812 17876
rect 43864 17824 43870 17876
rect 47486 17864 47492 17876
rect 46584 17836 47492 17864
rect 42610 17756 42616 17808
rect 42668 17796 42674 17808
rect 46584 17796 46612 17836
rect 47486 17824 47492 17836
rect 47544 17824 47550 17876
rect 48590 17824 48596 17876
rect 48648 17864 48654 17876
rect 49053 17867 49111 17873
rect 49053 17864 49065 17867
rect 48648 17836 49065 17864
rect 48648 17824 48654 17836
rect 49053 17833 49065 17836
rect 49099 17864 49111 17867
rect 49326 17864 49332 17876
rect 49099 17836 49332 17864
rect 49099 17833 49111 17836
rect 49053 17827 49111 17833
rect 49326 17824 49332 17836
rect 49384 17824 49390 17876
rect 49510 17824 49516 17876
rect 49568 17824 49574 17876
rect 49881 17867 49939 17873
rect 49881 17833 49893 17867
rect 49927 17864 49939 17867
rect 56594 17864 56600 17876
rect 49927 17836 56600 17864
rect 49927 17833 49939 17836
rect 49881 17827 49939 17833
rect 56594 17824 56600 17836
rect 56652 17824 56658 17876
rect 58158 17824 58164 17876
rect 58216 17864 58222 17876
rect 58253 17867 58311 17873
rect 58253 17864 58265 17867
rect 58216 17836 58265 17864
rect 58216 17824 58222 17836
rect 58253 17833 58265 17836
rect 58299 17833 58311 17867
rect 58253 17827 58311 17833
rect 42668 17768 46612 17796
rect 42668 17756 42674 17768
rect 47946 17756 47952 17808
rect 48004 17796 48010 17808
rect 49694 17796 49700 17808
rect 48004 17768 49700 17796
rect 48004 17756 48010 17768
rect 49694 17756 49700 17768
rect 49752 17796 49758 17808
rect 49752 17768 50660 17796
rect 49752 17756 49758 17768
rect 41506 17688 41512 17740
rect 41564 17688 41570 17740
rect 42978 17688 42984 17740
rect 43036 17728 43042 17740
rect 43036 17700 43209 17728
rect 43036 17688 43042 17700
rect 40865 17663 40923 17669
rect 40865 17660 40877 17663
rect 40644 17632 40877 17660
rect 40644 17620 40650 17632
rect 40865 17629 40877 17632
rect 40911 17629 40923 17663
rect 40865 17623 40923 17629
rect 40957 17663 41015 17669
rect 40957 17629 40969 17663
rect 41003 17629 41015 17663
rect 40957 17623 41015 17629
rect 41230 17620 41236 17672
rect 41288 17620 41294 17672
rect 43070 17620 43076 17672
rect 43128 17620 43134 17672
rect 43181 17669 43209 17700
rect 45002 17688 45008 17740
rect 45060 17728 45066 17740
rect 46477 17731 46535 17737
rect 46477 17728 46489 17731
rect 45060 17700 46489 17728
rect 45060 17688 45066 17700
rect 46477 17697 46489 17700
rect 46523 17697 46535 17731
rect 46477 17691 46535 17697
rect 48225 17731 48283 17737
rect 48225 17697 48237 17731
rect 48271 17728 48283 17731
rect 48271 17700 48912 17728
rect 48271 17697 48283 17700
rect 48225 17691 48283 17697
rect 43166 17663 43224 17669
rect 43166 17629 43178 17663
rect 43212 17629 43224 17663
rect 43166 17623 43224 17629
rect 43346 17620 43352 17672
rect 43404 17620 43410 17672
rect 43438 17620 43444 17672
rect 43496 17620 43502 17672
rect 43579 17663 43637 17669
rect 43579 17629 43591 17663
rect 43625 17660 43637 17663
rect 43806 17660 43812 17672
rect 43625 17632 43812 17660
rect 43625 17629 43637 17632
rect 43579 17623 43637 17629
rect 43806 17620 43812 17632
rect 43864 17620 43870 17672
rect 47854 17620 47860 17672
rect 47912 17620 47918 17672
rect 48884 17669 48912 17700
rect 48958 17688 48964 17740
rect 49016 17728 49022 17740
rect 49513 17731 49571 17737
rect 49513 17728 49525 17731
rect 49016 17700 49525 17728
rect 49016 17688 49022 17700
rect 49513 17697 49525 17700
rect 49559 17697 49571 17731
rect 49970 17728 49976 17740
rect 49513 17691 49571 17697
rect 49620 17700 49976 17728
rect 48869 17663 48927 17669
rect 48869 17629 48881 17663
rect 48915 17660 48927 17663
rect 49050 17660 49056 17672
rect 48915 17632 49056 17660
rect 48915 17629 48927 17632
rect 48869 17623 48927 17629
rect 49050 17620 49056 17632
rect 49108 17660 49114 17672
rect 49620 17660 49648 17700
rect 49970 17688 49976 17700
rect 50028 17688 50034 17740
rect 50632 17737 50660 17768
rect 54478 17756 54484 17808
rect 54536 17796 54542 17808
rect 54941 17799 54999 17805
rect 54941 17796 54953 17799
rect 54536 17768 54953 17796
rect 54536 17756 54542 17768
rect 54941 17765 54953 17768
rect 54987 17765 54999 17799
rect 54941 17759 54999 17765
rect 55950 17756 55956 17808
rect 56008 17796 56014 17808
rect 56045 17799 56103 17805
rect 56045 17796 56057 17799
rect 56008 17768 56057 17796
rect 56008 17756 56014 17768
rect 56045 17765 56057 17768
rect 56091 17765 56103 17799
rect 56045 17759 56103 17765
rect 50617 17731 50675 17737
rect 50617 17697 50629 17731
rect 50663 17697 50675 17731
rect 50617 17691 50675 17697
rect 52457 17731 52515 17737
rect 52457 17697 52469 17731
rect 52503 17728 52515 17731
rect 53926 17728 53932 17740
rect 52503 17700 53932 17728
rect 52503 17697 52515 17700
rect 52457 17691 52515 17697
rect 53926 17688 53932 17700
rect 53984 17688 53990 17740
rect 54754 17688 54760 17740
rect 54812 17688 54818 17740
rect 55214 17688 55220 17740
rect 55272 17728 55278 17740
rect 56689 17731 56747 17737
rect 56689 17728 56701 17731
rect 55272 17700 56701 17728
rect 55272 17688 55278 17700
rect 56689 17697 56701 17700
rect 56735 17697 56747 17731
rect 56689 17691 56747 17697
rect 49108 17632 49648 17660
rect 49108 17620 49114 17632
rect 49694 17620 49700 17672
rect 49752 17620 49758 17672
rect 53834 17620 53840 17672
rect 53892 17620 53898 17672
rect 54478 17620 54484 17672
rect 54536 17620 54542 17672
rect 54570 17620 54576 17672
rect 54628 17620 54634 17672
rect 54849 17663 54907 17669
rect 54849 17629 54861 17663
rect 54895 17629 54907 17663
rect 54849 17623 54907 17629
rect 55861 17663 55919 17669
rect 55861 17629 55873 17663
rect 55907 17629 55919 17663
rect 55861 17623 55919 17629
rect 37608 17564 38884 17592
rect 37608 17552 37614 17564
rect 39850 17552 39856 17604
rect 39908 17552 39914 17604
rect 40681 17595 40739 17601
rect 40681 17592 40693 17595
rect 40328 17564 40693 17592
rect 35308 17496 35388 17524
rect 35308 17484 35314 17496
rect 36446 17484 36452 17536
rect 36504 17524 36510 17536
rect 37016 17524 37044 17552
rect 36504 17496 37044 17524
rect 39577 17527 39635 17533
rect 36504 17484 36510 17496
rect 39577 17493 39589 17527
rect 39623 17524 39635 17527
rect 40126 17524 40132 17536
rect 39623 17496 40132 17524
rect 39623 17493 39635 17496
rect 39577 17487 39635 17493
rect 40126 17484 40132 17496
rect 40184 17484 40190 17536
rect 40328 17533 40356 17564
rect 40681 17561 40693 17564
rect 40727 17561 40739 17595
rect 44082 17592 44088 17604
rect 42734 17564 44088 17592
rect 40681 17555 40739 17561
rect 44082 17552 44088 17564
rect 44140 17552 44146 17604
rect 46750 17552 46756 17604
rect 46808 17552 46814 17604
rect 48406 17552 48412 17604
rect 48464 17592 48470 17604
rect 49421 17595 49479 17601
rect 49421 17592 49433 17595
rect 48464 17564 49433 17592
rect 48464 17552 48470 17564
rect 49421 17561 49433 17564
rect 49467 17561 49479 17595
rect 49421 17555 49479 17561
rect 50614 17552 50620 17604
rect 50672 17592 50678 17604
rect 50893 17595 50951 17601
rect 50893 17592 50905 17595
rect 50672 17564 50905 17592
rect 50672 17552 50678 17564
rect 50893 17561 50905 17564
rect 50939 17561 50951 17595
rect 50893 17555 50951 17561
rect 51350 17552 51356 17604
rect 51408 17552 51414 17604
rect 52730 17552 52736 17604
rect 52788 17552 52794 17604
rect 54864 17592 54892 17623
rect 55766 17592 55772 17604
rect 54036 17564 55772 17592
rect 40313 17527 40371 17533
rect 40313 17493 40325 17527
rect 40359 17493 40371 17527
rect 40313 17487 40371 17493
rect 41138 17484 41144 17536
rect 41196 17484 41202 17536
rect 41322 17484 41328 17536
rect 41380 17524 41386 17536
rect 47578 17524 47584 17536
rect 41380 17496 47584 17524
rect 41380 17484 41386 17496
rect 47578 17484 47584 17496
rect 47636 17524 47642 17536
rect 48222 17524 48228 17536
rect 47636 17496 48228 17524
rect 47636 17484 47642 17496
rect 48222 17484 48228 17496
rect 48280 17484 48286 17536
rect 48314 17484 48320 17536
rect 48372 17484 48378 17536
rect 52362 17484 52368 17536
rect 52420 17484 52426 17536
rect 53098 17484 53104 17536
rect 53156 17524 53162 17536
rect 54036 17524 54064 17564
rect 55766 17552 55772 17564
rect 55824 17552 55830 17604
rect 53156 17496 54064 17524
rect 53156 17484 53162 17496
rect 54202 17484 54208 17536
rect 54260 17484 54266 17536
rect 54297 17527 54355 17533
rect 54297 17493 54309 17527
rect 54343 17524 54355 17527
rect 54386 17524 54392 17536
rect 54343 17496 54392 17524
rect 54343 17493 54355 17496
rect 54297 17487 54355 17493
rect 54386 17484 54392 17496
rect 54444 17484 54450 17536
rect 55674 17484 55680 17536
rect 55732 17524 55738 17536
rect 55876 17524 55904 17623
rect 56410 17620 56416 17672
rect 56468 17620 56474 17672
rect 56505 17663 56563 17669
rect 56505 17629 56517 17663
rect 56551 17660 56563 17663
rect 56594 17660 56600 17672
rect 56551 17632 56600 17660
rect 56551 17629 56563 17632
rect 56505 17623 56563 17629
rect 56594 17620 56600 17632
rect 56652 17620 56658 17672
rect 56781 17663 56839 17669
rect 56781 17660 56793 17663
rect 56704 17632 56793 17660
rect 56704 17604 56732 17632
rect 56781 17629 56793 17632
rect 56827 17629 56839 17663
rect 56781 17623 56839 17629
rect 56870 17620 56876 17672
rect 56928 17620 56934 17672
rect 57140 17663 57198 17669
rect 57140 17629 57152 17663
rect 57186 17660 57198 17663
rect 57422 17660 57428 17672
rect 57186 17632 57428 17660
rect 57186 17629 57198 17632
rect 57140 17623 57198 17629
rect 57422 17620 57428 17632
rect 57480 17620 57486 17672
rect 56686 17552 56692 17604
rect 56744 17552 56750 17604
rect 55732 17496 55904 17524
rect 55732 17484 55738 17496
rect 56226 17484 56232 17536
rect 56284 17484 56290 17536
rect 1104 17434 58880 17456
rect 1104 17382 4874 17434
rect 4926 17382 4938 17434
rect 4990 17382 5002 17434
rect 5054 17382 5066 17434
rect 5118 17382 5130 17434
rect 5182 17382 35594 17434
rect 35646 17382 35658 17434
rect 35710 17382 35722 17434
rect 35774 17382 35786 17434
rect 35838 17382 35850 17434
rect 35902 17382 58880 17434
rect 1104 17360 58880 17382
rect 16758 17280 16764 17332
rect 16816 17320 16822 17332
rect 24857 17323 24915 17329
rect 24857 17320 24869 17323
rect 16816 17292 24869 17320
rect 16816 17280 16822 17292
rect 24857 17289 24869 17292
rect 24903 17289 24915 17323
rect 26513 17323 26571 17329
rect 26513 17320 26525 17323
rect 24857 17283 24915 17289
rect 26160 17292 26525 17320
rect 17954 17212 17960 17264
rect 18012 17212 18018 17264
rect 19705 17255 19763 17261
rect 19705 17221 19717 17255
rect 19751 17252 19763 17255
rect 21634 17252 21640 17264
rect 19751 17224 21640 17252
rect 19751 17221 19763 17224
rect 19705 17215 19763 17221
rect 21634 17212 21640 17224
rect 21692 17212 21698 17264
rect 22278 17212 22284 17264
rect 22336 17252 22342 17264
rect 24305 17255 24363 17261
rect 24305 17252 24317 17255
rect 22336 17224 24317 17252
rect 22336 17212 22342 17224
rect 24305 17221 24317 17224
rect 24351 17221 24363 17255
rect 24305 17215 24363 17221
rect 24670 17212 24676 17264
rect 24728 17212 24734 17264
rect 19061 17187 19119 17193
rect 19061 17153 19073 17187
rect 19107 17184 19119 17187
rect 19608 17187 19666 17193
rect 19107 17156 19472 17184
rect 19107 17153 19119 17156
rect 19061 17147 19119 17153
rect 16666 17076 16672 17128
rect 16724 17116 16730 17128
rect 17037 17119 17095 17125
rect 17037 17116 17049 17119
rect 16724 17088 17049 17116
rect 16724 17076 16730 17088
rect 17037 17085 17049 17088
rect 17083 17085 17095 17119
rect 17037 17079 17095 17085
rect 17313 17119 17371 17125
rect 17313 17085 17325 17119
rect 17359 17116 17371 17119
rect 18877 17119 18935 17125
rect 18877 17116 18889 17119
rect 17359 17088 18889 17116
rect 17359 17085 17371 17088
rect 17313 17079 17371 17085
rect 18877 17085 18889 17088
rect 18923 17085 18935 17119
rect 19334 17116 19340 17128
rect 18877 17079 18935 17085
rect 19306 17076 19340 17116
rect 19392 17076 19398 17128
rect 18785 17051 18843 17057
rect 18785 17017 18797 17051
rect 18831 17048 18843 17051
rect 19306 17048 19334 17076
rect 19444 17057 19472 17156
rect 19608 17153 19620 17187
rect 19654 17153 19666 17187
rect 19608 17147 19666 17153
rect 19623 17116 19651 17147
rect 19794 17144 19800 17196
rect 19852 17144 19858 17196
rect 19980 17187 20038 17193
rect 19980 17153 19992 17187
rect 20026 17153 20038 17187
rect 19980 17147 20038 17153
rect 20073 17187 20131 17193
rect 20073 17153 20085 17187
rect 20119 17184 20131 17187
rect 20346 17184 20352 17196
rect 20119 17156 20352 17184
rect 20119 17153 20131 17156
rect 20073 17147 20131 17153
rect 19702 17116 19708 17128
rect 19623 17088 19708 17116
rect 19702 17076 19708 17088
rect 19760 17076 19766 17128
rect 19996 17116 20024 17147
rect 20346 17144 20352 17156
rect 20404 17144 20410 17196
rect 23109 17187 23167 17193
rect 23109 17153 23121 17187
rect 23155 17184 23167 17187
rect 23198 17184 23204 17196
rect 23155 17156 23204 17184
rect 23155 17153 23167 17156
rect 23109 17147 23167 17153
rect 23198 17144 23204 17156
rect 23256 17144 23262 17196
rect 24026 17144 24032 17196
rect 24084 17144 24090 17196
rect 24213 17187 24271 17193
rect 24213 17153 24225 17187
rect 24259 17153 24271 17187
rect 24213 17147 24271 17153
rect 24397 17187 24455 17193
rect 24397 17153 24409 17187
rect 24443 17184 24455 17187
rect 24578 17184 24584 17196
rect 24443 17156 24584 17184
rect 24443 17153 24455 17156
rect 24397 17147 24455 17153
rect 20162 17116 20168 17128
rect 19996 17088 20168 17116
rect 20162 17076 20168 17088
rect 20220 17076 20226 17128
rect 23014 17076 23020 17128
rect 23072 17116 23078 17128
rect 23385 17119 23443 17125
rect 23385 17116 23397 17119
rect 23072 17088 23397 17116
rect 23072 17076 23078 17088
rect 23385 17085 23397 17088
rect 23431 17085 23443 17119
rect 24228 17116 24256 17147
rect 24578 17144 24584 17156
rect 24636 17144 24642 17196
rect 24688 17116 24716 17212
rect 24946 17144 24952 17196
rect 25004 17184 25010 17196
rect 26160 17193 26188 17292
rect 26513 17289 26525 17292
rect 26559 17320 26571 17323
rect 26786 17320 26792 17332
rect 26559 17292 26792 17320
rect 26559 17289 26571 17292
rect 26513 17283 26571 17289
rect 26786 17280 26792 17292
rect 26844 17280 26850 17332
rect 28994 17280 29000 17332
rect 29052 17320 29058 17332
rect 29181 17323 29239 17329
rect 29181 17320 29193 17323
rect 29052 17292 29193 17320
rect 29052 17280 29058 17292
rect 29181 17289 29193 17292
rect 29227 17289 29239 17323
rect 32214 17320 32220 17332
rect 29181 17283 29239 17289
rect 30760 17292 32220 17320
rect 26234 17212 26240 17264
rect 26292 17252 26298 17264
rect 30760 17261 30788 17292
rect 32214 17280 32220 17292
rect 32272 17280 32278 17332
rect 32398 17280 32404 17332
rect 32456 17280 32462 17332
rect 32490 17280 32496 17332
rect 32548 17280 32554 17332
rect 33336 17292 35112 17320
rect 26973 17255 27031 17261
rect 26973 17252 26985 17255
rect 26292 17224 26985 17252
rect 26292 17212 26298 17224
rect 26973 17221 26985 17224
rect 27019 17221 27031 17255
rect 26973 17215 27031 17221
rect 30745 17255 30803 17261
rect 30745 17221 30757 17255
rect 30791 17221 30803 17255
rect 31481 17255 31539 17261
rect 31481 17252 31493 17255
rect 30745 17215 30803 17221
rect 30944 17224 31493 17252
rect 25041 17187 25099 17193
rect 25041 17184 25053 17187
rect 25004 17156 25053 17184
rect 25004 17144 25010 17156
rect 25041 17153 25053 17156
rect 25087 17153 25099 17187
rect 25041 17147 25099 17153
rect 25317 17187 25375 17193
rect 25317 17153 25329 17187
rect 25363 17184 25375 17187
rect 25409 17187 25467 17193
rect 25409 17184 25421 17187
rect 25363 17156 25421 17184
rect 25363 17153 25375 17156
rect 25317 17147 25375 17153
rect 25409 17153 25421 17156
rect 25455 17153 25467 17187
rect 25961 17187 26019 17193
rect 25961 17184 25973 17187
rect 25409 17147 25467 17153
rect 25516 17156 25973 17184
rect 24228 17088 24716 17116
rect 23385 17079 23443 17085
rect 25222 17076 25228 17128
rect 25280 17076 25286 17128
rect 18831 17020 19334 17048
rect 19429 17051 19487 17057
rect 18831 17017 18843 17020
rect 18785 17011 18843 17017
rect 19429 17017 19441 17051
rect 19475 17017 19487 17051
rect 19429 17011 19487 17017
rect 22066 17020 23612 17048
rect 19242 16940 19248 16992
rect 19300 16980 19306 16992
rect 22066 16980 22094 17020
rect 19300 16952 22094 16980
rect 19300 16940 19306 16952
rect 22738 16940 22744 16992
rect 22796 16980 22802 16992
rect 22925 16983 22983 16989
rect 22925 16980 22937 16983
rect 22796 16952 22937 16980
rect 22796 16940 22802 16952
rect 22925 16949 22937 16952
rect 22971 16949 22983 16983
rect 22925 16943 22983 16949
rect 23106 16940 23112 16992
rect 23164 16980 23170 16992
rect 23293 16983 23351 16989
rect 23293 16980 23305 16983
rect 23164 16952 23305 16980
rect 23164 16940 23170 16952
rect 23293 16949 23305 16952
rect 23339 16949 23351 16983
rect 23584 16980 23612 17020
rect 23658 17008 23664 17060
rect 23716 17048 23722 17060
rect 25516 17048 25544 17156
rect 25961 17153 25973 17156
rect 26007 17153 26019 17187
rect 25961 17147 26019 17153
rect 26145 17187 26203 17193
rect 26145 17153 26157 17187
rect 26191 17153 26203 17187
rect 26145 17147 26203 17153
rect 27525 17187 27583 17193
rect 27525 17153 27537 17187
rect 27571 17184 27583 17187
rect 27890 17184 27896 17196
rect 27571 17156 27896 17184
rect 27571 17153 27583 17156
rect 27525 17147 27583 17153
rect 27890 17144 27896 17156
rect 27948 17144 27954 17196
rect 29641 17187 29699 17193
rect 29641 17153 29653 17187
rect 29687 17184 29699 17187
rect 29822 17184 29828 17196
rect 29687 17156 29828 17184
rect 29687 17153 29699 17156
rect 29641 17147 29699 17153
rect 29822 17144 29828 17156
rect 29880 17144 29886 17196
rect 29914 17144 29920 17196
rect 29972 17144 29978 17196
rect 30556 17187 30614 17193
rect 30556 17153 30568 17187
rect 30602 17153 30614 17187
rect 30556 17147 30614 17153
rect 25685 17119 25743 17125
rect 25685 17085 25697 17119
rect 25731 17116 25743 17119
rect 26326 17116 26332 17128
rect 25731 17088 26332 17116
rect 25731 17085 25743 17088
rect 25685 17079 25743 17085
rect 26326 17076 26332 17088
rect 26384 17076 26390 17128
rect 26418 17076 26424 17128
rect 26476 17116 26482 17128
rect 27709 17119 27767 17125
rect 27709 17116 27721 17119
rect 26476 17088 27721 17116
rect 26476 17076 26482 17088
rect 27709 17085 27721 17088
rect 27755 17085 27767 17119
rect 27709 17079 27767 17085
rect 27798 17076 27804 17128
rect 27856 17076 27862 17128
rect 29362 17076 29368 17128
rect 29420 17116 29426 17128
rect 30571 17116 30599 17147
rect 30650 17144 30656 17196
rect 30708 17144 30714 17196
rect 30944 17193 30972 17224
rect 31481 17221 31493 17224
rect 31527 17252 31539 17255
rect 32122 17252 32128 17264
rect 31527 17224 32128 17252
rect 31527 17221 31539 17224
rect 31481 17215 31539 17221
rect 32122 17212 32128 17224
rect 32180 17212 32186 17264
rect 30928 17187 30986 17193
rect 30928 17153 30940 17187
rect 30974 17153 30986 17187
rect 30928 17147 30986 17153
rect 31018 17144 31024 17196
rect 31076 17144 31082 17196
rect 31110 17144 31116 17196
rect 31168 17144 31174 17196
rect 31202 17144 31208 17196
rect 31260 17144 31266 17196
rect 31386 17144 31392 17196
rect 31444 17144 31450 17196
rect 31662 17193 31668 17196
rect 31619 17187 31668 17193
rect 31619 17153 31631 17187
rect 31665 17153 31668 17187
rect 31619 17147 31668 17153
rect 31662 17144 31668 17147
rect 31720 17184 31726 17196
rect 33336 17184 33364 17292
rect 33778 17212 33784 17264
rect 33836 17212 33842 17264
rect 34238 17212 34244 17264
rect 34296 17212 34302 17264
rect 35084 17252 35112 17292
rect 35158 17280 35164 17332
rect 35216 17320 35222 17332
rect 35713 17323 35771 17329
rect 35713 17320 35725 17323
rect 35216 17292 35725 17320
rect 35216 17280 35222 17292
rect 35713 17289 35725 17292
rect 35759 17289 35771 17323
rect 36078 17320 36084 17332
rect 35713 17283 35771 17289
rect 35912 17292 36084 17320
rect 35084 17224 35756 17252
rect 35728 17196 35756 17224
rect 35912 17196 35940 17292
rect 36078 17280 36084 17292
rect 36136 17320 36142 17332
rect 36814 17320 36820 17332
rect 36136 17292 36820 17320
rect 36136 17280 36142 17292
rect 36814 17280 36820 17292
rect 36872 17280 36878 17332
rect 37182 17280 37188 17332
rect 37240 17320 37246 17332
rect 37277 17323 37335 17329
rect 37277 17320 37289 17323
rect 37240 17292 37289 17320
rect 37240 17280 37246 17292
rect 37277 17289 37289 17292
rect 37323 17320 37335 17323
rect 37645 17323 37703 17329
rect 37645 17320 37657 17323
rect 37323 17292 37657 17320
rect 37323 17289 37335 17292
rect 37277 17283 37335 17289
rect 37645 17289 37657 17292
rect 37691 17289 37703 17323
rect 37645 17283 37703 17289
rect 38102 17280 38108 17332
rect 38160 17280 38166 17332
rect 38930 17280 38936 17332
rect 38988 17320 38994 17332
rect 39209 17323 39267 17329
rect 38988 17292 39068 17320
rect 38988 17280 38994 17292
rect 39040 17252 39068 17292
rect 39209 17289 39221 17323
rect 39255 17320 39267 17323
rect 39298 17320 39304 17332
rect 39255 17292 39304 17320
rect 39255 17289 39267 17292
rect 39209 17283 39267 17289
rect 39298 17280 39304 17292
rect 39356 17280 39362 17332
rect 39758 17280 39764 17332
rect 39816 17280 39822 17332
rect 40402 17280 40408 17332
rect 40460 17280 40466 17332
rect 40586 17280 40592 17332
rect 40644 17280 40650 17332
rect 40678 17280 40684 17332
rect 40736 17320 40742 17332
rect 41233 17323 41291 17329
rect 41233 17320 41245 17323
rect 40736 17292 41245 17320
rect 40736 17280 40742 17292
rect 41233 17289 41245 17292
rect 41279 17289 41291 17323
rect 41233 17283 41291 17289
rect 41509 17323 41567 17329
rect 41509 17289 41521 17323
rect 41555 17320 41567 17323
rect 41966 17320 41972 17332
rect 41555 17292 41972 17320
rect 41555 17289 41567 17292
rect 41509 17283 41567 17289
rect 41966 17280 41972 17292
rect 42024 17280 42030 17332
rect 42981 17323 43039 17329
rect 42981 17289 42993 17323
rect 43027 17320 43039 17323
rect 43070 17320 43076 17332
rect 43027 17292 43076 17320
rect 43027 17289 43039 17292
rect 42981 17283 43039 17289
rect 43070 17280 43076 17292
rect 43128 17280 43134 17332
rect 43349 17323 43407 17329
rect 43349 17289 43361 17323
rect 43395 17320 43407 17323
rect 43898 17320 43904 17332
rect 43395 17292 43904 17320
rect 43395 17289 43407 17292
rect 43349 17283 43407 17289
rect 39776 17252 39804 17280
rect 39040 17224 39804 17252
rect 40221 17255 40279 17261
rect 40221 17221 40233 17255
rect 40267 17252 40279 17255
rect 40420 17252 40448 17280
rect 41138 17252 41144 17264
rect 40267 17224 41144 17252
rect 40267 17221 40279 17224
rect 40221 17215 40279 17221
rect 41138 17212 41144 17224
rect 41196 17212 41202 17264
rect 42610 17212 42616 17264
rect 42668 17212 42674 17264
rect 42702 17212 42708 17264
rect 42760 17212 42766 17264
rect 31720 17156 33364 17184
rect 31720 17144 31726 17156
rect 33502 17144 33508 17196
rect 33560 17144 33566 17196
rect 35621 17187 35679 17193
rect 35621 17184 35633 17187
rect 35176 17156 35633 17184
rect 30742 17116 30748 17128
rect 29420 17088 30512 17116
rect 30571 17088 30748 17116
rect 29420 17076 29426 17088
rect 23716 17020 25544 17048
rect 25777 17051 25835 17057
rect 23716 17008 23722 17020
rect 25777 17017 25789 17051
rect 25823 17048 25835 17051
rect 30377 17051 30435 17057
rect 30377 17048 30389 17051
rect 25823 17020 30389 17048
rect 25823 17017 25835 17020
rect 25777 17011 25835 17017
rect 30377 17017 30389 17020
rect 30423 17017 30435 17051
rect 30484 17048 30512 17088
rect 30742 17076 30748 17088
rect 30800 17076 30806 17128
rect 34514 17076 34520 17128
rect 34572 17116 34578 17128
rect 35176 17116 35204 17156
rect 35621 17153 35633 17156
rect 35667 17153 35679 17187
rect 35621 17147 35679 17153
rect 35710 17144 35716 17196
rect 35768 17144 35774 17196
rect 35894 17144 35900 17196
rect 35952 17144 35958 17196
rect 35989 17187 36047 17193
rect 35989 17153 36001 17187
rect 36035 17153 36047 17187
rect 35989 17147 36047 17153
rect 34572 17088 35204 17116
rect 34572 17076 34578 17088
rect 35250 17076 35256 17128
rect 35308 17076 35314 17128
rect 35526 17076 35532 17128
rect 35584 17116 35590 17128
rect 36004 17116 36032 17147
rect 36078 17144 36084 17196
rect 36136 17144 36142 17196
rect 36265 17187 36323 17193
rect 36265 17153 36277 17187
rect 36311 17184 36323 17187
rect 36538 17184 36544 17196
rect 36311 17156 36544 17184
rect 36311 17153 36323 17156
rect 36265 17147 36323 17153
rect 36538 17144 36544 17156
rect 36596 17144 36602 17196
rect 38289 17187 38347 17193
rect 38289 17153 38301 17187
rect 38335 17184 38347 17187
rect 38335 17156 38700 17184
rect 38335 17153 38347 17156
rect 38289 17147 38347 17153
rect 35584 17088 36032 17116
rect 35584 17076 35590 17088
rect 37274 17076 37280 17128
rect 37332 17116 37338 17128
rect 37461 17119 37519 17125
rect 37461 17116 37473 17119
rect 37332 17088 37473 17116
rect 37332 17076 37338 17088
rect 37461 17085 37473 17088
rect 37507 17085 37519 17119
rect 37461 17079 37519 17085
rect 31202 17048 31208 17060
rect 30484 17020 31208 17048
rect 30377 17011 30435 17017
rect 31202 17008 31208 17020
rect 31260 17008 31266 17060
rect 31680 17020 33640 17048
rect 24210 16980 24216 16992
rect 23584 16952 24216 16980
rect 23293 16943 23351 16949
rect 24210 16940 24216 16952
rect 24268 16940 24274 16992
rect 24394 16940 24400 16992
rect 24452 16980 24458 16992
rect 24581 16983 24639 16989
rect 24581 16980 24593 16983
rect 24452 16952 24593 16980
rect 24452 16940 24458 16952
rect 24581 16949 24593 16952
rect 24627 16949 24639 16983
rect 24581 16943 24639 16949
rect 25317 16983 25375 16989
rect 25317 16949 25329 16983
rect 25363 16980 25375 16983
rect 25406 16980 25412 16992
rect 25363 16952 25412 16980
rect 25363 16949 25375 16952
rect 25317 16943 25375 16949
rect 25406 16940 25412 16952
rect 25464 16940 25470 16992
rect 25866 16940 25872 16992
rect 25924 16940 25930 16992
rect 27246 16940 27252 16992
rect 27304 16980 27310 16992
rect 27341 16983 27399 16989
rect 27341 16980 27353 16983
rect 27304 16952 27353 16980
rect 27304 16940 27310 16952
rect 27341 16949 27353 16952
rect 27387 16949 27399 16983
rect 27341 16943 27399 16949
rect 29454 16940 29460 16992
rect 29512 16940 29518 16992
rect 29638 16940 29644 16992
rect 29696 16980 29702 16992
rect 29825 16983 29883 16989
rect 29825 16980 29837 16983
rect 29696 16952 29837 16980
rect 29696 16940 29702 16952
rect 29825 16949 29837 16952
rect 29871 16949 29883 16983
rect 29825 16943 29883 16949
rect 30101 16983 30159 16989
rect 30101 16949 30113 16983
rect 30147 16980 30159 16983
rect 30282 16980 30288 16992
rect 30147 16952 30288 16980
rect 30147 16949 30159 16952
rect 30101 16943 30159 16949
rect 30282 16940 30288 16952
rect 30340 16980 30346 16992
rect 31680 16980 31708 17020
rect 30340 16952 31708 16980
rect 30340 16940 30346 16952
rect 31754 16940 31760 16992
rect 31812 16940 31818 16992
rect 31846 16940 31852 16992
rect 31904 16940 31910 16992
rect 33612 16980 33640 17020
rect 34882 17008 34888 17060
rect 34940 17048 34946 17060
rect 35437 17051 35495 17057
rect 35437 17048 35449 17051
rect 34940 17020 35449 17048
rect 34940 17008 34946 17020
rect 35437 17017 35449 17020
rect 35483 17048 35495 17051
rect 36170 17048 36176 17060
rect 35483 17020 36176 17048
rect 35483 17017 35495 17020
rect 35437 17011 35495 17017
rect 36170 17008 36176 17020
rect 36228 17008 36234 17060
rect 36538 17008 36544 17060
rect 36596 17048 36602 17060
rect 36725 17051 36783 17057
rect 36725 17048 36737 17051
rect 36596 17020 36737 17048
rect 36596 17008 36602 17020
rect 36725 17017 36737 17020
rect 36771 17017 36783 17051
rect 36725 17011 36783 17017
rect 38672 16992 38700 17156
rect 38746 17144 38752 17196
rect 38804 17144 38810 17196
rect 38933 17187 38991 17193
rect 38933 17153 38945 17187
rect 38979 17184 38991 17187
rect 39025 17187 39083 17193
rect 39025 17184 39037 17187
rect 38979 17156 39037 17184
rect 38979 17153 38991 17156
rect 38933 17147 38991 17153
rect 39025 17153 39037 17156
rect 39071 17184 39083 17187
rect 39485 17187 39543 17193
rect 39485 17184 39497 17187
rect 39071 17156 39497 17184
rect 39071 17153 39083 17156
rect 39025 17147 39083 17153
rect 39485 17153 39497 17156
rect 39531 17184 39543 17187
rect 39669 17187 39727 17193
rect 39669 17184 39681 17187
rect 39531 17156 39681 17184
rect 39531 17153 39543 17156
rect 39485 17147 39543 17153
rect 39669 17153 39681 17156
rect 39715 17184 39727 17187
rect 39758 17184 39764 17196
rect 39715 17156 39764 17184
rect 39715 17153 39727 17156
rect 39669 17147 39727 17153
rect 39758 17144 39764 17156
rect 39816 17144 39822 17196
rect 39942 17144 39948 17196
rect 40000 17144 40006 17196
rect 40093 17187 40151 17193
rect 40093 17153 40105 17187
rect 40139 17184 40151 17187
rect 40139 17153 40172 17184
rect 40093 17147 40172 17153
rect 40144 17116 40172 17147
rect 40310 17144 40316 17196
rect 40368 17144 40374 17196
rect 40451 17187 40509 17193
rect 40451 17153 40463 17187
rect 40497 17184 40509 17187
rect 40862 17184 40868 17196
rect 40497 17156 40868 17184
rect 40497 17153 40509 17156
rect 40451 17147 40509 17153
rect 40862 17144 40868 17156
rect 40920 17144 40926 17196
rect 41046 17144 41052 17196
rect 41104 17184 41110 17196
rect 41104 17156 41414 17184
rect 41104 17144 41110 17156
rect 40586 17116 40592 17128
rect 40144 17088 40592 17116
rect 40586 17076 40592 17088
rect 40644 17076 40650 17128
rect 41064 17116 41092 17144
rect 40788 17088 41092 17116
rect 41386 17116 41414 17156
rect 42334 17144 42340 17196
rect 42392 17184 42398 17196
rect 42429 17187 42487 17193
rect 42429 17184 42441 17187
rect 42392 17156 42441 17184
rect 42392 17144 42398 17156
rect 42429 17153 42441 17156
rect 42475 17153 42487 17187
rect 42429 17147 42487 17153
rect 42797 17187 42855 17193
rect 42797 17153 42809 17187
rect 42843 17184 42855 17187
rect 43364 17184 43392 17283
rect 43898 17280 43904 17292
rect 43956 17280 43962 17332
rect 44082 17280 44088 17332
rect 44140 17280 44146 17332
rect 44542 17280 44548 17332
rect 44600 17320 44606 17332
rect 44600 17292 45048 17320
rect 44600 17280 44606 17292
rect 44100 17252 44128 17280
rect 45020 17252 45048 17292
rect 46750 17280 46756 17332
rect 46808 17320 46814 17332
rect 47581 17323 47639 17329
rect 47581 17320 47593 17323
rect 46808 17292 47593 17320
rect 46808 17280 46814 17292
rect 47581 17289 47593 17292
rect 47627 17289 47639 17323
rect 47581 17283 47639 17289
rect 49050 17280 49056 17332
rect 49108 17320 49114 17332
rect 49108 17292 49280 17320
rect 49108 17280 49114 17292
rect 46566 17252 46572 17264
rect 44100 17224 44206 17252
rect 45020 17224 46572 17252
rect 46566 17212 46572 17224
rect 46624 17252 46630 17264
rect 48498 17252 48504 17264
rect 46624 17224 47072 17252
rect 46624 17212 46630 17224
rect 42843 17156 43392 17184
rect 42843 17153 42855 17156
rect 42797 17147 42855 17153
rect 46014 17144 46020 17196
rect 46072 17144 46078 17196
rect 46198 17193 46204 17196
rect 46165 17187 46204 17193
rect 46165 17153 46177 17187
rect 46165 17147 46204 17153
rect 46198 17144 46204 17147
rect 46256 17144 46262 17196
rect 46290 17144 46296 17196
rect 46348 17144 46354 17196
rect 46385 17187 46443 17193
rect 46385 17153 46397 17187
rect 46431 17153 46443 17187
rect 46385 17147 46443 17153
rect 42978 17116 42984 17128
rect 41386 17088 42984 17116
rect 39390 17008 39396 17060
rect 39448 17048 39454 17060
rect 40681 17051 40739 17057
rect 40681 17048 40693 17051
rect 39448 17020 40693 17048
rect 39448 17008 39454 17020
rect 40681 17017 40693 17020
rect 40727 17017 40739 17051
rect 40681 17011 40739 17017
rect 35894 16980 35900 16992
rect 33612 16952 35900 16980
rect 35894 16940 35900 16952
rect 35952 16940 35958 16992
rect 36630 16940 36636 16992
rect 36688 16940 36694 16992
rect 38470 16940 38476 16992
rect 38528 16940 38534 16992
rect 38654 16940 38660 16992
rect 38712 16980 38718 16992
rect 40788 16980 40816 17088
rect 42978 17076 42984 17088
rect 43036 17076 43042 17128
rect 43438 17076 43444 17128
rect 43496 17076 43502 17128
rect 43717 17119 43775 17125
rect 43717 17085 43729 17119
rect 43763 17116 43775 17119
rect 43806 17116 43812 17128
rect 43763 17088 43812 17116
rect 43763 17085 43775 17088
rect 43717 17079 43775 17085
rect 43806 17076 43812 17088
rect 43864 17076 43870 17128
rect 45833 17119 45891 17125
rect 45833 17116 45845 17119
rect 45204 17088 45845 17116
rect 40862 17008 40868 17060
rect 40920 17048 40926 17060
rect 41598 17048 41604 17060
rect 40920 17020 41604 17048
rect 40920 17008 40926 17020
rect 41598 17008 41604 17020
rect 41656 17008 41662 17060
rect 41782 17008 41788 17060
rect 41840 17048 41846 17060
rect 42610 17048 42616 17060
rect 41840 17020 42616 17048
rect 41840 17008 41846 17020
rect 42610 17008 42616 17020
rect 42668 17048 42674 17060
rect 43073 17051 43131 17057
rect 43073 17048 43085 17051
rect 42668 17020 43085 17048
rect 42668 17008 42674 17020
rect 43073 17017 43085 17020
rect 43119 17017 43131 17051
rect 43073 17011 43131 17017
rect 38712 16952 40816 16980
rect 38712 16940 38718 16952
rect 43530 16940 43536 16992
rect 43588 16980 43594 16992
rect 45204 16989 45232 17088
rect 45833 17085 45845 17088
rect 45879 17085 45891 17119
rect 46400 17116 46428 17147
rect 46474 17144 46480 17196
rect 46532 17193 46538 17196
rect 47044 17193 47072 17224
rect 47780 17224 48504 17252
rect 47780 17193 47808 17224
rect 48498 17212 48504 17224
rect 48556 17212 48562 17264
rect 49252 17261 49280 17292
rect 49510 17280 49516 17332
rect 49568 17280 49574 17332
rect 49694 17280 49700 17332
rect 49752 17280 49758 17332
rect 49786 17280 49792 17332
rect 49844 17320 49850 17332
rect 50433 17323 50491 17329
rect 50433 17320 50445 17323
rect 49844 17292 50445 17320
rect 49844 17280 49850 17292
rect 50433 17289 50445 17292
rect 50479 17289 50491 17323
rect 50433 17283 50491 17289
rect 50614 17280 50620 17332
rect 50672 17280 50678 17332
rect 53006 17280 53012 17332
rect 53064 17320 53070 17332
rect 53285 17323 53343 17329
rect 53285 17320 53297 17323
rect 53064 17292 53297 17320
rect 53064 17280 53070 17292
rect 53285 17289 53297 17292
rect 53331 17289 53343 17323
rect 53285 17283 53343 17289
rect 53466 17280 53472 17332
rect 53524 17320 53530 17332
rect 54021 17323 54079 17329
rect 53524 17292 53696 17320
rect 53524 17280 53530 17292
rect 48685 17255 48743 17261
rect 48685 17221 48697 17255
rect 48731 17252 48743 17255
rect 49145 17255 49203 17261
rect 49145 17252 49157 17255
rect 48731 17224 49157 17252
rect 48731 17221 48743 17224
rect 48685 17215 48743 17221
rect 49145 17221 49157 17224
rect 49191 17221 49203 17255
rect 49145 17215 49203 17221
rect 49237 17255 49295 17261
rect 49237 17221 49249 17255
rect 49283 17221 49295 17255
rect 49237 17215 49295 17221
rect 46532 17184 46540 17193
rect 47029 17187 47087 17193
rect 46532 17156 46577 17184
rect 46532 17147 46540 17156
rect 47029 17153 47041 17187
rect 47075 17153 47087 17187
rect 47029 17147 47087 17153
rect 47765 17187 47823 17193
rect 47765 17153 47777 17187
rect 47811 17153 47823 17187
rect 47765 17147 47823 17153
rect 47857 17187 47915 17193
rect 47857 17153 47869 17187
rect 47903 17153 47915 17187
rect 47857 17147 47915 17153
rect 48133 17187 48191 17193
rect 48133 17153 48145 17187
rect 48179 17184 48191 17187
rect 48314 17184 48320 17196
rect 48179 17156 48320 17184
rect 48179 17153 48191 17156
rect 48133 17147 48191 17153
rect 46532 17144 46538 17147
rect 46845 17119 46903 17125
rect 46845 17116 46857 17119
rect 46400 17088 46857 17116
rect 45833 17079 45891 17085
rect 46845 17085 46857 17088
rect 46891 17085 46903 17119
rect 46845 17079 46903 17085
rect 47213 17119 47271 17125
rect 47213 17085 47225 17119
rect 47259 17116 47271 17119
rect 47872 17116 47900 17147
rect 48314 17144 48320 17156
rect 48372 17144 48378 17196
rect 48866 17144 48872 17196
rect 48924 17144 48930 17196
rect 49050 17193 49056 17196
rect 49017 17187 49056 17193
rect 49017 17153 49029 17187
rect 49017 17147 49056 17153
rect 49050 17144 49056 17147
rect 49108 17144 49114 17196
rect 47259 17088 47900 17116
rect 48041 17119 48099 17125
rect 47259 17085 47271 17088
rect 47213 17079 47271 17085
rect 48041 17085 48053 17119
rect 48087 17116 48099 17119
rect 48774 17116 48780 17128
rect 48087 17088 48780 17116
rect 48087 17085 48099 17088
rect 48041 17079 48099 17085
rect 46860 17048 46888 17079
rect 48774 17076 48780 17088
rect 48832 17076 48838 17128
rect 49160 17116 49188 17215
rect 49326 17144 49332 17196
rect 49384 17193 49390 17196
rect 49384 17184 49392 17193
rect 49804 17184 49832 17280
rect 50062 17212 50068 17264
rect 50120 17212 50126 17264
rect 53374 17252 53380 17264
rect 50264 17224 53380 17252
rect 50264 17196 50292 17224
rect 53374 17212 53380 17224
rect 53432 17252 53438 17264
rect 53668 17261 53696 17292
rect 54021 17289 54033 17323
rect 54067 17320 54079 17323
rect 54570 17320 54576 17332
rect 54067 17292 54576 17320
rect 54067 17289 54079 17292
rect 54021 17283 54079 17289
rect 54570 17280 54576 17292
rect 54628 17280 54634 17332
rect 55766 17280 55772 17332
rect 55824 17320 55830 17332
rect 55861 17323 55919 17329
rect 55861 17320 55873 17323
rect 55824 17292 55873 17320
rect 55824 17280 55830 17292
rect 55861 17289 55873 17292
rect 55907 17289 55919 17323
rect 56870 17320 56876 17332
rect 55861 17283 55919 17289
rect 55968 17292 56876 17320
rect 53653 17255 53711 17261
rect 53432 17224 53512 17252
rect 53432 17212 53438 17224
rect 49876 17187 49934 17193
rect 49876 17184 49888 17187
rect 49384 17156 49429 17184
rect 49804 17156 49888 17184
rect 49384 17147 49392 17156
rect 49876 17153 49888 17156
rect 49922 17153 49934 17187
rect 49876 17147 49934 17153
rect 49973 17187 50031 17193
rect 49973 17153 49985 17187
rect 50019 17153 50031 17187
rect 50246 17184 50252 17196
rect 50207 17156 50252 17184
rect 49973 17147 50031 17153
rect 49384 17144 49390 17147
rect 49786 17116 49792 17128
rect 49160 17088 49792 17116
rect 49786 17076 49792 17088
rect 49844 17076 49850 17128
rect 49988 17116 50016 17147
rect 50246 17144 50252 17156
rect 50304 17144 50310 17196
rect 50338 17144 50344 17196
rect 50396 17144 50402 17196
rect 50798 17144 50804 17196
rect 50856 17144 50862 17196
rect 50890 17144 50896 17196
rect 50948 17144 50954 17196
rect 51169 17187 51227 17193
rect 51169 17153 51181 17187
rect 51215 17184 51227 17187
rect 51537 17187 51595 17193
rect 51537 17184 51549 17187
rect 51215 17156 51549 17184
rect 51215 17153 51227 17156
rect 51169 17147 51227 17153
rect 51537 17153 51549 17156
rect 51583 17153 51595 17187
rect 51537 17147 51595 17153
rect 51626 17144 51632 17196
rect 51684 17184 51690 17196
rect 52089 17187 52147 17193
rect 52089 17184 52101 17187
rect 51684 17156 52101 17184
rect 51684 17144 51690 17156
rect 52089 17153 52101 17156
rect 52135 17184 52147 17187
rect 52362 17184 52368 17196
rect 52135 17156 52368 17184
rect 52135 17153 52147 17156
rect 52089 17147 52147 17153
rect 52362 17144 52368 17156
rect 52420 17184 52426 17196
rect 52733 17187 52791 17193
rect 52733 17184 52745 17187
rect 52420 17156 52745 17184
rect 52420 17144 52426 17156
rect 52733 17153 52745 17156
rect 52779 17153 52791 17187
rect 52733 17147 52791 17153
rect 52914 17144 52920 17196
rect 52972 17144 52978 17196
rect 53006 17144 53012 17196
rect 53064 17144 53070 17196
rect 53101 17187 53159 17193
rect 53101 17153 53113 17187
rect 53147 17184 53159 17187
rect 53190 17184 53196 17196
rect 53147 17156 53196 17184
rect 53147 17153 53159 17156
rect 53101 17147 53159 17153
rect 53190 17144 53196 17156
rect 53248 17144 53254 17196
rect 53484 17193 53512 17224
rect 53653 17221 53665 17255
rect 53699 17221 53711 17255
rect 53653 17215 53711 17221
rect 54386 17212 54392 17264
rect 54444 17212 54450 17264
rect 54846 17212 54852 17264
rect 54904 17212 54910 17264
rect 53742 17193 53748 17196
rect 53469 17187 53527 17193
rect 53469 17153 53481 17187
rect 53515 17153 53527 17187
rect 53737 17184 53748 17193
rect 53469 17147 53527 17153
rect 53668 17156 53748 17184
rect 53668 17116 53696 17156
rect 53737 17147 53748 17156
rect 53742 17144 53748 17147
rect 53800 17144 53806 17196
rect 53837 17187 53895 17193
rect 53837 17153 53849 17187
rect 53883 17153 53895 17187
rect 53837 17147 53895 17153
rect 49988 17088 53696 17116
rect 51534 17048 51540 17060
rect 46860 17020 51540 17048
rect 51534 17008 51540 17020
rect 51592 17008 51598 17060
rect 51810 17008 51816 17060
rect 51868 17048 51874 17060
rect 53190 17048 53196 17060
rect 51868 17020 53196 17048
rect 51868 17008 51874 17020
rect 53190 17008 53196 17020
rect 53248 17048 53254 17060
rect 53558 17048 53564 17060
rect 53248 17020 53564 17048
rect 53248 17008 53254 17020
rect 53558 17008 53564 17020
rect 53616 17048 53622 17060
rect 53852 17048 53880 17147
rect 53926 17076 53932 17128
rect 53984 17116 53990 17128
rect 55968 17125 55996 17292
rect 56870 17280 56876 17292
rect 56928 17280 56934 17332
rect 56226 17212 56232 17264
rect 56284 17212 56290 17264
rect 56778 17212 56784 17264
rect 56836 17212 56842 17264
rect 54113 17119 54171 17125
rect 54113 17116 54125 17119
rect 53984 17088 54125 17116
rect 53984 17076 53990 17088
rect 54113 17085 54125 17088
rect 54159 17116 54171 17119
rect 55953 17119 56011 17125
rect 55953 17116 55965 17119
rect 54159 17088 55965 17116
rect 54159 17085 54171 17088
rect 54113 17079 54171 17085
rect 55953 17085 55965 17088
rect 55999 17085 56011 17119
rect 55953 17079 56011 17085
rect 56686 17076 56692 17128
rect 56744 17116 56750 17128
rect 57514 17116 57520 17128
rect 56744 17088 57520 17116
rect 56744 17076 56750 17088
rect 57514 17076 57520 17088
rect 57572 17116 57578 17128
rect 57701 17119 57759 17125
rect 57701 17116 57713 17119
rect 57572 17088 57713 17116
rect 57572 17076 57578 17088
rect 57701 17085 57713 17088
rect 57747 17085 57759 17119
rect 57701 17079 57759 17085
rect 53616 17020 53880 17048
rect 53616 17008 53622 17020
rect 45189 16983 45247 16989
rect 45189 16980 45201 16983
rect 43588 16952 45201 16980
rect 43588 16940 43594 16952
rect 45189 16949 45201 16952
rect 45235 16949 45247 16983
rect 45189 16943 45247 16949
rect 45278 16940 45284 16992
rect 45336 16940 45342 16992
rect 46661 16983 46719 16989
rect 46661 16949 46673 16983
rect 46707 16980 46719 16983
rect 47486 16980 47492 16992
rect 46707 16952 47492 16980
rect 46707 16949 46719 16952
rect 46661 16943 46719 16949
rect 47486 16940 47492 16952
rect 47544 16940 47550 16992
rect 48314 16940 48320 16992
rect 48372 16940 48378 16992
rect 48498 16940 48504 16992
rect 48556 16940 48562 16992
rect 51074 16940 51080 16992
rect 51132 16980 51138 16992
rect 51258 16980 51264 16992
rect 51132 16952 51264 16980
rect 51132 16940 51138 16952
rect 51258 16940 51264 16952
rect 51316 16940 51322 16992
rect 52914 16940 52920 16992
rect 52972 16980 52978 16992
rect 53466 16980 53472 16992
rect 52972 16952 53472 16980
rect 52972 16940 52978 16952
rect 53466 16940 53472 16952
rect 53524 16940 53530 16992
rect 1104 16890 58880 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 58880 16890
rect 1104 16816 58880 16838
rect 22636 16779 22694 16785
rect 22636 16745 22648 16779
rect 22682 16776 22694 16779
rect 22738 16776 22744 16788
rect 22682 16748 22744 16776
rect 22682 16745 22694 16748
rect 22636 16739 22694 16745
rect 22738 16736 22744 16748
rect 22796 16736 22802 16788
rect 23014 16736 23020 16788
rect 23072 16776 23078 16788
rect 24121 16779 24179 16785
rect 24121 16776 24133 16779
rect 23072 16748 24133 16776
rect 23072 16736 23078 16748
rect 24121 16745 24133 16748
rect 24167 16776 24179 16779
rect 25038 16776 25044 16788
rect 24167 16748 25044 16776
rect 24167 16745 24179 16748
rect 24121 16739 24179 16745
rect 25038 16736 25044 16748
rect 25096 16736 25102 16788
rect 25133 16779 25191 16785
rect 25133 16745 25145 16779
rect 25179 16776 25191 16779
rect 25314 16776 25320 16788
rect 25179 16748 25320 16776
rect 25179 16745 25191 16748
rect 25133 16739 25191 16745
rect 19245 16711 19303 16717
rect 19245 16677 19257 16711
rect 19291 16677 19303 16711
rect 19245 16671 19303 16677
rect 16666 16600 16672 16652
rect 16724 16600 16730 16652
rect 16945 16643 17003 16649
rect 16945 16609 16957 16643
rect 16991 16640 17003 16643
rect 18509 16643 18567 16649
rect 18509 16640 18521 16643
rect 16991 16612 18521 16640
rect 16991 16609 17003 16612
rect 16945 16603 17003 16609
rect 18509 16609 18521 16612
rect 18555 16609 18567 16643
rect 19260 16640 19288 16671
rect 18509 16603 18567 16609
rect 18708 16612 19288 16640
rect 18708 16581 18736 16612
rect 19518 16600 19524 16652
rect 19576 16640 19582 16652
rect 20533 16643 20591 16649
rect 19576 16612 19932 16640
rect 19576 16600 19582 16612
rect 18693 16575 18751 16581
rect 18693 16541 18705 16575
rect 18739 16541 18751 16575
rect 18693 16535 18751 16541
rect 18874 16532 18880 16584
rect 18932 16532 18938 16584
rect 18966 16532 18972 16584
rect 19024 16532 19030 16584
rect 19424 16575 19482 16581
rect 19424 16541 19436 16575
rect 19470 16572 19482 16575
rect 19702 16572 19708 16584
rect 19470 16544 19708 16572
rect 19470 16541 19482 16544
rect 19424 16535 19482 16541
rect 19702 16532 19708 16544
rect 19760 16532 19766 16584
rect 19904 16581 19932 16612
rect 20533 16609 20545 16643
rect 20579 16640 20591 16643
rect 22186 16640 22192 16652
rect 20579 16612 22192 16640
rect 20579 16609 20591 16612
rect 20533 16603 20591 16609
rect 22186 16600 22192 16612
rect 22244 16640 22250 16652
rect 22373 16643 22431 16649
rect 22373 16640 22385 16643
rect 22244 16612 22385 16640
rect 22244 16600 22250 16612
rect 22373 16609 22385 16612
rect 22419 16640 22431 16643
rect 24118 16640 24124 16652
rect 22419 16612 24124 16640
rect 22419 16609 22431 16612
rect 22373 16603 22431 16609
rect 24118 16600 24124 16612
rect 24176 16600 24182 16652
rect 25148 16640 25176 16739
rect 25314 16736 25320 16748
rect 25372 16736 25378 16788
rect 25866 16736 25872 16788
rect 25924 16736 25930 16788
rect 25958 16736 25964 16788
rect 26016 16776 26022 16788
rect 26053 16779 26111 16785
rect 26053 16776 26065 16779
rect 26016 16748 26065 16776
rect 26016 16736 26022 16748
rect 26053 16745 26065 16748
rect 26099 16776 26111 16779
rect 26878 16776 26884 16788
rect 26099 16748 26884 16776
rect 26099 16745 26111 16748
rect 26053 16739 26111 16745
rect 26878 16736 26884 16748
rect 26936 16736 26942 16788
rect 27798 16736 27804 16788
rect 27856 16776 27862 16788
rect 28721 16779 28779 16785
rect 28721 16776 28733 16779
rect 27856 16748 28733 16776
rect 27856 16736 27862 16748
rect 28721 16745 28733 16748
rect 28767 16776 28779 16779
rect 28767 16748 28994 16776
rect 28767 16745 28779 16748
rect 28721 16739 28779 16745
rect 25222 16668 25228 16720
rect 25280 16708 25286 16720
rect 26329 16711 26387 16717
rect 26329 16708 26341 16711
rect 25280 16680 26341 16708
rect 25280 16668 25286 16680
rect 26329 16677 26341 16680
rect 26375 16677 26387 16711
rect 26329 16671 26387 16677
rect 24688 16612 25176 16640
rect 19796 16575 19854 16581
rect 19796 16541 19808 16575
rect 19842 16541 19854 16575
rect 19796 16535 19854 16541
rect 19889 16575 19947 16581
rect 19889 16541 19901 16575
rect 19935 16572 19947 16575
rect 20346 16572 20352 16584
rect 19935 16544 20352 16572
rect 19935 16541 19947 16544
rect 19889 16535 19947 16541
rect 17954 16464 17960 16516
rect 18012 16464 18018 16516
rect 19334 16464 19340 16516
rect 19392 16504 19398 16516
rect 19521 16507 19579 16513
rect 19521 16504 19533 16507
rect 19392 16476 19533 16504
rect 19392 16464 19398 16476
rect 19521 16473 19533 16476
rect 19567 16473 19579 16507
rect 19521 16467 19579 16473
rect 18417 16439 18475 16445
rect 18417 16405 18429 16439
rect 18463 16436 18475 16439
rect 18966 16436 18972 16448
rect 18463 16408 18972 16436
rect 18463 16405 18475 16408
rect 18417 16399 18475 16405
rect 18966 16396 18972 16408
rect 19024 16396 19030 16448
rect 19536 16436 19564 16467
rect 19610 16464 19616 16516
rect 19668 16464 19674 16516
rect 19812 16504 19840 16535
rect 20346 16532 20352 16544
rect 20404 16532 20410 16584
rect 21910 16532 21916 16584
rect 21968 16572 21974 16584
rect 21968 16544 22140 16572
rect 21968 16532 21974 16544
rect 19978 16504 19984 16516
rect 19812 16476 19984 16504
rect 19978 16464 19984 16476
rect 20036 16464 20042 16516
rect 20806 16464 20812 16516
rect 20864 16464 20870 16516
rect 22112 16504 22140 16544
rect 24394 16532 24400 16584
rect 24452 16532 24458 16584
rect 24486 16532 24492 16584
rect 24544 16532 24550 16584
rect 24688 16581 24716 16612
rect 26418 16600 26424 16652
rect 26476 16640 26482 16652
rect 26476 16612 26648 16640
rect 26476 16600 26482 16612
rect 24673 16575 24731 16581
rect 24673 16541 24685 16575
rect 24719 16541 24731 16575
rect 24673 16535 24731 16541
rect 24903 16575 24961 16581
rect 24903 16541 24915 16575
rect 24949 16572 24961 16575
rect 25038 16572 25044 16584
rect 24949 16544 25044 16572
rect 24949 16541 24961 16544
rect 24903 16535 24961 16541
rect 25038 16532 25044 16544
rect 25096 16532 25102 16584
rect 25314 16532 25320 16584
rect 25372 16532 25378 16584
rect 25593 16575 25651 16581
rect 25593 16572 25605 16575
rect 25424 16544 25605 16572
rect 22112 16476 23138 16504
rect 24578 16464 24584 16516
rect 24636 16504 24642 16516
rect 24765 16507 24823 16513
rect 24765 16504 24777 16507
rect 24636 16476 24777 16504
rect 24636 16464 24642 16476
rect 24765 16473 24777 16476
rect 24811 16473 24823 16507
rect 25424 16504 25452 16544
rect 25593 16541 25605 16544
rect 25639 16541 25651 16575
rect 25593 16535 25651 16541
rect 25682 16532 25688 16584
rect 25740 16532 25746 16584
rect 25866 16532 25872 16584
rect 25924 16572 25930 16584
rect 26145 16575 26203 16581
rect 26145 16572 26157 16575
rect 25924 16544 26157 16572
rect 25924 16532 25930 16544
rect 26145 16541 26157 16544
rect 26191 16541 26203 16575
rect 26145 16535 26203 16541
rect 26234 16532 26240 16584
rect 26292 16572 26298 16584
rect 26620 16581 26648 16612
rect 26970 16600 26976 16652
rect 27028 16600 27034 16652
rect 27246 16600 27252 16652
rect 27304 16600 27310 16652
rect 28966 16640 28994 16748
rect 29822 16736 29828 16788
rect 29880 16776 29886 16788
rect 30193 16779 30251 16785
rect 30193 16776 30205 16779
rect 29880 16748 30205 16776
rect 29880 16736 29886 16748
rect 30193 16745 30205 16748
rect 30239 16745 30251 16779
rect 30193 16739 30251 16745
rect 30650 16736 30656 16788
rect 30708 16776 30714 16788
rect 30926 16776 30932 16788
rect 30708 16748 30932 16776
rect 30708 16736 30714 16748
rect 30926 16736 30932 16748
rect 30984 16736 30990 16788
rect 31018 16736 31024 16788
rect 31076 16776 31082 16788
rect 34238 16776 34244 16788
rect 31076 16748 34244 16776
rect 31076 16736 31082 16748
rect 34238 16736 34244 16748
rect 34296 16736 34302 16788
rect 35802 16736 35808 16788
rect 35860 16776 35866 16788
rect 35860 16748 35940 16776
rect 35860 16736 35866 16748
rect 30558 16708 30564 16720
rect 29840 16680 30564 16708
rect 28966 16612 29684 16640
rect 26513 16575 26571 16581
rect 26513 16572 26525 16575
rect 26292 16544 26525 16572
rect 26292 16532 26298 16544
rect 26513 16541 26525 16544
rect 26559 16541 26571 16575
rect 26513 16535 26571 16541
rect 26605 16575 26663 16581
rect 26605 16541 26617 16575
rect 26651 16541 26663 16575
rect 26605 16535 26663 16541
rect 24765 16467 24823 16473
rect 24872 16476 25452 16504
rect 22186 16436 22192 16448
rect 19536 16408 22192 16436
rect 22186 16396 22192 16408
rect 22244 16396 22250 16448
rect 22281 16439 22339 16445
rect 22281 16405 22293 16439
rect 22327 16436 22339 16439
rect 22370 16436 22376 16448
rect 22327 16408 22376 16436
rect 22327 16405 22339 16408
rect 22281 16399 22339 16405
rect 22370 16396 22376 16408
rect 22428 16436 22434 16448
rect 23658 16436 23664 16448
rect 22428 16408 23664 16436
rect 22428 16396 22434 16408
rect 23658 16396 23664 16408
rect 23716 16396 23722 16448
rect 24394 16396 24400 16448
rect 24452 16436 24458 16448
rect 24872 16436 24900 16476
rect 25498 16464 25504 16516
rect 25556 16464 25562 16516
rect 24452 16408 24900 16436
rect 25041 16439 25099 16445
rect 24452 16396 24458 16408
rect 25041 16405 25053 16439
rect 25087 16436 25099 16439
rect 25406 16436 25412 16448
rect 25087 16408 25412 16436
rect 25087 16405 25099 16408
rect 25041 16399 25099 16405
rect 25406 16396 25412 16408
rect 25464 16396 25470 16448
rect 25516 16436 25544 16464
rect 25866 16436 25872 16448
rect 25516 16408 25872 16436
rect 25866 16396 25872 16408
rect 25924 16396 25930 16448
rect 26620 16436 26648 16535
rect 26786 16532 26792 16584
rect 26844 16532 26850 16584
rect 26881 16575 26939 16581
rect 26881 16541 26893 16575
rect 26927 16572 26939 16575
rect 26927 16544 27016 16572
rect 26927 16541 26939 16544
rect 26881 16535 26939 16541
rect 26878 16436 26884 16448
rect 26620 16408 26884 16436
rect 26878 16396 26884 16408
rect 26936 16396 26942 16448
rect 26988 16436 27016 16544
rect 28350 16532 28356 16584
rect 28408 16572 28414 16584
rect 28902 16572 28908 16584
rect 28408 16544 28908 16572
rect 28408 16532 28414 16544
rect 28902 16532 28908 16544
rect 28960 16532 28966 16584
rect 28994 16532 29000 16584
rect 29052 16532 29058 16584
rect 29178 16532 29184 16584
rect 29236 16532 29242 16584
rect 29362 16532 29368 16584
rect 29420 16532 29426 16584
rect 29546 16532 29552 16584
rect 29604 16532 29610 16584
rect 29656 16581 29684 16612
rect 29840 16584 29868 16680
rect 30558 16668 30564 16680
rect 30616 16708 30622 16720
rect 31386 16708 31392 16720
rect 30616 16680 31392 16708
rect 30616 16668 30622 16680
rect 31386 16668 31392 16680
rect 31444 16668 31450 16720
rect 34054 16668 34060 16720
rect 34112 16708 34118 16720
rect 34112 16680 35296 16708
rect 34112 16668 34118 16680
rect 35268 16652 35296 16680
rect 30653 16643 30711 16649
rect 30653 16609 30665 16643
rect 30699 16640 30711 16643
rect 31297 16643 31355 16649
rect 31297 16640 31309 16643
rect 30699 16612 31309 16640
rect 30699 16609 30711 16612
rect 30653 16603 30711 16609
rect 31297 16609 31309 16612
rect 31343 16609 31355 16643
rect 31297 16603 31355 16609
rect 33045 16643 33103 16649
rect 33045 16609 33057 16643
rect 33091 16640 33103 16643
rect 33502 16640 33508 16652
rect 33091 16612 33508 16640
rect 33091 16609 33103 16612
rect 33045 16603 33103 16609
rect 29642 16575 29700 16581
rect 29642 16541 29654 16575
rect 29688 16541 29700 16575
rect 29642 16535 29700 16541
rect 29822 16532 29828 16584
rect 29880 16532 29886 16584
rect 30055 16575 30113 16581
rect 30055 16541 30067 16575
rect 30101 16572 30113 16575
rect 30466 16572 30472 16584
rect 30101 16544 30472 16572
rect 30101 16541 30113 16544
rect 30055 16535 30113 16541
rect 30466 16532 30472 16544
rect 30524 16532 30530 16584
rect 29089 16507 29147 16513
rect 29089 16473 29101 16507
rect 29135 16504 29147 16507
rect 29917 16507 29975 16513
rect 29917 16504 29929 16507
rect 29135 16476 29929 16504
rect 29135 16473 29147 16476
rect 29089 16467 29147 16473
rect 29917 16473 29929 16476
rect 29963 16504 29975 16507
rect 30190 16504 30196 16516
rect 29963 16476 30196 16504
rect 29963 16473 29975 16476
rect 29917 16467 29975 16473
rect 30190 16464 30196 16476
rect 30248 16504 30254 16516
rect 30668 16504 30696 16603
rect 33502 16600 33508 16612
rect 33560 16600 33566 16652
rect 34790 16600 34796 16652
rect 34848 16640 34854 16652
rect 34848 16612 35112 16640
rect 34848 16600 34854 16612
rect 35084 16581 35112 16612
rect 35250 16600 35256 16652
rect 35308 16640 35314 16652
rect 35345 16643 35403 16649
rect 35345 16640 35357 16643
rect 35308 16612 35357 16640
rect 35308 16600 35314 16612
rect 35345 16609 35357 16612
rect 35391 16609 35403 16643
rect 35345 16603 35403 16609
rect 35069 16575 35127 16581
rect 35069 16541 35081 16575
rect 35115 16541 35127 16575
rect 35069 16535 35127 16541
rect 35158 16532 35164 16584
rect 35216 16532 35222 16584
rect 35434 16532 35440 16584
rect 35492 16532 35498 16584
rect 35710 16532 35716 16584
rect 35768 16532 35774 16584
rect 35912 16581 35940 16748
rect 37090 16736 37096 16788
rect 37148 16736 37154 16788
rect 37182 16736 37188 16788
rect 37240 16776 37246 16788
rect 38013 16779 38071 16785
rect 37240 16748 37780 16776
rect 37240 16736 37246 16748
rect 36722 16708 36728 16720
rect 36464 16680 36728 16708
rect 35986 16600 35992 16652
rect 36044 16640 36050 16652
rect 36044 16612 36124 16640
rect 36044 16600 36050 16612
rect 36096 16581 36124 16612
rect 35897 16575 35955 16581
rect 35897 16541 35909 16575
rect 35943 16541 35955 16575
rect 35897 16535 35955 16541
rect 36081 16575 36139 16581
rect 36081 16541 36093 16575
rect 36127 16541 36139 16575
rect 36081 16535 36139 16541
rect 31478 16504 31484 16516
rect 30248 16476 30696 16504
rect 31128 16476 31484 16504
rect 30248 16464 30254 16476
rect 28813 16439 28871 16445
rect 28813 16436 28825 16439
rect 26988 16408 28825 16436
rect 28813 16405 28825 16408
rect 28859 16405 28871 16439
rect 28813 16399 28871 16405
rect 29546 16396 29552 16448
rect 29604 16436 29610 16448
rect 30098 16436 30104 16448
rect 29604 16408 30104 16436
rect 29604 16396 29610 16408
rect 30098 16396 30104 16408
rect 30156 16436 30162 16448
rect 30285 16439 30343 16445
rect 30285 16436 30297 16439
rect 30156 16408 30297 16436
rect 30156 16396 30162 16408
rect 30285 16405 30297 16408
rect 30331 16405 30343 16439
rect 30285 16399 30343 16405
rect 30650 16396 30656 16448
rect 30708 16436 30714 16448
rect 31128 16436 31156 16476
rect 31478 16464 31484 16476
rect 31536 16504 31542 16516
rect 31536 16476 31754 16504
rect 32338 16476 32536 16504
rect 31536 16464 31542 16476
rect 30708 16408 31156 16436
rect 30708 16396 30714 16408
rect 31202 16396 31208 16448
rect 31260 16396 31266 16448
rect 31726 16436 31754 16476
rect 32508 16436 32536 16476
rect 32766 16464 32772 16516
rect 32824 16464 32830 16516
rect 35342 16504 35348 16516
rect 34532 16476 35348 16504
rect 34532 16436 34560 16476
rect 35342 16464 35348 16476
rect 35400 16464 35406 16516
rect 35805 16507 35863 16513
rect 35805 16473 35817 16507
rect 35851 16504 35863 16507
rect 35851 16476 35940 16504
rect 35851 16473 35863 16476
rect 35805 16467 35863 16473
rect 31726 16408 34560 16436
rect 34882 16396 34888 16448
rect 34940 16396 34946 16448
rect 35158 16396 35164 16448
rect 35216 16436 35222 16448
rect 35529 16439 35587 16445
rect 35529 16436 35541 16439
rect 35216 16408 35541 16436
rect 35216 16396 35222 16408
rect 35529 16405 35541 16408
rect 35575 16405 35587 16439
rect 35912 16436 35940 16476
rect 35986 16464 35992 16516
rect 36044 16504 36050 16516
rect 36464 16504 36492 16680
rect 36722 16668 36728 16680
rect 36780 16668 36786 16720
rect 36814 16668 36820 16720
rect 36872 16708 36878 16720
rect 37108 16708 37136 16736
rect 37553 16711 37611 16717
rect 37553 16708 37565 16711
rect 36872 16680 37565 16708
rect 36872 16668 36878 16680
rect 37553 16677 37565 16680
rect 37599 16677 37611 16711
rect 37553 16671 37611 16677
rect 36630 16532 36636 16584
rect 36688 16572 36694 16584
rect 37752 16581 37780 16748
rect 38013 16745 38025 16779
rect 38059 16776 38071 16779
rect 38654 16776 38660 16788
rect 38059 16748 38660 16776
rect 38059 16745 38071 16748
rect 38013 16739 38071 16745
rect 38654 16736 38660 16748
rect 38712 16736 38718 16788
rect 39117 16779 39175 16785
rect 39117 16745 39129 16779
rect 39163 16776 39175 16779
rect 39942 16776 39948 16788
rect 39163 16748 39948 16776
rect 39163 16745 39175 16748
rect 39117 16739 39175 16745
rect 39942 16736 39948 16748
rect 40000 16736 40006 16788
rect 41322 16776 41328 16788
rect 40052 16748 41328 16776
rect 38470 16668 38476 16720
rect 38528 16708 38534 16720
rect 39669 16711 39727 16717
rect 39669 16708 39681 16711
rect 38528 16680 39681 16708
rect 38528 16668 38534 16680
rect 39669 16677 39681 16680
rect 39715 16708 39727 16711
rect 40052 16708 40080 16748
rect 41322 16736 41328 16748
rect 41380 16736 41386 16788
rect 43257 16779 43315 16785
rect 43257 16745 43269 16779
rect 43303 16776 43315 16779
rect 43625 16779 43683 16785
rect 43625 16776 43637 16779
rect 43303 16748 43637 16776
rect 43303 16745 43315 16748
rect 43257 16739 43315 16745
rect 43625 16745 43637 16748
rect 43671 16776 43683 16779
rect 44269 16779 44327 16785
rect 44269 16776 44281 16779
rect 43671 16748 44281 16776
rect 43671 16745 43683 16748
rect 43625 16739 43683 16745
rect 44269 16745 44281 16748
rect 44315 16776 44327 16779
rect 45370 16776 45376 16788
rect 44315 16748 45376 16776
rect 44315 16745 44327 16748
rect 44269 16739 44327 16745
rect 45370 16736 45376 16748
rect 45428 16736 45434 16788
rect 45925 16779 45983 16785
rect 45925 16745 45937 16779
rect 45971 16776 45983 16779
rect 46474 16776 46480 16788
rect 45971 16748 46480 16776
rect 45971 16745 45983 16748
rect 45925 16739 45983 16745
rect 46474 16736 46480 16748
rect 46532 16736 46538 16788
rect 47854 16736 47860 16788
rect 47912 16776 47918 16788
rect 48038 16776 48044 16788
rect 47912 16748 48044 16776
rect 47912 16736 47918 16748
rect 48038 16736 48044 16748
rect 48096 16736 48102 16788
rect 48314 16736 48320 16788
rect 48372 16736 48378 16788
rect 48409 16779 48467 16785
rect 48409 16745 48421 16779
rect 48455 16776 48467 16779
rect 48866 16776 48872 16788
rect 48455 16748 48872 16776
rect 48455 16745 48467 16748
rect 48409 16739 48467 16745
rect 48866 16736 48872 16748
rect 48924 16736 48930 16788
rect 49896 16748 51488 16776
rect 39715 16680 40080 16708
rect 39715 16677 39727 16680
rect 39669 16671 39727 16677
rect 40126 16668 40132 16720
rect 40184 16708 40190 16720
rect 40678 16708 40684 16720
rect 40184 16680 40684 16708
rect 40184 16668 40190 16680
rect 40678 16668 40684 16680
rect 40736 16668 40742 16720
rect 40770 16668 40776 16720
rect 40828 16708 40834 16720
rect 41046 16708 41052 16720
rect 40828 16680 41052 16708
rect 40828 16668 40834 16680
rect 41046 16668 41052 16680
rect 41104 16668 41110 16720
rect 41138 16668 41144 16720
rect 41196 16708 41202 16720
rect 41196 16680 41460 16708
rect 41196 16668 41202 16680
rect 40862 16640 40868 16652
rect 38856 16612 39068 16640
rect 36725 16575 36783 16581
rect 36725 16572 36737 16575
rect 36688 16544 36737 16572
rect 36688 16532 36694 16544
rect 36725 16541 36737 16544
rect 36771 16541 36783 16575
rect 36725 16535 36783 16541
rect 37737 16575 37795 16581
rect 37737 16541 37749 16575
rect 37783 16541 37795 16575
rect 37737 16535 37795 16541
rect 37826 16532 37832 16584
rect 37884 16572 37890 16584
rect 38565 16575 38623 16581
rect 38565 16572 38577 16575
rect 37884 16544 38577 16572
rect 37884 16532 37890 16544
rect 38565 16541 38577 16544
rect 38611 16541 38623 16575
rect 38856 16572 38884 16612
rect 38565 16535 38623 16541
rect 38672 16544 38884 16572
rect 36044 16476 36492 16504
rect 36044 16464 36050 16476
rect 36538 16464 36544 16516
rect 36596 16504 36602 16516
rect 36596 16476 36952 16504
rect 36596 16464 36602 16476
rect 36078 16436 36084 16448
rect 35912 16408 36084 16436
rect 35529 16399 35587 16405
rect 36078 16396 36084 16408
rect 36136 16396 36142 16448
rect 36449 16439 36507 16445
rect 36449 16405 36461 16439
rect 36495 16436 36507 16439
rect 36722 16436 36728 16448
rect 36495 16408 36728 16436
rect 36495 16405 36507 16408
rect 36449 16399 36507 16405
rect 36722 16396 36728 16408
rect 36780 16396 36786 16448
rect 36924 16445 36952 16476
rect 37274 16464 37280 16516
rect 37332 16464 37338 16516
rect 37921 16507 37979 16513
rect 37921 16473 37933 16507
rect 37967 16473 37979 16507
rect 37921 16467 37979 16473
rect 36909 16439 36967 16445
rect 36909 16405 36921 16439
rect 36955 16436 36967 16439
rect 37458 16436 37464 16448
rect 36955 16408 37464 16436
rect 36955 16405 36967 16408
rect 36909 16399 36967 16405
rect 37458 16396 37464 16408
rect 37516 16396 37522 16448
rect 37936 16436 37964 16467
rect 38286 16464 38292 16516
rect 38344 16464 38350 16516
rect 38378 16464 38384 16516
rect 38436 16504 38442 16516
rect 38672 16504 38700 16544
rect 38930 16532 38936 16584
rect 38988 16532 38994 16584
rect 39040 16572 39068 16612
rect 39961 16612 40172 16640
rect 39301 16575 39359 16581
rect 39301 16572 39313 16575
rect 39040 16544 39313 16572
rect 39301 16541 39313 16544
rect 39347 16541 39359 16575
rect 39301 16535 39359 16541
rect 38436 16476 38700 16504
rect 38436 16464 38442 16476
rect 38746 16464 38752 16516
rect 38804 16464 38810 16516
rect 38838 16464 38844 16516
rect 38896 16464 38902 16516
rect 39961 16504 39989 16612
rect 40034 16532 40040 16584
rect 40092 16532 40098 16584
rect 40144 16572 40172 16612
rect 40696 16612 40868 16640
rect 40696 16581 40724 16612
rect 40862 16600 40868 16612
rect 40920 16600 40926 16652
rect 40954 16600 40960 16652
rect 41012 16640 41018 16652
rect 41322 16640 41328 16652
rect 41012 16612 41328 16640
rect 41012 16600 41018 16612
rect 41322 16600 41328 16612
rect 41380 16600 41386 16652
rect 41432 16640 41460 16680
rect 41506 16668 41512 16720
rect 41564 16708 41570 16720
rect 43990 16708 43996 16720
rect 41564 16680 43996 16708
rect 41564 16668 41570 16680
rect 43990 16668 43996 16680
rect 44048 16668 44054 16720
rect 46842 16668 46848 16720
rect 46900 16708 46906 16720
rect 48498 16708 48504 16720
rect 46900 16680 48504 16708
rect 46900 16668 46906 16680
rect 48498 16668 48504 16680
rect 48556 16708 48562 16720
rect 49896 16708 49924 16748
rect 48556 16680 49924 16708
rect 49973 16711 50031 16717
rect 48556 16668 48562 16680
rect 49973 16677 49985 16711
rect 50019 16708 50031 16711
rect 50062 16708 50068 16720
rect 50019 16680 50068 16708
rect 50019 16677 50031 16680
rect 49973 16671 50031 16677
rect 50062 16668 50068 16680
rect 50120 16668 50126 16720
rect 51350 16708 51356 16720
rect 51046 16680 51356 16708
rect 45649 16643 45707 16649
rect 45649 16640 45661 16643
rect 41432 16612 43852 16640
rect 40405 16575 40463 16581
rect 40405 16572 40417 16575
rect 40144 16544 40417 16572
rect 40405 16541 40417 16544
rect 40451 16541 40463 16575
rect 40405 16535 40463 16541
rect 40681 16575 40739 16581
rect 40681 16541 40693 16575
rect 40727 16541 40739 16575
rect 40681 16535 40739 16541
rect 40770 16532 40776 16584
rect 40828 16532 40834 16584
rect 41049 16575 41107 16581
rect 41049 16541 41061 16575
rect 41095 16572 41107 16575
rect 41417 16575 41475 16581
rect 41417 16572 41429 16575
rect 41095 16544 41429 16572
rect 41095 16541 41107 16544
rect 41049 16535 41107 16541
rect 41417 16541 41429 16544
rect 41463 16541 41475 16575
rect 41417 16535 41475 16541
rect 41782 16532 41788 16584
rect 41840 16572 41846 16584
rect 41969 16575 42027 16581
rect 41969 16572 41981 16575
rect 41840 16544 41981 16572
rect 41840 16532 41846 16544
rect 41969 16541 41981 16544
rect 42015 16541 42027 16575
rect 41969 16535 42027 16541
rect 42794 16532 42800 16584
rect 42852 16532 42858 16584
rect 42978 16532 42984 16584
rect 43036 16532 43042 16584
rect 43070 16532 43076 16584
rect 43128 16532 43134 16584
rect 43162 16532 43168 16584
rect 43220 16572 43226 16584
rect 43303 16575 43361 16581
rect 43303 16572 43315 16575
rect 43220 16544 43315 16572
rect 43220 16532 43226 16544
rect 43303 16541 43315 16544
rect 43349 16541 43361 16575
rect 43303 16535 43361 16541
rect 39316 16476 39989 16504
rect 38470 16436 38476 16448
rect 37936 16408 38476 16436
rect 38470 16396 38476 16408
rect 38528 16396 38534 16448
rect 38654 16396 38660 16448
rect 38712 16436 38718 16448
rect 39316 16436 39344 16476
rect 40126 16464 40132 16516
rect 40184 16464 40190 16516
rect 40221 16507 40279 16513
rect 40221 16473 40233 16507
rect 40267 16504 40279 16507
rect 41874 16504 41880 16516
rect 40267 16476 41880 16504
rect 40267 16473 40279 16476
rect 40221 16467 40279 16473
rect 41874 16464 41880 16476
rect 41932 16464 41938 16516
rect 43533 16507 43591 16513
rect 43533 16473 43545 16507
rect 43579 16473 43591 16507
rect 43824 16504 43852 16612
rect 44284 16612 45661 16640
rect 43898 16532 43904 16584
rect 43956 16572 43962 16584
rect 43993 16575 44051 16581
rect 43993 16572 44005 16575
rect 43956 16544 44005 16572
rect 43956 16532 43962 16544
rect 43993 16541 44005 16544
rect 44039 16541 44051 16575
rect 43993 16535 44051 16541
rect 44085 16575 44143 16581
rect 44085 16541 44097 16575
rect 44131 16572 44143 16575
rect 44174 16572 44180 16584
rect 44131 16544 44180 16572
rect 44131 16541 44143 16544
rect 44085 16535 44143 16541
rect 44174 16532 44180 16544
rect 44232 16532 44238 16584
rect 44284 16504 44312 16612
rect 45649 16609 45661 16612
rect 45695 16640 45707 16643
rect 46290 16640 46296 16652
rect 45695 16612 46296 16640
rect 45695 16609 45707 16612
rect 45649 16603 45707 16609
rect 46290 16600 46296 16612
rect 46348 16600 46354 16652
rect 47397 16643 47455 16649
rect 47397 16609 47409 16643
rect 47443 16640 47455 16643
rect 47946 16640 47952 16652
rect 47443 16612 47952 16640
rect 47443 16609 47455 16612
rect 47397 16603 47455 16609
rect 44361 16575 44419 16581
rect 44361 16541 44373 16575
rect 44407 16572 44419 16575
rect 45278 16572 45284 16584
rect 44407 16544 45284 16572
rect 44407 16541 44419 16544
rect 44361 16535 44419 16541
rect 45278 16532 45284 16544
rect 45336 16532 45342 16584
rect 46385 16575 46443 16581
rect 46385 16541 46397 16575
rect 46431 16572 46443 16575
rect 47412 16572 47440 16603
rect 47946 16600 47952 16612
rect 48004 16600 48010 16652
rect 48038 16600 48044 16652
rect 48096 16640 48102 16652
rect 51046 16640 51074 16680
rect 51350 16668 51356 16680
rect 51408 16668 51414 16720
rect 48096 16612 51074 16640
rect 51460 16640 51488 16748
rect 53834 16736 53840 16788
rect 53892 16776 53898 16788
rect 54846 16776 54852 16788
rect 53892 16748 54852 16776
rect 53892 16736 53898 16748
rect 54846 16736 54852 16748
rect 54904 16736 54910 16788
rect 56594 16736 56600 16788
rect 56652 16776 56658 16788
rect 56873 16779 56931 16785
rect 56873 16776 56885 16779
rect 56652 16748 56885 16776
rect 56652 16736 56658 16748
rect 56873 16745 56885 16748
rect 56919 16745 56931 16779
rect 56873 16739 56931 16745
rect 53558 16668 53564 16720
rect 53616 16708 53622 16720
rect 53616 16680 56456 16708
rect 53616 16668 53622 16680
rect 55306 16640 55312 16652
rect 51460 16612 55312 16640
rect 48096 16600 48102 16612
rect 55306 16600 55312 16612
rect 55364 16600 55370 16652
rect 55766 16600 55772 16652
rect 55824 16640 55830 16652
rect 55824 16612 56364 16640
rect 55824 16600 55830 16612
rect 46431 16544 47440 16572
rect 46431 16541 46443 16544
rect 46385 16535 46443 16541
rect 47486 16532 47492 16584
rect 47544 16572 47550 16584
rect 47673 16575 47731 16581
rect 47673 16572 47685 16575
rect 47544 16544 47685 16572
rect 47544 16532 47550 16544
rect 47673 16541 47685 16544
rect 47719 16541 47731 16575
rect 47673 16535 47731 16541
rect 47762 16532 47768 16584
rect 47820 16572 47826 16584
rect 48157 16575 48215 16581
rect 48157 16572 48169 16575
rect 47820 16544 47865 16572
rect 47820 16532 47826 16544
rect 48153 16541 48169 16572
rect 48203 16541 48215 16575
rect 48153 16535 48215 16541
rect 43824 16476 44312 16504
rect 46569 16507 46627 16513
rect 43533 16467 43591 16473
rect 46569 16473 46581 16507
rect 46615 16504 46627 16507
rect 46842 16504 46848 16516
rect 46615 16476 46848 16504
rect 46615 16473 46627 16476
rect 46569 16467 46627 16473
rect 38712 16408 39344 16436
rect 38712 16396 38718 16408
rect 39390 16396 39396 16448
rect 39448 16396 39454 16448
rect 39666 16396 39672 16448
rect 39724 16436 39730 16448
rect 39853 16439 39911 16445
rect 39853 16436 39865 16439
rect 39724 16408 39865 16436
rect 39724 16396 39730 16408
rect 39853 16405 39865 16408
rect 39899 16405 39911 16439
rect 39853 16399 39911 16405
rect 40310 16396 40316 16448
rect 40368 16436 40374 16448
rect 40497 16439 40555 16445
rect 40497 16436 40509 16439
rect 40368 16408 40509 16436
rect 40368 16396 40374 16408
rect 40497 16405 40509 16408
rect 40543 16405 40555 16439
rect 40497 16399 40555 16405
rect 41138 16396 41144 16448
rect 41196 16396 41202 16448
rect 42058 16396 42064 16448
rect 42116 16436 42122 16448
rect 42610 16436 42616 16448
rect 42116 16408 42616 16436
rect 42116 16396 42122 16408
rect 42610 16396 42616 16408
rect 42668 16436 42674 16448
rect 43548 16436 43576 16467
rect 46842 16464 46848 16476
rect 46900 16464 46906 16516
rect 47578 16464 47584 16516
rect 47636 16504 47642 16516
rect 47949 16507 48007 16513
rect 47949 16504 47961 16507
rect 47636 16476 47961 16504
rect 47636 16464 47642 16476
rect 47949 16473 47961 16476
rect 47995 16473 48007 16507
rect 47949 16467 48007 16473
rect 48038 16464 48044 16516
rect 48096 16464 48102 16516
rect 48153 16504 48181 16535
rect 48590 16532 48596 16584
rect 48648 16572 48654 16584
rect 48866 16572 48872 16584
rect 48648 16544 48872 16572
rect 48648 16532 48654 16544
rect 48866 16532 48872 16544
rect 48924 16532 48930 16584
rect 48961 16575 49019 16581
rect 48961 16541 48973 16575
rect 49007 16572 49019 16575
rect 49326 16572 49332 16584
rect 49007 16544 49332 16572
rect 49007 16541 49019 16544
rect 48961 16535 49019 16541
rect 49326 16532 49332 16544
rect 49384 16532 49390 16584
rect 49418 16532 49424 16584
rect 49476 16532 49482 16584
rect 49602 16532 49608 16584
rect 49660 16532 49666 16584
rect 49789 16575 49847 16581
rect 49789 16541 49801 16575
rect 49835 16572 49847 16575
rect 54110 16572 54116 16584
rect 49835 16544 54116 16572
rect 49835 16541 49847 16544
rect 49789 16535 49847 16541
rect 54110 16532 54116 16544
rect 54168 16532 54174 16584
rect 56336 16581 56364 16612
rect 56045 16575 56103 16581
rect 56045 16572 56057 16575
rect 54220 16544 56057 16572
rect 48153 16476 48268 16504
rect 48240 16448 48268 16476
rect 48314 16464 48320 16516
rect 48372 16504 48378 16516
rect 48685 16507 48743 16513
rect 48685 16504 48697 16507
rect 48372 16476 48697 16504
rect 48372 16464 48378 16476
rect 48685 16473 48697 16476
rect 48731 16473 48743 16507
rect 48685 16467 48743 16473
rect 48777 16507 48835 16513
rect 48777 16473 48789 16507
rect 48823 16504 48835 16507
rect 49050 16504 49056 16516
rect 48823 16476 49056 16504
rect 48823 16473 48835 16476
rect 48777 16467 48835 16473
rect 49050 16464 49056 16476
rect 49108 16464 49114 16516
rect 49142 16464 49148 16516
rect 49200 16504 49206 16516
rect 49513 16507 49571 16513
rect 49513 16504 49525 16507
rect 49200 16476 49525 16504
rect 49200 16464 49206 16476
rect 49513 16473 49525 16476
rect 49559 16473 49571 16507
rect 50338 16504 50344 16516
rect 49513 16467 49571 16473
rect 49804 16476 50344 16504
rect 42668 16408 43576 16436
rect 42668 16396 42674 16408
rect 43806 16396 43812 16448
rect 43864 16396 43870 16448
rect 48222 16396 48228 16448
rect 48280 16436 48286 16448
rect 48590 16436 48596 16448
rect 48280 16408 48596 16436
rect 48280 16396 48286 16408
rect 48590 16396 48596 16408
rect 48648 16396 48654 16448
rect 49237 16439 49295 16445
rect 49237 16405 49249 16439
rect 49283 16436 49295 16439
rect 49804 16436 49832 16476
rect 50338 16464 50344 16476
rect 50396 16464 50402 16516
rect 53926 16464 53932 16516
rect 53984 16504 53990 16516
rect 54220 16513 54248 16544
rect 56045 16541 56057 16544
rect 56091 16541 56103 16575
rect 56045 16535 56103 16541
rect 56321 16575 56379 16581
rect 56321 16541 56333 16575
rect 56367 16541 56379 16575
rect 56428 16572 56456 16680
rect 56689 16575 56747 16581
rect 56689 16572 56701 16575
rect 56428 16544 56701 16572
rect 56321 16535 56379 16541
rect 56689 16541 56701 16544
rect 56735 16572 56747 16575
rect 57149 16575 57207 16581
rect 57149 16572 57161 16575
rect 56735 16544 57161 16572
rect 56735 16541 56747 16544
rect 56689 16535 56747 16541
rect 57149 16541 57161 16544
rect 57195 16541 57207 16575
rect 57149 16535 57207 16541
rect 57514 16532 57520 16584
rect 57572 16532 57578 16584
rect 54205 16507 54263 16513
rect 54205 16504 54217 16507
rect 53984 16476 54217 16504
rect 53984 16464 53990 16476
rect 54205 16473 54217 16476
rect 54251 16473 54263 16507
rect 54205 16467 54263 16473
rect 55306 16464 55312 16516
rect 55364 16464 55370 16516
rect 55950 16464 55956 16516
rect 56008 16504 56014 16516
rect 56505 16507 56563 16513
rect 56505 16504 56517 16507
rect 56008 16476 56517 16504
rect 56008 16464 56014 16476
rect 56505 16473 56517 16476
rect 56551 16473 56563 16507
rect 56505 16467 56563 16473
rect 56597 16507 56655 16513
rect 56597 16473 56609 16507
rect 56643 16473 56655 16507
rect 56597 16467 56655 16473
rect 49283 16408 49832 16436
rect 49283 16405 49295 16408
rect 49237 16399 49295 16405
rect 54110 16396 54116 16448
rect 54168 16436 54174 16448
rect 56612 16436 56640 16467
rect 57238 16464 57244 16516
rect 57296 16464 57302 16516
rect 57330 16464 57336 16516
rect 57388 16464 57394 16516
rect 54168 16408 56640 16436
rect 54168 16396 54174 16408
rect 56962 16396 56968 16448
rect 57020 16396 57026 16448
rect 1104 16346 58880 16368
rect 1104 16294 4874 16346
rect 4926 16294 4938 16346
rect 4990 16294 5002 16346
rect 5054 16294 5066 16346
rect 5118 16294 5130 16346
rect 5182 16294 35594 16346
rect 35646 16294 35658 16346
rect 35710 16294 35722 16346
rect 35774 16294 35786 16346
rect 35838 16294 35850 16346
rect 35902 16294 58880 16346
rect 1104 16272 58880 16294
rect 19518 16232 19524 16244
rect 19260 16204 19524 16232
rect 19260 16105 19288 16204
rect 19518 16192 19524 16204
rect 19576 16192 19582 16244
rect 19794 16192 19800 16244
rect 19852 16192 19858 16244
rect 19889 16235 19947 16241
rect 19889 16201 19901 16235
rect 19935 16232 19947 16235
rect 20254 16232 20260 16244
rect 19935 16204 20260 16232
rect 19935 16201 19947 16204
rect 19889 16195 19947 16201
rect 20254 16192 20260 16204
rect 20312 16192 20318 16244
rect 20806 16192 20812 16244
rect 20864 16232 20870 16244
rect 21177 16235 21235 16241
rect 21177 16232 21189 16235
rect 20864 16204 21189 16232
rect 20864 16192 20870 16204
rect 21177 16201 21189 16204
rect 21223 16201 21235 16235
rect 21177 16195 21235 16201
rect 21634 16192 21640 16244
rect 21692 16232 21698 16244
rect 22370 16232 22376 16244
rect 21692 16204 22376 16232
rect 21692 16192 21698 16204
rect 22370 16192 22376 16204
rect 22428 16192 22434 16244
rect 23109 16235 23167 16241
rect 23109 16201 23121 16235
rect 23155 16232 23167 16235
rect 23198 16232 23204 16244
rect 23155 16204 23204 16232
rect 23155 16201 23167 16204
rect 23109 16195 23167 16201
rect 23198 16192 23204 16204
rect 23256 16192 23262 16244
rect 24946 16192 24952 16244
rect 25004 16192 25010 16244
rect 25130 16192 25136 16244
rect 25188 16232 25194 16244
rect 25317 16235 25375 16241
rect 25317 16232 25329 16235
rect 25188 16204 25329 16232
rect 25188 16192 25194 16204
rect 25317 16201 25329 16204
rect 25363 16201 25375 16235
rect 27893 16235 27951 16241
rect 27893 16232 27905 16235
rect 25317 16195 25375 16201
rect 27092 16204 27905 16232
rect 19812 16164 19840 16192
rect 22097 16167 22155 16173
rect 19444 16136 19840 16164
rect 19904 16136 21956 16164
rect 19444 16105 19472 16136
rect 19245 16099 19303 16105
rect 19245 16065 19257 16099
rect 19291 16065 19303 16099
rect 19245 16059 19303 16065
rect 19393 16099 19472 16105
rect 19393 16065 19405 16099
rect 19439 16068 19472 16099
rect 19439 16065 19451 16068
rect 19393 16059 19451 16065
rect 19518 16056 19524 16108
rect 19576 16056 19582 16108
rect 19613 16099 19671 16105
rect 19613 16065 19625 16099
rect 19659 16065 19671 16099
rect 19613 16059 19671 16065
rect 18966 15988 18972 16040
rect 19024 16028 19030 16040
rect 19628 16028 19656 16059
rect 19702 16056 19708 16108
rect 19760 16105 19766 16108
rect 19760 16099 19809 16105
rect 19760 16065 19763 16099
rect 19797 16096 19809 16099
rect 19904 16096 19932 16136
rect 19797 16068 19932 16096
rect 21361 16099 21419 16105
rect 19797 16065 19809 16068
rect 19760 16059 19809 16065
rect 21361 16065 21373 16099
rect 21407 16096 21419 16099
rect 21928 16096 21956 16136
rect 22097 16133 22109 16167
rect 22143 16164 22155 16167
rect 23014 16164 23020 16176
rect 22143 16136 23020 16164
rect 22143 16133 22155 16136
rect 22097 16127 22155 16133
rect 23014 16124 23020 16136
rect 23072 16124 23078 16176
rect 23385 16167 23443 16173
rect 23385 16133 23397 16167
rect 23431 16164 23443 16167
rect 24670 16164 24676 16176
rect 23431 16136 24676 16164
rect 23431 16133 23443 16136
rect 23385 16127 23443 16133
rect 24670 16124 24676 16136
rect 24728 16124 24734 16176
rect 27092 16164 27120 16204
rect 27893 16201 27905 16204
rect 27939 16201 27951 16235
rect 27893 16195 27951 16201
rect 29178 16192 29184 16244
rect 29236 16192 29242 16244
rect 30374 16232 30380 16244
rect 29380 16204 30380 16232
rect 25332 16136 27120 16164
rect 22000 16099 22058 16105
rect 22000 16096 22012 16099
rect 21407 16068 21864 16096
rect 21928 16068 22012 16096
rect 21407 16065 21419 16068
rect 21361 16059 21419 16065
rect 19760 16056 19766 16059
rect 20162 16028 20168 16040
rect 19024 16000 20168 16028
rect 19024 15988 19030 16000
rect 19996 15892 20024 16000
rect 20162 15988 20168 16000
rect 20220 15988 20226 16040
rect 21634 15988 21640 16040
rect 21692 15988 21698 16040
rect 20070 15920 20076 15972
rect 20128 15960 20134 15972
rect 21542 15960 21548 15972
rect 20128 15932 21548 15960
rect 20128 15920 20134 15932
rect 21542 15920 21548 15932
rect 21600 15920 21606 15972
rect 21836 15969 21864 16068
rect 22000 16065 22012 16068
rect 22046 16065 22058 16099
rect 22000 16059 22058 16065
rect 22020 16028 22048 16059
rect 22186 16056 22192 16108
rect 22244 16056 22250 16108
rect 22278 16056 22284 16108
rect 22336 16105 22342 16108
rect 22336 16099 22375 16105
rect 22363 16065 22375 16099
rect 22336 16059 22375 16065
rect 22336 16056 22342 16059
rect 22462 16056 22468 16108
rect 22520 16056 22526 16108
rect 23290 16105 23296 16108
rect 23288 16096 23296 16105
rect 22572 16068 23296 16096
rect 22572 16028 22600 16068
rect 23288 16059 23296 16068
rect 23290 16056 23296 16059
rect 23348 16056 23354 16108
rect 23474 16056 23480 16108
rect 23532 16056 23538 16108
rect 23658 16096 23664 16108
rect 23619 16068 23664 16096
rect 23658 16056 23664 16068
rect 23716 16056 23722 16108
rect 23753 16099 23811 16105
rect 23753 16065 23765 16099
rect 23799 16065 23811 16099
rect 23753 16059 23811 16065
rect 22020 16000 22600 16028
rect 23768 15972 23796 16059
rect 23842 16056 23848 16108
rect 23900 16096 23906 16108
rect 24397 16099 24455 16105
rect 24397 16096 24409 16099
rect 23900 16068 24409 16096
rect 23900 16056 23906 16068
rect 24397 16065 24409 16068
rect 24443 16065 24455 16099
rect 24397 16059 24455 16065
rect 24581 16099 24639 16105
rect 24581 16065 24593 16099
rect 24627 16065 24639 16099
rect 24581 16059 24639 16065
rect 24596 16028 24624 16059
rect 24762 16056 24768 16108
rect 24820 16056 24826 16108
rect 25038 16056 25044 16108
rect 25096 16096 25102 16108
rect 25225 16099 25283 16105
rect 25225 16096 25237 16099
rect 25096 16068 25237 16096
rect 25096 16056 25102 16068
rect 25225 16065 25237 16068
rect 25271 16065 25283 16099
rect 25225 16059 25283 16065
rect 25130 16028 25136 16040
rect 24596 16000 25136 16028
rect 25130 15988 25136 16000
rect 25188 15988 25194 16040
rect 21821 15963 21879 15969
rect 21821 15929 21833 15963
rect 21867 15929 21879 15963
rect 21821 15923 21879 15929
rect 22462 15920 22468 15972
rect 22520 15960 22526 15972
rect 22830 15960 22836 15972
rect 22520 15932 22836 15960
rect 22520 15920 22526 15932
rect 22830 15920 22836 15932
rect 22888 15960 22894 15972
rect 23750 15960 23756 15972
rect 22888 15932 23756 15960
rect 22888 15920 22894 15932
rect 23750 15920 23756 15932
rect 23808 15960 23814 15972
rect 25332 15960 25360 16136
rect 25866 16056 25872 16108
rect 25924 16096 25930 16108
rect 26237 16099 26295 16105
rect 26237 16096 26249 16099
rect 25924 16068 26249 16096
rect 25924 16056 25930 16068
rect 26237 16065 26249 16068
rect 26283 16065 26295 16099
rect 26237 16059 26295 16065
rect 26418 16056 26424 16108
rect 26476 16056 26482 16108
rect 27092 16105 27120 16136
rect 27338 16124 27344 16176
rect 27396 16124 27402 16176
rect 27433 16167 27491 16173
rect 27433 16133 27445 16167
rect 27479 16164 27491 16167
rect 29270 16164 29276 16176
rect 27479 16136 29276 16164
rect 27479 16133 27491 16136
rect 27433 16127 27491 16133
rect 29270 16124 29276 16136
rect 29328 16124 29334 16176
rect 26513 16099 26571 16105
rect 26513 16065 26525 16099
rect 26559 16065 26571 16099
rect 26513 16059 26571 16065
rect 26605 16099 26663 16105
rect 26605 16065 26617 16099
rect 26651 16096 26663 16099
rect 27065 16099 27123 16105
rect 26651 16068 26740 16096
rect 26651 16065 26663 16068
rect 26605 16059 26663 16065
rect 26528 15972 26556 16059
rect 26712 16040 26740 16068
rect 27065 16065 27077 16099
rect 27111 16065 27123 16099
rect 27065 16059 27123 16065
rect 27158 16099 27216 16105
rect 27158 16065 27170 16099
rect 27204 16065 27216 16099
rect 27158 16059 27216 16065
rect 26694 15988 26700 16040
rect 26752 15988 26758 16040
rect 26878 15988 26884 16040
rect 26936 16028 26942 16040
rect 27173 16028 27201 16059
rect 27522 16056 27528 16108
rect 27580 16105 27586 16108
rect 29380 16105 29408 16204
rect 30374 16192 30380 16204
rect 30432 16192 30438 16244
rect 31110 16192 31116 16244
rect 31168 16192 31174 16244
rect 31665 16235 31723 16241
rect 31665 16201 31677 16235
rect 31711 16232 31723 16235
rect 32766 16232 32772 16244
rect 31711 16204 32772 16232
rect 31711 16201 31723 16204
rect 31665 16195 31723 16201
rect 32766 16192 32772 16204
rect 32824 16192 32830 16244
rect 35250 16192 35256 16244
rect 35308 16232 35314 16244
rect 35802 16232 35808 16244
rect 35308 16204 35808 16232
rect 35308 16192 35314 16204
rect 35802 16192 35808 16204
rect 35860 16192 35866 16244
rect 36170 16232 36176 16244
rect 35912 16204 36176 16232
rect 29638 16124 29644 16176
rect 29696 16124 29702 16176
rect 30650 16124 30656 16176
rect 30708 16124 30714 16176
rect 33229 16167 33287 16173
rect 33229 16133 33241 16167
rect 33275 16164 33287 16167
rect 33502 16164 33508 16176
rect 33275 16136 33508 16164
rect 33275 16133 33287 16136
rect 33229 16127 33287 16133
rect 33502 16124 33508 16136
rect 33560 16164 33566 16176
rect 35342 16164 35348 16176
rect 33560 16136 33640 16164
rect 35098 16136 35348 16164
rect 33560 16124 33566 16136
rect 27580 16096 27588 16105
rect 28077 16099 28135 16105
rect 27580 16068 27625 16096
rect 27580 16059 27588 16068
rect 28077 16065 28089 16099
rect 28123 16065 28135 16099
rect 28077 16059 28135 16065
rect 29365 16099 29423 16105
rect 29365 16065 29377 16099
rect 29411 16065 29423 16099
rect 29365 16059 29423 16065
rect 27580 16056 27586 16059
rect 28092 16028 28120 16059
rect 31202 16056 31208 16108
rect 31260 16056 31266 16108
rect 31481 16099 31539 16105
rect 31481 16065 31493 16099
rect 31527 16096 31539 16099
rect 31754 16096 31760 16108
rect 31527 16068 31760 16096
rect 31527 16065 31539 16068
rect 31481 16059 31539 16065
rect 31754 16056 31760 16068
rect 31812 16056 31818 16108
rect 33612 16105 33640 16136
rect 35342 16124 35348 16136
rect 35400 16124 35406 16176
rect 35912 16105 35940 16204
rect 36170 16192 36176 16204
rect 36228 16192 36234 16244
rect 36449 16235 36507 16241
rect 36449 16201 36461 16235
rect 36495 16201 36507 16235
rect 38654 16232 38660 16244
rect 36449 16195 36507 16201
rect 36556 16204 38660 16232
rect 36464 16164 36492 16195
rect 36004 16136 36492 16164
rect 36004 16105 36032 16136
rect 36556 16108 36584 16204
rect 38654 16192 38660 16204
rect 38712 16192 38718 16244
rect 38930 16192 38936 16244
rect 38988 16232 38994 16244
rect 38988 16204 39712 16232
rect 38988 16192 38994 16204
rect 36725 16167 36783 16173
rect 36725 16133 36737 16167
rect 36771 16164 36783 16167
rect 39022 16164 39028 16176
rect 36771 16136 39028 16164
rect 36771 16133 36783 16136
rect 36725 16127 36783 16133
rect 39022 16124 39028 16136
rect 39080 16164 39086 16176
rect 39080 16136 39344 16164
rect 39080 16124 39086 16136
rect 32401 16099 32459 16105
rect 32401 16096 32413 16099
rect 32232 16068 32413 16096
rect 28169 16031 28227 16037
rect 28169 16028 28181 16031
rect 26936 16000 27201 16028
rect 27632 16000 28181 16028
rect 26936 15988 26942 16000
rect 23808 15932 25360 15960
rect 23808 15920 23814 15932
rect 26510 15920 26516 15972
rect 26568 15920 26574 15972
rect 26786 15920 26792 15972
rect 26844 15920 26850 15972
rect 24578 15892 24584 15904
rect 19996 15864 24584 15892
rect 24578 15852 24584 15864
rect 24636 15852 24642 15904
rect 24762 15852 24768 15904
rect 24820 15892 24826 15904
rect 25501 15895 25559 15901
rect 25501 15892 25513 15895
rect 24820 15864 25513 15892
rect 24820 15852 24826 15864
rect 25501 15861 25513 15864
rect 25547 15892 25559 15895
rect 26050 15892 26056 15904
rect 25547 15864 26056 15892
rect 25547 15861 25559 15864
rect 25501 15855 25559 15861
rect 26050 15852 26056 15864
rect 26108 15852 26114 15904
rect 26142 15852 26148 15904
rect 26200 15892 26206 15904
rect 27632 15892 27660 16000
rect 28169 15997 28181 16000
rect 28215 15997 28227 16031
rect 28169 15991 28227 15997
rect 32232 15969 32260 16068
rect 32401 16065 32413 16068
rect 32447 16065 32459 16099
rect 32401 16059 32459 16065
rect 33597 16099 33655 16105
rect 33597 16065 33609 16099
rect 33643 16065 33655 16099
rect 33597 16059 33655 16065
rect 35897 16099 35955 16105
rect 35897 16065 35909 16099
rect 35943 16065 35955 16099
rect 35897 16059 35955 16065
rect 35989 16099 36047 16105
rect 35989 16065 36001 16099
rect 36035 16065 36047 16099
rect 35989 16059 36047 16065
rect 36078 16056 36084 16108
rect 36136 16096 36142 16108
rect 36265 16099 36323 16105
rect 36265 16096 36277 16099
rect 36136 16068 36277 16096
rect 36136 16056 36142 16068
rect 36265 16065 36277 16068
rect 36311 16096 36323 16099
rect 36538 16096 36544 16108
rect 36311 16068 36544 16096
rect 36311 16065 36323 16068
rect 36265 16059 36323 16065
rect 36538 16056 36544 16068
rect 36596 16056 36602 16108
rect 36633 16099 36691 16105
rect 36633 16065 36645 16099
rect 36679 16065 36691 16099
rect 36633 16059 36691 16065
rect 33873 16031 33931 16037
rect 33873 15997 33885 16031
rect 33919 16028 33931 16031
rect 34882 16028 34888 16040
rect 33919 16000 34888 16028
rect 33919 15997 33931 16000
rect 33873 15991 33931 15997
rect 34882 15988 34888 16000
rect 34940 15988 34946 16040
rect 35345 16031 35403 16037
rect 35345 15997 35357 16031
rect 35391 16028 35403 16031
rect 35434 16028 35440 16040
rect 35391 16000 35440 16028
rect 35391 15997 35403 16000
rect 35345 15991 35403 15997
rect 35434 15988 35440 16000
rect 35492 15988 35498 16040
rect 36648 16028 36676 16059
rect 36814 16056 36820 16108
rect 36872 16056 36878 16108
rect 36998 16056 37004 16108
rect 37056 16096 37062 16108
rect 37826 16096 37832 16108
rect 37056 16068 37832 16096
rect 37056 16056 37062 16068
rect 37826 16056 37832 16068
rect 37884 16056 37890 16108
rect 37921 16099 37979 16105
rect 37921 16065 37933 16099
rect 37967 16065 37979 16099
rect 37921 16059 37979 16065
rect 37369 16031 37427 16037
rect 36648 16000 37044 16028
rect 32217 15963 32275 15969
rect 32217 15960 32229 15963
rect 30668 15932 32229 15960
rect 26200 15864 27660 15892
rect 27709 15895 27767 15901
rect 26200 15852 26206 15864
rect 27709 15861 27721 15895
rect 27755 15892 27767 15895
rect 27890 15892 27896 15904
rect 27755 15864 27896 15892
rect 27755 15861 27767 15864
rect 27709 15855 27767 15861
rect 27890 15852 27896 15864
rect 27948 15852 27954 15904
rect 27982 15852 27988 15904
rect 28040 15892 28046 15904
rect 29730 15892 29736 15904
rect 28040 15864 29736 15892
rect 28040 15852 28046 15864
rect 29730 15852 29736 15864
rect 29788 15892 29794 15904
rect 30668 15892 30696 15932
rect 32217 15929 32229 15932
rect 32263 15929 32275 15963
rect 32217 15923 32275 15929
rect 35986 15920 35992 15972
rect 36044 15960 36050 15972
rect 36648 15960 36676 16000
rect 37016 15972 37044 16000
rect 37369 15997 37381 16031
rect 37415 16028 37427 16031
rect 37458 16028 37464 16040
rect 37415 16000 37464 16028
rect 37415 15997 37427 16000
rect 37369 15991 37427 15997
rect 37458 15988 37464 16000
rect 37516 15988 37522 16040
rect 36044 15932 36676 15960
rect 36044 15920 36050 15932
rect 36998 15920 37004 15972
rect 37056 15920 37062 15972
rect 37936 15960 37964 16059
rect 38194 16056 38200 16108
rect 38252 16096 38258 16108
rect 38289 16099 38347 16105
rect 38289 16096 38301 16099
rect 38252 16068 38301 16096
rect 38252 16056 38258 16068
rect 38289 16065 38301 16068
rect 38335 16065 38347 16099
rect 38289 16059 38347 16065
rect 38381 16099 38439 16105
rect 38381 16065 38393 16099
rect 38427 16065 38439 16099
rect 38381 16059 38439 16065
rect 38473 16099 38531 16105
rect 38473 16065 38485 16099
rect 38519 16096 38531 16099
rect 38562 16096 38568 16108
rect 38519 16068 38568 16096
rect 38519 16065 38531 16068
rect 38473 16059 38531 16065
rect 38396 16028 38424 16059
rect 38562 16056 38568 16068
rect 38620 16056 38626 16108
rect 38654 16056 38660 16108
rect 38712 16056 38718 16108
rect 39316 16105 39344 16136
rect 39482 16124 39488 16176
rect 39540 16124 39546 16176
rect 39684 16105 39712 16204
rect 39850 16192 39856 16244
rect 39908 16192 39914 16244
rect 41230 16232 41236 16244
rect 40052 16204 41236 16232
rect 39117 16099 39175 16105
rect 39117 16065 39129 16099
rect 39163 16065 39175 16099
rect 39117 16059 39175 16065
rect 39301 16099 39359 16105
rect 39301 16065 39313 16099
rect 39347 16065 39359 16099
rect 39301 16059 39359 16065
rect 39577 16099 39635 16105
rect 39577 16065 39589 16099
rect 39623 16065 39635 16099
rect 39577 16059 39635 16065
rect 39669 16099 39727 16105
rect 39669 16065 39681 16099
rect 39715 16096 39727 16099
rect 39942 16096 39948 16108
rect 39715 16068 39948 16096
rect 39715 16065 39727 16068
rect 39669 16059 39727 16065
rect 38838 16028 38844 16040
rect 38396 16000 38844 16028
rect 38838 15988 38844 16000
rect 38896 16028 38902 16040
rect 38896 16000 38976 16028
rect 38896 15988 38902 16000
rect 37936 15932 38608 15960
rect 38580 15904 38608 15932
rect 29788 15864 30696 15892
rect 29788 15852 29794 15864
rect 31018 15852 31024 15904
rect 31076 15892 31082 15904
rect 31297 15895 31355 15901
rect 31297 15892 31309 15895
rect 31076 15864 31309 15892
rect 31076 15852 31082 15864
rect 31297 15861 31309 15864
rect 31343 15892 31355 15895
rect 34054 15892 34060 15904
rect 31343 15864 34060 15892
rect 31343 15861 31355 15864
rect 31297 15855 31355 15861
rect 34054 15852 34060 15864
rect 34112 15852 34118 15904
rect 35710 15852 35716 15904
rect 35768 15852 35774 15904
rect 35802 15852 35808 15904
rect 35860 15892 35866 15904
rect 36173 15895 36231 15901
rect 36173 15892 36185 15895
rect 35860 15864 36185 15892
rect 35860 15852 35866 15864
rect 36173 15861 36185 15864
rect 36219 15892 36231 15895
rect 36814 15892 36820 15904
rect 36219 15864 36820 15892
rect 36219 15861 36231 15864
rect 36173 15855 36231 15861
rect 36814 15852 36820 15864
rect 36872 15852 36878 15904
rect 37826 15852 37832 15904
rect 37884 15852 37890 15904
rect 38102 15852 38108 15904
rect 38160 15852 38166 15904
rect 38562 15852 38568 15904
rect 38620 15892 38626 15904
rect 38841 15895 38899 15901
rect 38841 15892 38853 15895
rect 38620 15864 38853 15892
rect 38620 15852 38626 15864
rect 38841 15861 38853 15864
rect 38887 15861 38899 15895
rect 38948 15892 38976 16000
rect 39132 15960 39160 16059
rect 39592 16028 39620 16059
rect 39942 16056 39948 16068
rect 40000 16056 40006 16108
rect 40052 16105 40080 16204
rect 41230 16192 41236 16204
rect 41288 16192 41294 16244
rect 44174 16192 44180 16244
rect 44232 16232 44238 16244
rect 44453 16235 44511 16241
rect 44453 16232 44465 16235
rect 44232 16204 44465 16232
rect 44232 16192 44238 16204
rect 44453 16201 44465 16204
rect 44499 16201 44511 16235
rect 44453 16195 44511 16201
rect 47397 16235 47455 16241
rect 47397 16201 47409 16235
rect 47443 16232 47455 16235
rect 47578 16232 47584 16244
rect 47443 16204 47584 16232
rect 47443 16201 47455 16204
rect 47397 16195 47455 16201
rect 47578 16192 47584 16204
rect 47636 16192 47642 16244
rect 47670 16192 47676 16244
rect 47728 16232 47734 16244
rect 48406 16232 48412 16244
rect 47728 16204 48412 16232
rect 47728 16192 47734 16204
rect 48406 16192 48412 16204
rect 48464 16192 48470 16244
rect 49329 16235 49387 16241
rect 49329 16201 49341 16235
rect 49375 16232 49387 16235
rect 49602 16232 49608 16244
rect 49375 16204 49608 16232
rect 49375 16201 49387 16204
rect 49329 16195 49387 16201
rect 49602 16192 49608 16204
rect 49660 16192 49666 16244
rect 49694 16192 49700 16244
rect 49752 16192 49758 16244
rect 49789 16235 49847 16241
rect 49789 16201 49801 16235
rect 49835 16201 49847 16235
rect 49789 16195 49847 16201
rect 40310 16124 40316 16176
rect 40368 16124 40374 16176
rect 40862 16124 40868 16176
rect 40920 16124 40926 16176
rect 42794 16124 42800 16176
rect 42852 16164 42858 16176
rect 42889 16167 42947 16173
rect 42889 16164 42901 16167
rect 42852 16136 42901 16164
rect 42852 16124 42858 16136
rect 42889 16133 42901 16136
rect 42935 16133 42947 16167
rect 49804 16164 49832 16195
rect 50246 16192 50252 16244
rect 50304 16232 50310 16244
rect 50433 16235 50491 16241
rect 50433 16232 50445 16235
rect 50304 16204 50445 16232
rect 50304 16192 50310 16204
rect 50433 16201 50445 16204
rect 50479 16201 50491 16235
rect 53282 16232 53288 16244
rect 50433 16195 50491 16201
rect 52840 16204 53288 16232
rect 52840 16173 52868 16204
rect 53282 16192 53288 16204
rect 53340 16192 53346 16244
rect 53374 16192 53380 16244
rect 53432 16232 53438 16244
rect 54754 16232 54760 16244
rect 53432 16204 54760 16232
rect 53432 16192 53438 16204
rect 54754 16192 54760 16204
rect 54812 16232 54818 16244
rect 56042 16232 56048 16244
rect 54812 16204 56048 16232
rect 54812 16192 54818 16204
rect 56042 16192 56048 16204
rect 56100 16192 56106 16244
rect 50157 16167 50215 16173
rect 50157 16164 50169 16167
rect 42889 16127 42947 16133
rect 44376 16136 45048 16164
rect 40037 16099 40095 16105
rect 40037 16065 40049 16099
rect 40083 16065 40095 16099
rect 40037 16059 40095 16065
rect 43990 16056 43996 16108
rect 44048 16056 44054 16108
rect 40402 16028 40408 16040
rect 39592 16000 40408 16028
rect 40402 15988 40408 16000
rect 40460 15988 40466 16040
rect 42613 16031 42671 16037
rect 42613 15997 42625 16031
rect 42659 16028 42671 16031
rect 42659 16000 42748 16028
rect 42659 15997 42671 16000
rect 42613 15991 42671 15997
rect 39390 15960 39396 15972
rect 39132 15932 39396 15960
rect 39390 15920 39396 15932
rect 39448 15960 39454 15972
rect 39666 15960 39672 15972
rect 39448 15932 39672 15960
rect 39448 15920 39454 15932
rect 39666 15920 39672 15932
rect 39724 15920 39730 15972
rect 41782 15892 41788 15904
rect 38948 15864 41788 15892
rect 38841 15855 38899 15861
rect 41782 15852 41788 15864
rect 41840 15852 41846 15904
rect 42720 15892 42748 16000
rect 43254 15988 43260 16040
rect 43312 16028 43318 16040
rect 44376 16037 44404 16136
rect 44637 16099 44695 16105
rect 44637 16065 44649 16099
rect 44683 16065 44695 16099
rect 44637 16059 44695 16065
rect 44361 16031 44419 16037
rect 44361 16028 44373 16031
rect 43312 16000 44373 16028
rect 43312 15988 43318 16000
rect 44361 15997 44373 16000
rect 44407 15997 44419 16031
rect 44361 15991 44419 15997
rect 44542 15988 44548 16040
rect 44600 16028 44606 16040
rect 44652 16028 44680 16059
rect 44726 16056 44732 16108
rect 44784 16056 44790 16108
rect 45020 16105 45048 16136
rect 48332 16136 49832 16164
rect 49896 16136 50169 16164
rect 44821 16099 44879 16105
rect 44821 16065 44833 16099
rect 44867 16065 44879 16099
rect 44821 16059 44879 16065
rect 45005 16099 45063 16105
rect 45005 16065 45017 16099
rect 45051 16065 45063 16099
rect 45005 16059 45063 16065
rect 44836 16028 44864 16059
rect 46566 16056 46572 16108
rect 46624 16056 46630 16108
rect 47394 16056 47400 16108
rect 47452 16096 47458 16108
rect 47762 16096 47768 16108
rect 47452 16068 47768 16096
rect 47452 16056 47458 16068
rect 47762 16056 47768 16068
rect 47820 16096 47826 16108
rect 48332 16105 48360 16136
rect 48133 16099 48191 16105
rect 48133 16096 48145 16099
rect 47820 16068 48145 16096
rect 47820 16056 47826 16068
rect 48133 16065 48145 16068
rect 48179 16065 48191 16099
rect 48133 16059 48191 16065
rect 48317 16099 48375 16105
rect 48317 16065 48329 16099
rect 48363 16065 48375 16099
rect 48317 16059 48375 16065
rect 48410 16099 48468 16105
rect 48410 16065 48422 16099
rect 48456 16065 48468 16099
rect 48410 16059 48468 16065
rect 44600 16000 44680 16028
rect 44744 16000 44864 16028
rect 44600 15988 44606 16000
rect 43438 15892 43444 15904
rect 42720 15864 43444 15892
rect 43438 15852 43444 15864
rect 43496 15852 43502 15904
rect 43622 15852 43628 15904
rect 43680 15892 43686 15904
rect 44744 15892 44772 16000
rect 45370 15988 45376 16040
rect 45428 16028 45434 16040
rect 46753 16031 46811 16037
rect 46753 16028 46765 16031
rect 45428 16000 46765 16028
rect 45428 15988 45434 16000
rect 46753 15997 46765 16000
rect 46799 15997 46811 16031
rect 46753 15991 46811 15997
rect 46845 16031 46903 16037
rect 46845 15997 46857 16031
rect 46891 16028 46903 16031
rect 47581 16031 47639 16037
rect 47581 16028 47593 16031
rect 46891 16000 47593 16028
rect 46891 15997 46903 16000
rect 46845 15991 46903 15997
rect 47581 15997 47593 16000
rect 47627 15997 47639 16031
rect 47581 15991 47639 15997
rect 48222 15988 48228 16040
rect 48280 16028 48286 16040
rect 48424 16028 48452 16059
rect 48590 16056 48596 16108
rect 48648 16056 48654 16108
rect 48682 16056 48688 16108
rect 48740 16056 48746 16108
rect 48782 16099 48840 16105
rect 48782 16065 48794 16099
rect 48828 16065 48840 16099
rect 48782 16059 48840 16065
rect 48280 16000 48452 16028
rect 48280 15988 48286 16000
rect 48038 15920 48044 15972
rect 48096 15960 48102 15972
rect 48096 15932 48314 15960
rect 48096 15920 48102 15932
rect 45646 15892 45652 15904
rect 43680 15864 45652 15892
rect 43680 15852 43686 15864
rect 45646 15852 45652 15864
rect 45704 15852 45710 15904
rect 45922 15852 45928 15904
rect 45980 15892 45986 15904
rect 46385 15895 46443 15901
rect 46385 15892 46397 15895
rect 45980 15864 46397 15892
rect 45980 15852 45986 15864
rect 46385 15861 46397 15864
rect 46431 15861 46443 15895
rect 48286 15892 48314 15932
rect 48406 15920 48412 15972
rect 48464 15960 48470 15972
rect 48797 15960 48825 16059
rect 48958 16056 48964 16108
rect 49016 16096 49022 16108
rect 49053 16099 49111 16105
rect 49053 16096 49065 16099
rect 49016 16068 49065 16096
rect 49016 16056 49022 16068
rect 49053 16065 49065 16068
rect 49099 16065 49111 16099
rect 49053 16059 49111 16065
rect 49418 16056 49424 16108
rect 49476 16056 49482 16108
rect 49694 16056 49700 16108
rect 49752 16096 49758 16108
rect 49896 16096 49924 16136
rect 50157 16133 50169 16136
rect 50203 16133 50215 16167
rect 50157 16127 50215 16133
rect 52825 16167 52883 16173
rect 52825 16133 52837 16167
rect 52871 16133 52883 16167
rect 55217 16167 55275 16173
rect 55217 16164 55229 16167
rect 52825 16127 52883 16133
rect 54588 16136 55229 16164
rect 49752 16068 49924 16096
rect 49973 16099 50031 16105
rect 49752 16056 49758 16068
rect 49973 16065 49985 16099
rect 50019 16065 50031 16099
rect 49973 16059 50031 16065
rect 49988 16028 50016 16059
rect 50062 16056 50068 16108
rect 50120 16056 50126 16108
rect 50341 16099 50399 16105
rect 50341 16065 50353 16099
rect 50387 16096 50399 16099
rect 51350 16096 51356 16108
rect 50387 16068 51356 16096
rect 50387 16065 50399 16068
rect 50341 16059 50399 16065
rect 51350 16056 51356 16068
rect 51408 16056 51414 16108
rect 54588 16105 54616 16136
rect 55217 16133 55229 16136
rect 55263 16133 55275 16167
rect 55217 16127 55275 16133
rect 54297 16099 54355 16105
rect 54297 16096 54309 16099
rect 53760 16068 54309 16096
rect 50154 16028 50160 16040
rect 49988 16000 50160 16028
rect 50154 15988 50160 16000
rect 50212 15988 50218 16040
rect 51074 15988 51080 16040
rect 51132 16028 51138 16040
rect 53760 16028 53788 16068
rect 54297 16065 54309 16068
rect 54343 16096 54355 16099
rect 54573 16099 54631 16105
rect 54573 16096 54585 16099
rect 54343 16068 54585 16096
rect 54343 16065 54355 16068
rect 54297 16059 54355 16065
rect 54573 16065 54585 16068
rect 54619 16065 54631 16099
rect 54573 16059 54631 16065
rect 54754 16056 54760 16108
rect 54812 16096 54818 16108
rect 54938 16096 54944 16108
rect 54812 16068 54944 16096
rect 54812 16056 54818 16068
rect 54938 16056 54944 16068
rect 54996 16096 55002 16108
rect 55033 16099 55091 16105
rect 55033 16096 55045 16099
rect 54996 16068 55045 16096
rect 54996 16056 55002 16068
rect 55033 16065 55045 16068
rect 55079 16065 55091 16099
rect 55232 16096 55260 16127
rect 55306 16124 55312 16176
rect 55364 16124 55370 16176
rect 56686 16124 56692 16176
rect 56744 16124 56750 16176
rect 55493 16099 55551 16105
rect 55493 16096 55505 16099
rect 55232 16068 55505 16096
rect 55033 16059 55091 16065
rect 55493 16065 55505 16068
rect 55539 16096 55551 16099
rect 55674 16096 55680 16108
rect 55539 16068 55680 16096
rect 55539 16065 55551 16068
rect 55493 16059 55551 16065
rect 55674 16056 55680 16068
rect 55732 16056 55738 16108
rect 51132 16000 53788 16028
rect 51132 15988 51138 16000
rect 53926 15988 53932 16040
rect 53984 16028 53990 16040
rect 55953 16031 56011 16037
rect 55953 16028 55965 16031
rect 53984 16000 55965 16028
rect 53984 15988 53990 16000
rect 55953 15997 55965 16000
rect 55999 15997 56011 16031
rect 55953 15991 56011 15997
rect 56229 16031 56287 16037
rect 56229 15997 56241 16031
rect 56275 16028 56287 16031
rect 56594 16028 56600 16040
rect 56275 16000 56600 16028
rect 56275 15997 56287 16000
rect 56229 15991 56287 15997
rect 56594 15988 56600 16000
rect 56652 15988 56658 16040
rect 48464 15932 48825 15960
rect 48961 15963 49019 15969
rect 48464 15920 48470 15932
rect 48961 15929 48973 15963
rect 49007 15960 49019 15963
rect 49050 15960 49056 15972
rect 49007 15932 49056 15960
rect 49007 15929 49019 15932
rect 48961 15923 49019 15929
rect 49050 15920 49056 15932
rect 49108 15920 49114 15972
rect 52914 15920 52920 15972
rect 52972 15960 52978 15972
rect 54481 15963 54539 15969
rect 54481 15960 54493 15963
rect 52972 15932 54493 15960
rect 52972 15920 52978 15932
rect 54481 15929 54493 15932
rect 54527 15960 54539 15963
rect 55398 15960 55404 15972
rect 54527 15932 55404 15960
rect 54527 15929 54539 15932
rect 54481 15923 54539 15929
rect 55398 15920 55404 15932
rect 55456 15920 55462 15972
rect 52822 15892 52828 15904
rect 48286 15864 52828 15892
rect 46385 15855 46443 15861
rect 52822 15852 52828 15864
rect 52880 15852 52886 15904
rect 53101 15895 53159 15901
rect 53101 15861 53113 15895
rect 53147 15892 53159 15895
rect 53742 15892 53748 15904
rect 53147 15864 53748 15892
rect 53147 15861 53159 15864
rect 53101 15855 53159 15861
rect 53742 15852 53748 15864
rect 53800 15852 53806 15904
rect 55950 15852 55956 15904
rect 56008 15892 56014 15904
rect 57238 15892 57244 15904
rect 56008 15864 57244 15892
rect 56008 15852 56014 15864
rect 57238 15852 57244 15864
rect 57296 15852 57302 15904
rect 57698 15852 57704 15904
rect 57756 15852 57762 15904
rect 1104 15802 58880 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 58880 15802
rect 1104 15728 58880 15750
rect 13265 15691 13323 15697
rect 13265 15657 13277 15691
rect 13311 15688 13323 15691
rect 13311 15660 14780 15688
rect 13311 15657 13323 15660
rect 13265 15651 13323 15657
rect 12437 15555 12495 15561
rect 12437 15521 12449 15555
rect 12483 15521 12495 15555
rect 12437 15515 12495 15521
rect 12897 15555 12955 15561
rect 12897 15521 12909 15555
rect 12943 15552 12955 15555
rect 13262 15552 13268 15564
rect 12943 15524 13268 15552
rect 12943 15521 12955 15524
rect 12897 15515 12955 15521
rect 12452 15416 12480 15515
rect 13262 15512 13268 15524
rect 13320 15512 13326 15564
rect 14752 15493 14780 15660
rect 18874 15648 18880 15700
rect 18932 15688 18938 15700
rect 19613 15691 19671 15697
rect 19613 15688 19625 15691
rect 18932 15660 19625 15688
rect 18932 15648 18938 15660
rect 19613 15657 19625 15660
rect 19659 15688 19671 15691
rect 19889 15691 19947 15697
rect 19889 15688 19901 15691
rect 19659 15660 19901 15688
rect 19659 15657 19671 15660
rect 19613 15651 19671 15657
rect 19889 15657 19901 15660
rect 19935 15688 19947 15691
rect 20070 15688 20076 15700
rect 19935 15660 20076 15688
rect 19935 15657 19947 15660
rect 19889 15651 19947 15657
rect 20070 15648 20076 15660
rect 20128 15648 20134 15700
rect 20162 15648 20168 15700
rect 20220 15688 20226 15700
rect 22186 15688 22192 15700
rect 20220 15660 22192 15688
rect 20220 15648 20226 15660
rect 22186 15648 22192 15660
rect 22244 15688 22250 15700
rect 22554 15688 22560 15700
rect 22244 15660 22560 15688
rect 22244 15648 22250 15660
rect 22554 15648 22560 15660
rect 22612 15688 22618 15700
rect 23474 15688 23480 15700
rect 22612 15660 23480 15688
rect 22612 15648 22618 15660
rect 23474 15648 23480 15660
rect 23532 15648 23538 15700
rect 24210 15648 24216 15700
rect 24268 15688 24274 15700
rect 24670 15688 24676 15700
rect 24268 15660 24676 15688
rect 24268 15648 24274 15660
rect 24670 15648 24676 15660
rect 24728 15688 24734 15700
rect 24728 15660 24808 15688
rect 24728 15648 24734 15660
rect 19978 15620 19984 15632
rect 19720 15592 19984 15620
rect 19720 15561 19748 15592
rect 19978 15580 19984 15592
rect 20036 15620 20042 15632
rect 24486 15620 24492 15632
rect 20036 15592 24492 15620
rect 20036 15580 20042 15592
rect 24486 15580 24492 15592
rect 24544 15580 24550 15632
rect 24780 15620 24808 15660
rect 24854 15648 24860 15700
rect 24912 15648 24918 15700
rect 26602 15648 26608 15700
rect 26660 15688 26666 15700
rect 27065 15691 27123 15697
rect 27065 15688 27077 15691
rect 26660 15660 27077 15688
rect 26660 15648 26666 15660
rect 27065 15657 27077 15660
rect 27111 15657 27123 15691
rect 27065 15651 27123 15657
rect 28966 15660 30328 15688
rect 25501 15623 25559 15629
rect 25501 15620 25513 15623
rect 24780 15592 25513 15620
rect 25501 15589 25513 15592
rect 25547 15620 25559 15623
rect 26326 15620 26332 15632
rect 25547 15592 26332 15620
rect 25547 15589 25559 15592
rect 25501 15583 25559 15589
rect 26326 15580 26332 15592
rect 26384 15580 26390 15632
rect 26694 15580 26700 15632
rect 26752 15620 26758 15632
rect 26973 15623 27031 15629
rect 26973 15620 26985 15623
rect 26752 15592 26985 15620
rect 26752 15580 26758 15592
rect 26973 15589 26985 15592
rect 27019 15620 27031 15623
rect 28718 15620 28724 15632
rect 27019 15592 28724 15620
rect 27019 15589 27031 15592
rect 26973 15583 27031 15589
rect 28718 15580 28724 15592
rect 28776 15580 28782 15632
rect 19705 15555 19763 15561
rect 19705 15521 19717 15555
rect 19751 15521 19763 15555
rect 19705 15515 19763 15521
rect 21542 15512 21548 15564
rect 21600 15552 21606 15564
rect 22465 15555 22523 15561
rect 21600 15524 22416 15552
rect 21600 15512 21606 15524
rect 22388 15496 22416 15524
rect 22465 15521 22477 15555
rect 22511 15552 22523 15555
rect 23566 15552 23572 15564
rect 22511 15524 23572 15552
rect 22511 15521 22523 15524
rect 22465 15515 22523 15521
rect 23566 15512 23572 15524
rect 23624 15552 23630 15564
rect 23842 15552 23848 15564
rect 23624 15524 23848 15552
rect 23624 15512 23630 15524
rect 23842 15512 23848 15524
rect 23900 15512 23906 15564
rect 24026 15512 24032 15564
rect 24084 15552 24090 15564
rect 24762 15552 24768 15564
rect 24084 15524 24768 15552
rect 24084 15512 24090 15524
rect 24762 15512 24768 15524
rect 24820 15552 24826 15564
rect 25409 15555 25467 15561
rect 25409 15552 25421 15555
rect 24820 15524 25421 15552
rect 24820 15512 24826 15524
rect 25409 15521 25421 15524
rect 25455 15521 25467 15555
rect 25409 15515 25467 15521
rect 26510 15512 26516 15564
rect 26568 15552 26574 15564
rect 28966 15552 28994 15660
rect 26568 15524 28994 15552
rect 26568 15512 26574 15524
rect 30190 15512 30196 15564
rect 30248 15512 30254 15564
rect 12529 15487 12587 15493
rect 12529 15453 12541 15487
rect 12575 15484 12587 15487
rect 14093 15487 14151 15493
rect 14093 15484 14105 15487
rect 12575 15456 14105 15484
rect 12575 15453 12587 15456
rect 12529 15447 12587 15453
rect 14093 15453 14105 15456
rect 14139 15453 14151 15487
rect 14093 15447 14151 15453
rect 14737 15487 14795 15493
rect 14737 15453 14749 15487
rect 14783 15484 14795 15487
rect 14918 15484 14924 15496
rect 14783 15456 14924 15484
rect 14783 15453 14795 15456
rect 14737 15447 14795 15453
rect 14918 15444 14924 15456
rect 14976 15444 14982 15496
rect 19429 15487 19487 15493
rect 19429 15453 19441 15487
rect 19475 15453 19487 15487
rect 19429 15447 19487 15453
rect 12618 15416 12624 15428
rect 12452 15388 12624 15416
rect 12618 15376 12624 15388
rect 12676 15416 12682 15428
rect 12676 15388 13216 15416
rect 12676 15376 12682 15388
rect 12710 15308 12716 15360
rect 12768 15348 12774 15360
rect 13081 15351 13139 15357
rect 13081 15348 13093 15351
rect 12768 15320 13093 15348
rect 12768 15308 12774 15320
rect 13081 15317 13093 15320
rect 13127 15317 13139 15351
rect 13188 15348 13216 15388
rect 13446 15376 13452 15428
rect 13504 15376 13510 15428
rect 19444 15416 19472 15447
rect 19794 15444 19800 15496
rect 19852 15444 19858 15496
rect 20070 15444 20076 15496
rect 20128 15444 20134 15496
rect 20254 15444 20260 15496
rect 20312 15444 20318 15496
rect 22186 15444 22192 15496
rect 22244 15444 22250 15496
rect 22370 15444 22376 15496
rect 22428 15444 22434 15496
rect 22922 15444 22928 15496
rect 22980 15444 22986 15496
rect 23106 15444 23112 15496
rect 23164 15444 23170 15496
rect 23201 15487 23259 15493
rect 23201 15453 23213 15487
rect 23247 15484 23259 15487
rect 23382 15484 23388 15496
rect 23247 15456 23388 15484
rect 23247 15453 23259 15456
rect 23201 15447 23259 15453
rect 23382 15444 23388 15456
rect 23440 15444 23446 15496
rect 24486 15444 24492 15496
rect 24544 15484 24550 15496
rect 24673 15487 24731 15493
rect 24673 15484 24685 15487
rect 24544 15456 24685 15484
rect 24544 15444 24550 15456
rect 24673 15453 24685 15456
rect 24719 15453 24731 15487
rect 24673 15447 24731 15453
rect 20272 15416 20300 15444
rect 19444 15388 20300 15416
rect 23290 15376 23296 15428
rect 23348 15376 23354 15428
rect 24118 15376 24124 15428
rect 24176 15376 24182 15428
rect 24688 15416 24716 15447
rect 25682 15444 25688 15496
rect 25740 15444 25746 15496
rect 29638 15444 29644 15496
rect 29696 15484 29702 15496
rect 29917 15487 29975 15493
rect 29917 15484 29929 15487
rect 29696 15456 29929 15484
rect 29696 15444 29702 15456
rect 25958 15416 25964 15428
rect 24688 15388 25964 15416
rect 25958 15376 25964 15388
rect 26016 15416 26022 15428
rect 26694 15416 26700 15428
rect 26016 15388 26700 15416
rect 26016 15376 26022 15388
rect 26694 15376 26700 15388
rect 26752 15416 26758 15428
rect 27338 15416 27344 15428
rect 26752 15388 27344 15416
rect 26752 15376 26758 15388
rect 27338 15376 27344 15388
rect 27396 15376 27402 15428
rect 13249 15351 13307 15357
rect 13249 15348 13261 15351
rect 13188 15320 13261 15348
rect 13081 15311 13139 15317
rect 13249 15317 13261 15320
rect 13295 15348 13307 15351
rect 15102 15348 15108 15360
rect 13295 15320 15108 15348
rect 13295 15317 13307 15320
rect 13249 15311 13307 15317
rect 15102 15308 15108 15320
rect 15160 15308 15166 15360
rect 18138 15308 18144 15360
rect 18196 15348 18202 15360
rect 19245 15351 19303 15357
rect 19245 15348 19257 15351
rect 18196 15320 19257 15348
rect 18196 15308 18202 15320
rect 19245 15317 19257 15320
rect 19291 15317 19303 15351
rect 19245 15311 19303 15317
rect 20257 15351 20315 15357
rect 20257 15317 20269 15351
rect 20303 15348 20315 15351
rect 20714 15348 20720 15360
rect 20303 15320 20720 15348
rect 20303 15317 20315 15320
rect 20257 15311 20315 15317
rect 20714 15308 20720 15320
rect 20772 15308 20778 15360
rect 21726 15308 21732 15360
rect 21784 15348 21790 15360
rect 22005 15351 22063 15357
rect 22005 15348 22017 15351
rect 21784 15320 22017 15348
rect 21784 15308 21790 15320
rect 22005 15317 22017 15320
rect 22051 15317 22063 15351
rect 22005 15311 22063 15317
rect 22094 15308 22100 15360
rect 22152 15348 22158 15360
rect 22741 15351 22799 15357
rect 22741 15348 22753 15351
rect 22152 15320 22753 15348
rect 22152 15308 22158 15320
rect 22741 15317 22753 15320
rect 22787 15317 22799 15351
rect 22741 15311 22799 15317
rect 23474 15308 23480 15360
rect 23532 15348 23538 15360
rect 24489 15351 24547 15357
rect 24489 15348 24501 15351
rect 23532 15320 24501 15348
rect 23532 15308 23538 15320
rect 24489 15317 24501 15320
rect 24535 15317 24547 15351
rect 24489 15311 24547 15317
rect 25869 15351 25927 15357
rect 25869 15317 25881 15351
rect 25915 15348 25927 15351
rect 26234 15348 26240 15360
rect 25915 15320 26240 15348
rect 25915 15317 25927 15320
rect 25869 15311 25927 15317
rect 26234 15308 26240 15320
rect 26292 15308 26298 15360
rect 29748 15348 29776 15456
rect 29917 15453 29929 15456
rect 29963 15453 29975 15487
rect 29917 15447 29975 15453
rect 30065 15487 30123 15493
rect 30065 15453 30077 15487
rect 30111 15484 30123 15487
rect 30208 15484 30236 15512
rect 30300 15496 30328 15660
rect 34514 15648 34520 15700
rect 34572 15688 34578 15700
rect 34572 15660 36492 15688
rect 34572 15648 34578 15660
rect 30561 15623 30619 15629
rect 30561 15589 30573 15623
rect 30607 15589 30619 15623
rect 30561 15583 30619 15589
rect 30111 15456 30236 15484
rect 30111 15453 30123 15456
rect 30065 15447 30123 15453
rect 30282 15444 30288 15496
rect 30340 15444 30346 15496
rect 30466 15493 30472 15496
rect 30423 15487 30472 15493
rect 30423 15453 30435 15487
rect 30469 15453 30472 15487
rect 30423 15447 30472 15453
rect 30466 15444 30472 15447
rect 30524 15444 30530 15496
rect 30576 15484 30604 15583
rect 31018 15580 31024 15632
rect 31076 15580 31082 15632
rect 36464 15620 36492 15660
rect 36538 15648 36544 15700
rect 36596 15688 36602 15700
rect 36633 15691 36691 15697
rect 36633 15688 36645 15691
rect 36596 15660 36645 15688
rect 36596 15648 36602 15660
rect 36633 15657 36645 15660
rect 36679 15657 36691 15691
rect 38286 15688 38292 15700
rect 36633 15651 36691 15657
rect 37384 15660 38292 15688
rect 37384 15620 37412 15660
rect 38286 15648 38292 15660
rect 38344 15648 38350 15700
rect 38580 15660 38976 15688
rect 36464 15592 37412 15620
rect 30742 15512 30748 15564
rect 30800 15552 30806 15564
rect 31113 15555 31171 15561
rect 31113 15552 31125 15555
rect 30800 15524 31125 15552
rect 30800 15512 30806 15524
rect 31113 15521 31125 15524
rect 31159 15552 31171 15555
rect 31573 15555 31631 15561
rect 31573 15552 31585 15555
rect 31159 15524 31585 15552
rect 31159 15521 31171 15524
rect 31113 15515 31171 15521
rect 31573 15521 31585 15524
rect 31619 15521 31631 15555
rect 31573 15515 31631 15521
rect 32122 15512 32128 15564
rect 32180 15512 32186 15564
rect 33502 15552 33508 15564
rect 33060 15524 33508 15552
rect 30837 15487 30895 15493
rect 30837 15484 30849 15487
rect 30576 15456 30849 15484
rect 30837 15453 30849 15456
rect 30883 15453 30895 15487
rect 30837 15447 30895 15453
rect 32582 15444 32588 15496
rect 32640 15484 32646 15496
rect 33060 15493 33088 15524
rect 33502 15512 33508 15524
rect 33560 15552 33566 15564
rect 34885 15555 34943 15561
rect 34885 15552 34897 15555
rect 33560 15524 34897 15552
rect 33560 15512 33566 15524
rect 34885 15521 34897 15524
rect 34931 15521 34943 15555
rect 34885 15515 34943 15521
rect 35161 15555 35219 15561
rect 35161 15521 35173 15555
rect 35207 15552 35219 15555
rect 35710 15552 35716 15564
rect 35207 15524 35716 15552
rect 35207 15521 35219 15524
rect 35161 15515 35219 15521
rect 35710 15512 35716 15524
rect 35768 15512 35774 15564
rect 38194 15512 38200 15564
rect 38252 15552 38258 15564
rect 38580 15552 38608 15660
rect 38654 15580 38660 15632
rect 38712 15580 38718 15632
rect 38948 15620 38976 15660
rect 39022 15648 39028 15700
rect 39080 15648 39086 15700
rect 39393 15691 39451 15697
rect 39393 15657 39405 15691
rect 39439 15688 39451 15691
rect 40310 15688 40316 15700
rect 39439 15660 40316 15688
rect 39439 15657 39451 15660
rect 39393 15651 39451 15657
rect 39114 15620 39120 15632
rect 38948 15592 39120 15620
rect 39114 15580 39120 15592
rect 39172 15620 39178 15632
rect 39408 15620 39436 15651
rect 40310 15648 40316 15660
rect 40368 15648 40374 15700
rect 40497 15691 40555 15697
rect 40497 15657 40509 15691
rect 40543 15688 40555 15691
rect 40678 15688 40684 15700
rect 40543 15660 40684 15688
rect 40543 15657 40555 15660
rect 40497 15651 40555 15657
rect 40678 15648 40684 15660
rect 40736 15648 40742 15700
rect 42981 15691 43039 15697
rect 42981 15657 42993 15691
rect 43027 15688 43039 15691
rect 43070 15688 43076 15700
rect 43027 15660 43076 15688
rect 43027 15657 43039 15660
rect 42981 15651 43039 15657
rect 43070 15648 43076 15660
rect 43128 15648 43134 15700
rect 47670 15648 47676 15700
rect 47728 15688 47734 15700
rect 48133 15691 48191 15697
rect 48133 15688 48145 15691
rect 47728 15660 48145 15688
rect 47728 15648 47734 15660
rect 48133 15657 48145 15660
rect 48179 15657 48191 15691
rect 48133 15651 48191 15657
rect 48774 15648 48780 15700
rect 48832 15688 48838 15700
rect 48961 15691 49019 15697
rect 48961 15688 48973 15691
rect 48832 15660 48973 15688
rect 48832 15648 48838 15660
rect 48961 15657 48973 15660
rect 49007 15688 49019 15691
rect 49234 15688 49240 15700
rect 49007 15660 49240 15688
rect 49007 15657 49019 15660
rect 48961 15651 49019 15657
rect 49234 15648 49240 15660
rect 49292 15648 49298 15700
rect 51350 15648 51356 15700
rect 51408 15688 51414 15700
rect 54754 15688 54760 15700
rect 51408 15660 54760 15688
rect 51408 15648 51414 15660
rect 54754 15648 54760 15660
rect 54812 15688 54818 15700
rect 55861 15691 55919 15697
rect 54812 15660 55076 15688
rect 54812 15648 54818 15660
rect 39172 15592 39436 15620
rect 39172 15580 39178 15592
rect 39482 15580 39488 15632
rect 39540 15620 39546 15632
rect 42610 15620 42616 15632
rect 39540 15592 42616 15620
rect 39540 15580 39546 15592
rect 42610 15580 42616 15592
rect 42668 15580 42674 15632
rect 48038 15580 48044 15632
rect 48096 15620 48102 15632
rect 48590 15620 48596 15632
rect 48096 15592 48596 15620
rect 48096 15580 48102 15592
rect 48590 15580 48596 15592
rect 48648 15580 48654 15632
rect 48682 15580 48688 15632
rect 48740 15620 48746 15632
rect 48740 15592 49924 15620
rect 48740 15580 48746 15592
rect 38252 15524 38608 15552
rect 38672 15552 38700 15580
rect 49896 15564 49924 15592
rect 51902 15580 51908 15632
rect 51960 15580 51966 15632
rect 52012 15592 52408 15620
rect 40034 15552 40040 15564
rect 38672 15524 40040 15552
rect 38252 15512 38258 15524
rect 40034 15512 40040 15524
rect 40092 15552 40098 15564
rect 40865 15555 40923 15561
rect 40092 15524 40172 15552
rect 40092 15512 40098 15524
rect 33045 15487 33103 15493
rect 33045 15484 33057 15487
rect 32640 15456 33057 15484
rect 32640 15444 32646 15456
rect 33045 15453 33057 15456
rect 33091 15453 33103 15487
rect 33045 15447 33103 15453
rect 37274 15444 37280 15496
rect 37332 15444 37338 15496
rect 39022 15444 39028 15496
rect 39080 15484 39086 15496
rect 40144 15493 40172 15524
rect 40865 15521 40877 15555
rect 40911 15521 40923 15555
rect 40865 15515 40923 15521
rect 39945 15487 40003 15493
rect 39945 15484 39957 15487
rect 39080 15456 39957 15484
rect 39080 15444 39086 15456
rect 39945 15453 39957 15456
rect 39991 15453 40003 15487
rect 39945 15447 40003 15453
rect 40129 15487 40187 15493
rect 40129 15453 40141 15487
rect 40175 15453 40187 15487
rect 40129 15447 40187 15453
rect 40218 15444 40224 15496
rect 40276 15444 40282 15496
rect 40310 15444 40316 15496
rect 40368 15444 40374 15496
rect 40880 15484 40908 15515
rect 43438 15512 43444 15564
rect 43496 15552 43502 15564
rect 44910 15552 44916 15564
rect 43496 15524 44916 15552
rect 43496 15512 43502 15524
rect 44910 15512 44916 15524
rect 44968 15552 44974 15564
rect 45649 15555 45707 15561
rect 45649 15552 45661 15555
rect 44968 15524 45661 15552
rect 44968 15512 44974 15524
rect 45649 15521 45661 15524
rect 45695 15552 45707 15555
rect 47946 15552 47952 15564
rect 45695 15524 47952 15552
rect 45695 15521 45707 15524
rect 45649 15515 45707 15521
rect 47946 15512 47952 15524
rect 48004 15512 48010 15564
rect 49878 15512 49884 15564
rect 49936 15552 49942 15564
rect 50709 15555 50767 15561
rect 50709 15552 50721 15555
rect 49936 15524 50721 15552
rect 49936 15512 49942 15524
rect 50709 15521 50721 15524
rect 50755 15521 50767 15555
rect 52012 15552 52040 15592
rect 50709 15515 50767 15521
rect 51552 15524 52040 15552
rect 40420 15456 40908 15484
rect 29822 15376 29828 15428
rect 29880 15416 29886 15428
rect 30193 15419 30251 15425
rect 30193 15416 30205 15419
rect 29880 15388 30205 15416
rect 29880 15376 29886 15388
rect 30193 15385 30205 15388
rect 30239 15385 30251 15419
rect 31297 15419 31355 15425
rect 31297 15416 31309 15419
rect 30193 15379 30251 15385
rect 30397 15388 31309 15416
rect 30397 15348 30425 15388
rect 31297 15385 31309 15388
rect 31343 15416 31355 15419
rect 32766 15416 32772 15428
rect 31343 15388 32772 15416
rect 31343 15385 31355 15388
rect 31297 15379 31355 15385
rect 32766 15376 32772 15388
rect 32824 15376 32830 15428
rect 36386 15388 36676 15416
rect 29748 15320 30425 15348
rect 30466 15308 30472 15360
rect 30524 15348 30530 15360
rect 30653 15351 30711 15357
rect 30653 15348 30665 15351
rect 30524 15320 30665 15348
rect 30524 15308 30530 15320
rect 30653 15317 30665 15320
rect 30699 15317 30711 15351
rect 36648 15348 36676 15388
rect 36722 15376 36728 15428
rect 36780 15416 36786 15428
rect 36817 15419 36875 15425
rect 36817 15416 36829 15419
rect 36780 15388 36829 15416
rect 36780 15376 36786 15388
rect 36817 15385 36829 15388
rect 36863 15385 36875 15419
rect 36817 15379 36875 15385
rect 37550 15376 37556 15428
rect 37608 15376 37614 15428
rect 39206 15416 39212 15428
rect 38778 15388 39212 15416
rect 37093 15351 37151 15357
rect 37093 15348 37105 15351
rect 36648 15320 37105 15348
rect 30653 15311 30711 15317
rect 37093 15317 37105 15320
rect 37139 15348 37151 15351
rect 37366 15348 37372 15360
rect 37139 15320 37372 15348
rect 37139 15317 37151 15320
rect 37093 15311 37151 15317
rect 37366 15308 37372 15320
rect 37424 15348 37430 15360
rect 38856 15348 38884 15388
rect 39206 15376 39212 15388
rect 39264 15376 39270 15428
rect 39298 15376 39304 15428
rect 39356 15416 39362 15428
rect 39485 15419 39543 15425
rect 39485 15416 39497 15419
rect 39356 15388 39497 15416
rect 39356 15376 39362 15388
rect 39485 15385 39497 15388
rect 39531 15416 39543 15419
rect 39850 15416 39856 15428
rect 39531 15388 39856 15416
rect 39531 15385 39543 15388
rect 39485 15379 39543 15385
rect 39850 15376 39856 15388
rect 39908 15376 39914 15428
rect 40420 15416 40448 15456
rect 41782 15444 41788 15496
rect 41840 15484 41846 15496
rect 42429 15487 42487 15493
rect 42429 15484 42441 15487
rect 41840 15456 42441 15484
rect 41840 15444 41846 15456
rect 42429 15453 42441 15456
rect 42475 15453 42487 15487
rect 42429 15447 42487 15453
rect 42797 15487 42855 15493
rect 42797 15453 42809 15487
rect 42843 15484 42855 15487
rect 43346 15484 43352 15496
rect 42843 15456 43352 15484
rect 42843 15453 42855 15456
rect 42797 15447 42855 15453
rect 43346 15444 43352 15456
rect 43404 15444 43410 15496
rect 43530 15444 43536 15496
rect 43588 15444 43594 15496
rect 43622 15444 43628 15496
rect 43680 15484 43686 15496
rect 43717 15487 43775 15493
rect 43717 15484 43729 15487
rect 43680 15456 43729 15484
rect 43680 15444 43686 15456
rect 43717 15453 43729 15456
rect 43763 15453 43775 15487
rect 43717 15447 43775 15453
rect 43901 15487 43959 15493
rect 43901 15453 43913 15487
rect 43947 15484 43959 15487
rect 44082 15484 44088 15496
rect 43947 15456 44088 15484
rect 43947 15453 43959 15456
rect 43901 15447 43959 15453
rect 44082 15444 44088 15456
rect 44140 15484 44146 15496
rect 48685 15487 48743 15493
rect 44140 15456 44680 15484
rect 44140 15444 44146 15456
rect 40236 15388 40448 15416
rect 37424 15320 38884 15348
rect 37424 15308 37430 15320
rect 39574 15308 39580 15360
rect 39632 15348 39638 15360
rect 40236 15348 40264 15388
rect 40494 15376 40500 15428
rect 40552 15416 40558 15428
rect 40862 15416 40868 15428
rect 40552 15388 40868 15416
rect 40552 15376 40558 15388
rect 40862 15376 40868 15388
rect 40920 15376 40926 15428
rect 40954 15376 40960 15428
rect 41012 15416 41018 15428
rect 42518 15416 42524 15428
rect 41012 15388 42524 15416
rect 41012 15376 41018 15388
rect 42518 15376 42524 15388
rect 42576 15376 42582 15428
rect 42613 15419 42671 15425
rect 42613 15385 42625 15419
rect 42659 15385 42671 15419
rect 42613 15379 42671 15385
rect 42705 15419 42763 15425
rect 42705 15385 42717 15419
rect 42751 15416 42763 15419
rect 43548 15416 43576 15444
rect 42751 15388 43576 15416
rect 42751 15385 42763 15388
rect 42705 15379 42763 15385
rect 39632 15320 40264 15348
rect 39632 15308 39638 15320
rect 40678 15308 40684 15360
rect 40736 15308 40742 15360
rect 40880 15348 40908 15376
rect 41506 15348 41512 15360
rect 40880 15320 41512 15348
rect 41506 15308 41512 15320
rect 41564 15308 41570 15360
rect 42628 15348 42656 15379
rect 43640 15348 43668 15444
rect 43809 15419 43867 15425
rect 43809 15385 43821 15419
rect 43855 15416 43867 15419
rect 43990 15416 43996 15428
rect 43855 15388 43996 15416
rect 43855 15385 43867 15388
rect 43809 15379 43867 15385
rect 43990 15376 43996 15388
rect 44048 15376 44054 15428
rect 42628 15320 43668 15348
rect 44085 15351 44143 15357
rect 44085 15317 44097 15351
rect 44131 15348 44143 15351
rect 44542 15348 44548 15360
rect 44131 15320 44548 15348
rect 44131 15317 44143 15320
rect 44085 15311 44143 15317
rect 44542 15308 44548 15320
rect 44600 15308 44606 15360
rect 44652 15348 44680 15456
rect 48685 15453 48697 15487
rect 48731 15453 48743 15487
rect 48685 15447 48743 15453
rect 45922 15376 45928 15428
rect 45980 15376 45986 15428
rect 47302 15416 47308 15428
rect 47150 15388 47308 15416
rect 47302 15376 47308 15388
rect 47360 15416 47366 15428
rect 47854 15416 47860 15428
rect 47360 15388 47860 15416
rect 47360 15376 47366 15388
rect 47854 15376 47860 15388
rect 47912 15376 47918 15428
rect 48700 15416 48728 15447
rect 48774 15444 48780 15496
rect 48832 15444 48838 15496
rect 49053 15487 49111 15493
rect 49053 15453 49065 15487
rect 49099 15484 49111 15487
rect 50157 15487 50215 15493
rect 50157 15484 50169 15487
rect 49099 15456 50169 15484
rect 49099 15453 49111 15456
rect 49053 15447 49111 15453
rect 50157 15453 50169 15456
rect 50203 15453 50215 15487
rect 50157 15447 50215 15453
rect 51350 15444 51356 15496
rect 51408 15444 51414 15496
rect 51552 15493 51580 15524
rect 52086 15512 52092 15564
rect 52144 15552 52150 15564
rect 52380 15552 52408 15592
rect 52454 15580 52460 15632
rect 52512 15620 52518 15632
rect 53282 15620 53288 15632
rect 52512 15592 53288 15620
rect 52512 15580 52518 15592
rect 53282 15580 53288 15592
rect 53340 15580 53346 15632
rect 53377 15623 53435 15629
rect 53377 15589 53389 15623
rect 53423 15589 53435 15623
rect 53377 15583 53435 15589
rect 53392 15552 53420 15583
rect 53929 15555 53987 15561
rect 52144 15524 52316 15552
rect 52380 15524 52500 15552
rect 52144 15512 52150 15524
rect 51537 15487 51595 15493
rect 51537 15453 51549 15487
rect 51583 15453 51595 15487
rect 51537 15447 51595 15453
rect 51718 15444 51724 15496
rect 51776 15444 51782 15496
rect 52288 15493 52316 15524
rect 52181 15487 52239 15493
rect 52181 15453 52193 15487
rect 52227 15453 52239 15487
rect 52181 15447 52239 15453
rect 52273 15487 52331 15493
rect 52273 15453 52285 15487
rect 52319 15453 52331 15487
rect 52273 15447 52331 15453
rect 48700 15388 49096 15416
rect 49068 15360 49096 15388
rect 49326 15376 49332 15428
rect 49384 15416 49390 15428
rect 51629 15419 51687 15425
rect 51629 15416 51641 15419
rect 49384 15388 51641 15416
rect 49384 15376 49390 15388
rect 51629 15385 51641 15388
rect 51675 15416 51687 15419
rect 51902 15416 51908 15428
rect 51675 15388 51908 15416
rect 51675 15385 51687 15388
rect 51629 15379 51687 15385
rect 51902 15376 51908 15388
rect 51960 15376 51966 15428
rect 46658 15348 46664 15360
rect 44652 15320 46664 15348
rect 46658 15308 46664 15320
rect 46716 15308 46722 15360
rect 47394 15308 47400 15360
rect 47452 15308 47458 15360
rect 48501 15351 48559 15357
rect 48501 15317 48513 15351
rect 48547 15348 48559 15351
rect 48682 15348 48688 15360
rect 48547 15320 48688 15348
rect 48547 15317 48559 15320
rect 48501 15311 48559 15317
rect 48682 15308 48688 15320
rect 48740 15308 48746 15360
rect 49050 15308 49056 15360
rect 49108 15308 49114 15360
rect 51718 15308 51724 15360
rect 51776 15348 51782 15360
rect 51997 15351 52055 15357
rect 51997 15348 52009 15351
rect 51776 15320 52009 15348
rect 51776 15308 51782 15320
rect 51997 15317 52009 15320
rect 52043 15317 52055 15351
rect 52196 15348 52224 15447
rect 52472 15416 52500 15524
rect 52564 15524 53144 15552
rect 53392 15524 53788 15552
rect 52564 15496 52592 15524
rect 52546 15444 52552 15496
rect 52604 15444 52610 15496
rect 52822 15444 52828 15496
rect 52880 15444 52886 15496
rect 53116 15493 53144 15524
rect 53101 15487 53159 15493
rect 53101 15453 53113 15487
rect 53147 15453 53159 15487
rect 53101 15447 53159 15453
rect 53190 15444 53196 15496
rect 53248 15444 53254 15496
rect 53558 15444 53564 15496
rect 53616 15484 53622 15496
rect 53760 15493 53788 15524
rect 53929 15521 53941 15555
rect 53975 15521 53987 15555
rect 53929 15515 53987 15521
rect 53653 15487 53711 15493
rect 53653 15484 53665 15487
rect 53616 15456 53665 15484
rect 53616 15444 53622 15456
rect 53653 15453 53665 15456
rect 53699 15453 53711 15487
rect 53653 15447 53711 15453
rect 53745 15487 53803 15493
rect 53745 15453 53757 15487
rect 53791 15453 53803 15487
rect 53745 15447 53803 15453
rect 52914 15416 52920 15428
rect 52472 15388 52920 15416
rect 52914 15376 52920 15388
rect 52972 15416 52978 15428
rect 53009 15419 53067 15425
rect 53009 15416 53021 15419
rect 52972 15388 53021 15416
rect 52972 15376 52978 15388
rect 53009 15385 53021 15388
rect 53055 15385 53067 15419
rect 53009 15379 53067 15385
rect 53282 15376 53288 15428
rect 53340 15416 53346 15428
rect 53469 15419 53527 15425
rect 53469 15416 53481 15419
rect 53340 15388 53481 15416
rect 53340 15376 53346 15388
rect 53469 15385 53481 15388
rect 53515 15385 53527 15419
rect 53944 15416 53972 15515
rect 54110 15512 54116 15564
rect 54168 15552 54174 15564
rect 55048 15561 55076 15660
rect 55861 15657 55873 15691
rect 55907 15688 55919 15691
rect 56226 15688 56232 15700
rect 55907 15660 56232 15688
rect 55907 15657 55919 15660
rect 55861 15651 55919 15657
rect 56226 15648 56232 15660
rect 56284 15648 56290 15700
rect 56594 15648 56600 15700
rect 56652 15648 56658 15700
rect 57330 15620 57336 15632
rect 55784 15592 57336 15620
rect 55033 15555 55091 15561
rect 54168 15524 54892 15552
rect 54168 15512 54174 15524
rect 54021 15487 54079 15493
rect 54021 15453 54033 15487
rect 54067 15484 54079 15487
rect 54389 15487 54447 15493
rect 54389 15484 54401 15487
rect 54067 15456 54401 15484
rect 54067 15453 54079 15456
rect 54021 15447 54079 15453
rect 54389 15453 54401 15456
rect 54435 15453 54447 15487
rect 54864 15484 54892 15524
rect 55033 15521 55045 15555
rect 55079 15552 55091 15555
rect 55079 15524 55628 15552
rect 55079 15521 55091 15524
rect 55033 15515 55091 15521
rect 55600 15493 55628 15524
rect 55309 15487 55367 15493
rect 55309 15484 55321 15487
rect 54864 15456 55321 15484
rect 54389 15447 54447 15453
rect 55309 15453 55321 15456
rect 55355 15453 55367 15487
rect 55309 15447 55367 15453
rect 55585 15487 55643 15493
rect 55585 15453 55597 15487
rect 55631 15453 55643 15487
rect 55585 15447 55643 15453
rect 53944 15388 54064 15416
rect 53469 15379 53527 15385
rect 52730 15348 52736 15360
rect 52196 15320 52736 15348
rect 51997 15311 52055 15317
rect 52730 15308 52736 15320
rect 52788 15308 52794 15360
rect 53834 15308 53840 15360
rect 53892 15348 53898 15360
rect 54036 15348 54064 15388
rect 55214 15348 55220 15360
rect 53892 15320 55220 15348
rect 53892 15308 53898 15320
rect 55214 15308 55220 15320
rect 55272 15308 55278 15360
rect 55324 15348 55352 15447
rect 55674 15444 55680 15496
rect 55732 15444 55738 15496
rect 55398 15376 55404 15428
rect 55456 15416 55462 15428
rect 55493 15419 55551 15425
rect 55493 15416 55505 15419
rect 55456 15388 55505 15416
rect 55456 15376 55462 15388
rect 55493 15385 55505 15388
rect 55539 15416 55551 15419
rect 55784 15416 55812 15592
rect 57330 15580 57336 15592
rect 57388 15580 57394 15632
rect 56042 15512 56048 15564
rect 56100 15552 56106 15564
rect 57057 15555 57115 15561
rect 57057 15552 57069 15555
rect 56100 15524 57069 15552
rect 56100 15512 56106 15524
rect 57057 15521 57069 15524
rect 57103 15521 57115 15555
rect 57057 15515 57115 15521
rect 55950 15444 55956 15496
rect 56008 15444 56014 15496
rect 56226 15444 56232 15496
rect 56284 15444 56290 15496
rect 56318 15444 56324 15496
rect 56376 15484 56382 15496
rect 56781 15487 56839 15493
rect 56781 15484 56793 15487
rect 56376 15456 56793 15484
rect 56376 15444 56382 15456
rect 56781 15453 56793 15456
rect 56827 15453 56839 15487
rect 56781 15447 56839 15453
rect 56873 15487 56931 15493
rect 56873 15453 56885 15487
rect 56919 15484 56931 15487
rect 56962 15484 56968 15496
rect 56919 15456 56968 15484
rect 56919 15453 56931 15456
rect 56873 15447 56931 15453
rect 56962 15444 56968 15456
rect 57020 15444 57026 15496
rect 57149 15487 57207 15493
rect 57149 15453 57161 15487
rect 57195 15484 57207 15487
rect 57698 15484 57704 15496
rect 57195 15456 57704 15484
rect 57195 15453 57207 15456
rect 57149 15447 57207 15453
rect 57164 15416 57192 15447
rect 57698 15444 57704 15456
rect 57756 15444 57762 15496
rect 55539 15388 55812 15416
rect 56428 15388 57192 15416
rect 55539 15385 55551 15388
rect 55493 15379 55551 15385
rect 56428 15348 56456 15388
rect 55324 15320 56456 15348
rect 56502 15308 56508 15360
rect 56560 15308 56566 15360
rect 1104 15258 58880 15280
rect 1104 15206 4874 15258
rect 4926 15206 4938 15258
rect 4990 15206 5002 15258
rect 5054 15206 5066 15258
rect 5118 15206 5130 15258
rect 5182 15206 35594 15258
rect 35646 15206 35658 15258
rect 35710 15206 35722 15258
rect 35774 15206 35786 15258
rect 35838 15206 35850 15258
rect 35902 15206 58880 15258
rect 1104 15184 58880 15206
rect 16666 15144 16672 15156
rect 13004 15116 16672 15144
rect 12618 14968 12624 15020
rect 12676 14968 12682 15020
rect 12713 15011 12771 15017
rect 12713 14977 12725 15011
rect 12759 14977 12771 15011
rect 12713 14971 12771 14977
rect 12728 14872 12756 14971
rect 12894 14968 12900 15020
rect 12952 14968 12958 15020
rect 13004 15017 13032 15116
rect 16666 15104 16672 15116
rect 16724 15104 16730 15156
rect 19613 15147 19671 15153
rect 19613 15113 19625 15147
rect 19659 15113 19671 15147
rect 19613 15107 19671 15113
rect 19705 15147 19763 15153
rect 19705 15113 19717 15147
rect 19751 15144 19763 15147
rect 20070 15144 20076 15156
rect 19751 15116 20076 15144
rect 19751 15113 19763 15116
rect 19705 15107 19763 15113
rect 13262 15036 13268 15088
rect 13320 15036 13326 15088
rect 18046 15076 18052 15088
rect 14490 15048 18052 15076
rect 18046 15036 18052 15048
rect 18104 15036 18110 15088
rect 18138 15036 18144 15088
rect 18196 15036 18202 15088
rect 19628 15076 19656 15107
rect 20070 15104 20076 15116
rect 20128 15104 20134 15156
rect 22186 15104 22192 15156
rect 22244 15104 22250 15156
rect 22370 15104 22376 15156
rect 22428 15144 22434 15156
rect 23106 15144 23112 15156
rect 22428 15116 23112 15144
rect 22428 15104 22434 15116
rect 23106 15104 23112 15116
rect 23164 15104 23170 15156
rect 23198 15104 23204 15156
rect 23256 15104 23262 15156
rect 25593 15147 25651 15153
rect 25593 15113 25605 15147
rect 25639 15144 25651 15147
rect 25682 15144 25688 15156
rect 25639 15116 25688 15144
rect 25639 15113 25651 15116
rect 25593 15107 25651 15113
rect 25682 15104 25688 15116
rect 25740 15104 25746 15156
rect 26142 15104 26148 15156
rect 26200 15144 26206 15156
rect 26329 15147 26387 15153
rect 26329 15144 26341 15147
rect 26200 15116 26341 15144
rect 26200 15104 26206 15116
rect 19978 15076 19984 15088
rect 19628 15048 19984 15076
rect 19978 15036 19984 15048
rect 20036 15036 20042 15088
rect 23216 15076 23244 15104
rect 22383 15048 23244 15076
rect 23492 15048 24854 15076
rect 12989 15011 13047 15017
rect 12989 14977 13001 15011
rect 13035 14977 13047 15011
rect 12989 14971 13047 14977
rect 14734 14968 14740 15020
rect 14792 15008 14798 15020
rect 15105 15011 15163 15017
rect 15105 15008 15117 15011
rect 14792 14980 15117 15008
rect 14792 14968 14798 14980
rect 15105 14977 15117 14980
rect 15151 14977 15163 15011
rect 15381 15011 15439 15017
rect 15381 15008 15393 15011
rect 15105 14971 15163 14977
rect 15212 14980 15393 15008
rect 13630 14900 13636 14952
rect 13688 14940 13694 14952
rect 15212 14940 15240 14980
rect 15381 14977 15393 14980
rect 15427 14977 15439 15011
rect 19274 14980 19334 15008
rect 15381 14971 15439 14977
rect 13688 14912 15240 14940
rect 15289 14943 15347 14949
rect 13688 14900 13694 14912
rect 15289 14909 15301 14943
rect 15335 14940 15347 14943
rect 15470 14940 15476 14952
rect 15335 14912 15476 14940
rect 15335 14909 15347 14912
rect 15289 14903 15347 14909
rect 15470 14900 15476 14912
rect 15528 14900 15534 14952
rect 17862 14900 17868 14952
rect 17920 14900 17926 14952
rect 12728 14844 13032 14872
rect 12342 14764 12348 14816
rect 12400 14804 12406 14816
rect 12897 14807 12955 14813
rect 12897 14804 12909 14807
rect 12400 14776 12909 14804
rect 12400 14764 12406 14776
rect 12897 14773 12909 14776
rect 12943 14773 12955 14807
rect 13004 14804 13032 14844
rect 14737 14807 14795 14813
rect 14737 14804 14749 14807
rect 13004 14776 14749 14804
rect 12897 14767 12955 14773
rect 14737 14773 14749 14776
rect 14783 14804 14795 14807
rect 14918 14804 14924 14816
rect 14783 14776 14924 14804
rect 14783 14773 14795 14776
rect 14737 14767 14795 14773
rect 14918 14764 14924 14776
rect 14976 14804 14982 14816
rect 15105 14807 15163 14813
rect 15105 14804 15117 14807
rect 14976 14776 15117 14804
rect 14976 14764 14982 14776
rect 15105 14773 15117 14776
rect 15151 14773 15163 14807
rect 15105 14767 15163 14773
rect 15565 14807 15623 14813
rect 15565 14773 15577 14807
rect 15611 14804 15623 14807
rect 16114 14804 16120 14816
rect 15611 14776 16120 14804
rect 15611 14773 15623 14776
rect 15565 14767 15623 14773
rect 16114 14764 16120 14776
rect 16172 14764 16178 14816
rect 19306 14804 19334 14980
rect 19702 14968 19708 15020
rect 19760 15008 19766 15020
rect 19843 15011 19901 15017
rect 19843 15008 19855 15011
rect 19760 14980 19855 15008
rect 19760 14968 19766 14980
rect 19843 14977 19855 14980
rect 19889 14977 19901 15011
rect 19843 14971 19901 14977
rect 20073 15011 20131 15017
rect 20073 14977 20085 15011
rect 20119 15008 20131 15011
rect 20162 15008 20168 15020
rect 20119 14980 20168 15008
rect 20119 14977 20131 14980
rect 20073 14971 20131 14977
rect 19610 14900 19616 14952
rect 19668 14940 19674 14952
rect 20088 14940 20116 14971
rect 20162 14968 20168 14980
rect 20220 14968 20226 15020
rect 20254 14968 20260 15020
rect 20312 14968 20318 15020
rect 20346 14968 20352 15020
rect 20404 14968 20410 15020
rect 20533 15011 20591 15017
rect 20533 14977 20545 15011
rect 20579 15008 20591 15011
rect 20622 15008 20628 15020
rect 20579 14980 20628 15008
rect 20579 14977 20591 14980
rect 20533 14971 20591 14977
rect 20622 14968 20628 14980
rect 20680 14968 20686 15020
rect 20901 15011 20959 15017
rect 20901 14977 20913 15011
rect 20947 15008 20959 15011
rect 21910 15008 21916 15020
rect 20947 14980 21916 15008
rect 20947 14977 20959 14980
rect 20901 14971 20959 14977
rect 21910 14968 21916 14980
rect 21968 14968 21974 15020
rect 22383 15017 22411 15048
rect 22368 15011 22426 15017
rect 22368 14977 22380 15011
rect 22414 14977 22426 15011
rect 22368 14971 22426 14977
rect 22465 15011 22523 15017
rect 22465 14977 22477 15011
rect 22511 14977 22523 15011
rect 22465 14971 22523 14977
rect 22480 14940 22508 14971
rect 22554 14968 22560 15020
rect 22612 14968 22618 15020
rect 22738 15008 22744 15020
rect 22699 14980 22744 15008
rect 22738 14968 22744 14980
rect 22796 14968 22802 15020
rect 22830 14968 22836 15020
rect 22888 14968 22894 15020
rect 23014 14968 23020 15020
rect 23072 15008 23078 15020
rect 23492 15008 23520 15048
rect 24826 15020 24854 15048
rect 25866 15036 25872 15088
rect 25924 15036 25930 15088
rect 25958 15036 25964 15088
rect 26016 15036 26022 15088
rect 23072 14980 23520 15008
rect 23569 15011 23627 15017
rect 23072 14968 23078 14980
rect 23569 14977 23581 15011
rect 23615 15008 23627 15011
rect 24118 15008 24124 15020
rect 23615 14980 24124 15008
rect 23615 14977 23627 14980
rect 23569 14971 23627 14977
rect 24118 14968 24124 14980
rect 24176 14968 24182 15020
rect 24826 14980 24860 15020
rect 24854 14968 24860 14980
rect 24912 15008 24918 15020
rect 26252 15017 26280 15116
rect 26329 15113 26341 15116
rect 26375 15113 26387 15147
rect 26329 15107 26387 15113
rect 31941 15147 31999 15153
rect 31941 15113 31953 15147
rect 31987 15144 31999 15147
rect 32122 15144 32128 15156
rect 31987 15116 32128 15144
rect 31987 15113 31999 15116
rect 31941 15107 31999 15113
rect 32122 15104 32128 15116
rect 32180 15104 32186 15156
rect 37550 15104 37556 15156
rect 37608 15144 37614 15156
rect 37737 15147 37795 15153
rect 37737 15144 37749 15147
rect 37608 15116 37749 15144
rect 37608 15104 37614 15116
rect 37737 15113 37749 15116
rect 37783 15113 37795 15147
rect 37737 15107 37795 15113
rect 38473 15147 38531 15153
rect 38473 15113 38485 15147
rect 38519 15144 38531 15147
rect 38562 15144 38568 15156
rect 38519 15116 38568 15144
rect 38519 15113 38531 15116
rect 38473 15107 38531 15113
rect 38562 15104 38568 15116
rect 38620 15144 38626 15156
rect 39482 15144 39488 15156
rect 38620 15116 39488 15144
rect 38620 15104 38626 15116
rect 39482 15104 39488 15116
rect 39540 15104 39546 15156
rect 39666 15104 39672 15156
rect 39724 15104 39730 15156
rect 42058 15144 42064 15156
rect 41386 15116 42064 15144
rect 30466 15036 30472 15088
rect 30524 15036 30530 15088
rect 30558 15036 30564 15088
rect 30616 15076 30622 15088
rect 33413 15079 33471 15085
rect 30616 15048 30958 15076
rect 30616 15036 30622 15048
rect 33413 15045 33425 15079
rect 33459 15076 33471 15079
rect 33597 15079 33655 15085
rect 33597 15076 33609 15079
rect 33459 15048 33609 15076
rect 33459 15045 33471 15048
rect 33413 15039 33471 15045
rect 33597 15045 33609 15048
rect 33643 15076 33655 15079
rect 34238 15076 34244 15088
rect 33643 15048 34244 15076
rect 33643 15045 33655 15048
rect 33597 15039 33655 15045
rect 34238 15036 34244 15048
rect 34296 15076 34302 15088
rect 41386 15076 41414 15116
rect 42058 15104 42064 15116
rect 42116 15104 42122 15156
rect 42150 15104 42156 15156
rect 42208 15144 42214 15156
rect 43070 15144 43076 15156
rect 42208 15116 43076 15144
rect 42208 15104 42214 15116
rect 43070 15104 43076 15116
rect 43128 15104 43134 15156
rect 43990 15144 43996 15156
rect 43180 15116 43996 15144
rect 34296 15048 41414 15076
rect 34296 15036 34302 15048
rect 41506 15036 41512 15088
rect 41564 15076 41570 15088
rect 43180 15076 43208 15116
rect 43990 15104 43996 15116
rect 44048 15104 44054 15156
rect 46477 15147 46535 15153
rect 46477 15113 46489 15147
rect 46523 15144 46535 15147
rect 46566 15144 46572 15156
rect 46523 15116 46572 15144
rect 46523 15113 46535 15116
rect 46477 15107 46535 15113
rect 46566 15104 46572 15116
rect 46624 15104 46630 15156
rect 49878 15104 49884 15156
rect 49936 15104 49942 15156
rect 49970 15104 49976 15156
rect 50028 15144 50034 15156
rect 51629 15147 51687 15153
rect 51629 15144 51641 15147
rect 50028 15116 51641 15144
rect 50028 15104 50034 15116
rect 51629 15113 51641 15116
rect 51675 15144 51687 15147
rect 52273 15147 52331 15153
rect 51675 15116 52040 15144
rect 51675 15113 51687 15116
rect 51629 15107 51687 15113
rect 41564 15048 43208 15076
rect 41564 15036 41570 15048
rect 25731 15011 25789 15017
rect 25731 15008 25743 15011
rect 24912 14980 25743 15008
rect 24912 14968 24918 14980
rect 25731 14977 25743 14980
rect 25777 14977 25789 15011
rect 25731 14971 25789 14977
rect 26144 15011 26202 15017
rect 26144 14977 26156 15011
rect 26190 14977 26202 15011
rect 26144 14971 26202 14977
rect 26237 15011 26295 15017
rect 26237 14977 26249 15011
rect 26283 14977 26295 15011
rect 26237 14971 26295 14977
rect 33229 15011 33287 15017
rect 33229 14977 33241 15011
rect 33275 15008 33287 15011
rect 35434 15008 35440 15020
rect 33275 14980 35440 15008
rect 33275 14977 33287 14980
rect 33229 14971 33287 14977
rect 25314 14940 25320 14952
rect 19668 14912 20116 14940
rect 22066 14912 25320 14940
rect 19668 14900 19674 14912
rect 19794 14832 19800 14884
rect 19852 14872 19858 14884
rect 22066 14872 22094 14912
rect 25314 14900 25320 14912
rect 25372 14900 25378 14952
rect 19852 14844 22094 14872
rect 19852 14832 19858 14844
rect 22738 14832 22744 14884
rect 22796 14872 22802 14884
rect 23382 14872 23388 14884
rect 22796 14844 23388 14872
rect 22796 14832 22802 14844
rect 23382 14832 23388 14844
rect 23440 14872 23446 14884
rect 26159 14872 26187 14971
rect 35434 14968 35440 14980
rect 35492 14968 35498 15020
rect 36633 15011 36691 15017
rect 36633 14977 36645 15011
rect 36679 14977 36691 15011
rect 36633 14971 36691 14977
rect 30190 14900 30196 14952
rect 30248 14900 30254 14952
rect 30926 14940 30932 14952
rect 30300 14912 30932 14940
rect 26786 14872 26792 14884
rect 23440 14844 24072 14872
rect 26159 14844 26792 14872
rect 23440 14832 23446 14844
rect 20438 14804 20444 14816
rect 19306 14776 20444 14804
rect 20438 14764 20444 14776
rect 20496 14764 20502 14816
rect 24044 14804 24072 14844
rect 26786 14832 26792 14844
rect 26844 14872 26850 14884
rect 30300 14872 30328 14912
rect 30926 14900 30932 14912
rect 30984 14900 30990 14952
rect 36648 14940 36676 14971
rect 37918 14968 37924 15020
rect 37976 14968 37982 15020
rect 38013 15011 38071 15017
rect 38013 14977 38025 15011
rect 38059 15008 38071 15011
rect 38102 15008 38108 15020
rect 38059 14980 38108 15008
rect 38059 14977 38071 14980
rect 38013 14971 38071 14977
rect 38102 14968 38108 14980
rect 38160 14968 38166 15020
rect 38289 15011 38347 15017
rect 38289 14977 38301 15011
rect 38335 15008 38347 15011
rect 38657 15011 38715 15017
rect 38657 15008 38669 15011
rect 38335 14980 38669 15008
rect 38335 14977 38347 14980
rect 38289 14971 38347 14977
rect 38657 14977 38669 14980
rect 38703 14977 38715 15011
rect 38657 14971 38715 14977
rect 39022 14968 39028 15020
rect 39080 15008 39086 15020
rect 39209 15011 39267 15017
rect 39209 15008 39221 15011
rect 39080 14980 39221 15008
rect 39080 14968 39086 14980
rect 39209 14977 39221 14980
rect 39255 14977 39267 15011
rect 39209 14971 39267 14977
rect 41230 14968 41236 15020
rect 41288 15008 41294 15020
rect 42610 15008 42616 15020
rect 41288 14980 42616 15008
rect 41288 14968 41294 14980
rect 42610 14968 42616 14980
rect 42668 15008 42674 15020
rect 42705 15011 42763 15017
rect 42705 15008 42717 15011
rect 42668 14980 42717 15008
rect 42668 14968 42674 14980
rect 42705 14977 42717 14980
rect 42751 14977 42763 15011
rect 42705 14971 42763 14977
rect 42794 14968 42800 15020
rect 42852 14968 42858 15020
rect 43073 15011 43131 15017
rect 43073 14977 43085 15011
rect 43119 15008 43131 15011
rect 43180 15008 43208 15048
rect 46014 15036 46020 15088
rect 46072 15076 46078 15088
rect 46382 15076 46388 15088
rect 46072 15048 46388 15076
rect 46072 15036 46078 15048
rect 46382 15036 46388 15048
rect 46440 15076 46446 15088
rect 46845 15079 46903 15085
rect 46845 15076 46857 15079
rect 46440 15048 46857 15076
rect 46440 15036 46446 15048
rect 46845 15045 46857 15048
rect 46891 15045 46903 15079
rect 46845 15039 46903 15045
rect 47854 15036 47860 15088
rect 47912 15076 47918 15088
rect 52012 15085 52040 15116
rect 52273 15113 52285 15147
rect 52319 15144 52331 15147
rect 52454 15144 52460 15156
rect 52319 15116 52460 15144
rect 52319 15113 52331 15116
rect 52273 15107 52331 15113
rect 52454 15104 52460 15116
rect 52512 15104 52518 15156
rect 53926 15144 53932 15156
rect 53024 15116 53932 15144
rect 51997 15079 52055 15085
rect 47912 15048 48898 15076
rect 47912 15036 47918 15048
rect 51997 15045 52009 15079
rect 52043 15045 52055 15079
rect 51997 15039 52055 15045
rect 52362 15036 52368 15088
rect 52420 15076 52426 15088
rect 52733 15079 52791 15085
rect 52733 15076 52745 15079
rect 52420 15048 52745 15076
rect 52420 15036 52426 15048
rect 52733 15045 52745 15048
rect 52779 15045 52791 15079
rect 52733 15039 52791 15045
rect 43119 14980 43208 15008
rect 43119 14977 43131 14980
rect 43073 14971 43131 14977
rect 37458 14940 37464 14952
rect 36648 14912 37464 14940
rect 37458 14900 37464 14912
rect 37516 14940 37522 14952
rect 38378 14940 38384 14952
rect 37516 14912 38384 14940
rect 37516 14900 37522 14912
rect 38378 14900 38384 14912
rect 38436 14900 38442 14952
rect 40126 14900 40132 14952
rect 40184 14940 40190 14952
rect 41414 14940 41420 14952
rect 40184 14912 41420 14940
rect 40184 14900 40190 14912
rect 41414 14900 41420 14912
rect 41472 14900 41478 14952
rect 41506 14900 41512 14952
rect 41564 14940 41570 14952
rect 43438 14940 43444 14952
rect 41564 14912 43444 14940
rect 41564 14900 41570 14912
rect 43438 14900 43444 14912
rect 43496 14940 43502 14952
rect 43548 14940 43576 14994
rect 44910 14968 44916 15020
rect 44968 14968 44974 15020
rect 46658 15017 46664 15020
rect 46656 15008 46664 15017
rect 46619 14980 46664 15008
rect 46656 14971 46664 14980
rect 46658 14968 46664 14971
rect 46716 14968 46722 15020
rect 46753 15011 46811 15017
rect 46753 14977 46765 15011
rect 46799 14977 46811 15011
rect 46753 14971 46811 14977
rect 47028 15011 47086 15017
rect 47028 14977 47040 15011
rect 47074 14977 47086 15011
rect 47028 14971 47086 14977
rect 47121 15011 47179 15017
rect 47121 14977 47133 15011
rect 47167 15008 47179 15011
rect 47210 15008 47216 15020
rect 47167 14980 47216 15008
rect 47167 14977 47179 14980
rect 47121 14971 47179 14977
rect 44174 14940 44180 14952
rect 43496 14912 43576 14940
rect 43640 14912 44180 14940
rect 43496 14900 43502 14912
rect 26844 14844 30328 14872
rect 26844 14832 26850 14844
rect 34330 14832 34336 14884
rect 34388 14872 34394 14884
rect 34609 14875 34667 14881
rect 34609 14872 34621 14875
rect 34388 14844 34621 14872
rect 34388 14832 34394 14844
rect 34609 14841 34621 14844
rect 34655 14872 34667 14875
rect 34655 14844 39712 14872
rect 34655 14841 34667 14844
rect 34609 14835 34667 14841
rect 25866 14804 25872 14816
rect 24044 14776 25872 14804
rect 25866 14764 25872 14776
rect 25924 14764 25930 14816
rect 27154 14764 27160 14816
rect 27212 14804 27218 14816
rect 34698 14804 34704 14816
rect 27212 14776 34704 14804
rect 27212 14764 27218 14776
rect 34698 14764 34704 14776
rect 34756 14804 34762 14816
rect 36446 14804 36452 14816
rect 34756 14776 36452 14804
rect 34756 14764 34762 14776
rect 36446 14764 36452 14776
rect 36504 14804 36510 14816
rect 36541 14807 36599 14813
rect 36541 14804 36553 14807
rect 36504 14776 36553 14804
rect 36504 14764 36510 14776
rect 36541 14773 36553 14776
rect 36587 14773 36599 14807
rect 36541 14767 36599 14773
rect 37826 14764 37832 14816
rect 37884 14804 37890 14816
rect 38194 14804 38200 14816
rect 37884 14776 38200 14804
rect 37884 14764 37890 14776
rect 38194 14764 38200 14776
rect 38252 14764 38258 14816
rect 39684 14804 39712 14844
rect 40034 14832 40040 14884
rect 40092 14872 40098 14884
rect 40954 14872 40960 14884
rect 40092 14844 40960 14872
rect 40092 14832 40098 14844
rect 40954 14832 40960 14844
rect 41012 14872 41018 14884
rect 42150 14872 42156 14884
rect 41012 14844 42156 14872
rect 41012 14832 41018 14844
rect 42150 14832 42156 14844
rect 42208 14832 42214 14884
rect 42334 14832 42340 14884
rect 42392 14872 42398 14884
rect 43165 14875 43223 14881
rect 43165 14872 43177 14875
rect 42392 14844 43177 14872
rect 42392 14832 42398 14844
rect 43165 14841 43177 14844
rect 43211 14841 43223 14875
rect 43165 14835 43223 14841
rect 42426 14804 42432 14816
rect 39684 14776 42432 14804
rect 42426 14764 42432 14776
rect 42484 14764 42490 14816
rect 42521 14807 42579 14813
rect 42521 14773 42533 14807
rect 42567 14804 42579 14807
rect 42702 14804 42708 14816
rect 42567 14776 42708 14804
rect 42567 14773 42579 14776
rect 42521 14767 42579 14773
rect 42702 14764 42708 14776
rect 42760 14764 42766 14816
rect 42981 14807 43039 14813
rect 42981 14773 42993 14807
rect 43027 14804 43039 14807
rect 43070 14804 43076 14816
rect 43027 14776 43076 14804
rect 43027 14773 43039 14776
rect 42981 14767 43039 14773
rect 43070 14764 43076 14776
rect 43128 14764 43134 14816
rect 43180 14804 43208 14835
rect 43254 14832 43260 14884
rect 43312 14872 43318 14884
rect 43640 14872 43668 14912
rect 44174 14900 44180 14912
rect 44232 14900 44238 14952
rect 44266 14900 44272 14952
rect 44324 14940 44330 14952
rect 44637 14943 44695 14949
rect 44637 14940 44649 14943
rect 44324 14912 44649 14940
rect 44324 14900 44330 14912
rect 44637 14909 44649 14912
rect 44683 14909 44695 14943
rect 46768 14940 46796 14971
rect 47044 14940 47072 14971
rect 47210 14968 47216 14980
rect 47268 14968 47274 15020
rect 47946 14968 47952 15020
rect 48004 15008 48010 15020
rect 48133 15011 48191 15017
rect 48133 15008 48145 15011
rect 48004 14980 48145 15008
rect 48004 14968 48010 14980
rect 48133 14977 48145 14980
rect 48179 14977 48191 15011
rect 48133 14971 48191 14977
rect 51810 14968 51816 15020
rect 51868 14968 51874 15020
rect 53024 14952 53052 15116
rect 53926 15104 53932 15116
rect 53984 15144 53990 15156
rect 55122 15144 55128 15156
rect 53984 15116 55128 15144
rect 53984 15104 53990 15116
rect 55122 15104 55128 15116
rect 55180 15144 55186 15156
rect 55180 15116 56732 15144
rect 55180 15104 55186 15116
rect 53282 15036 53288 15088
rect 53340 15036 53346 15088
rect 53742 15036 53748 15088
rect 53800 15036 53806 15088
rect 56413 15079 56471 15085
rect 56413 15045 56425 15079
rect 56459 15076 56471 15079
rect 56502 15076 56508 15088
rect 56459 15048 56508 15076
rect 56459 15045 56471 15048
rect 56413 15039 56471 15045
rect 56502 15036 56508 15048
rect 56560 15036 56566 15088
rect 56704 15017 56732 15116
rect 56689 15011 56747 15017
rect 54680 14980 55338 15008
rect 49694 14940 49700 14952
rect 46768 14912 46888 14940
rect 47044 14912 49700 14940
rect 44637 14903 44695 14909
rect 43312 14844 43668 14872
rect 46860 14872 46888 14912
rect 49694 14900 49700 14912
rect 49752 14900 49758 14952
rect 50062 14900 50068 14952
rect 50120 14940 50126 14952
rect 52546 14940 52552 14952
rect 50120 14912 52552 14940
rect 50120 14900 50126 14912
rect 52546 14900 52552 14912
rect 52604 14900 52610 14952
rect 53006 14900 53012 14952
rect 53064 14900 53070 14952
rect 53742 14900 53748 14952
rect 53800 14940 53806 14952
rect 54680 14940 54708 14980
rect 56689 14977 56701 15011
rect 56735 14977 56747 15011
rect 56689 14971 56747 14977
rect 53800 14912 54708 14940
rect 53800 14900 53806 14912
rect 46860 14844 48268 14872
rect 43312 14832 43318 14844
rect 48240 14816 48268 14844
rect 44082 14804 44088 14816
rect 43180 14776 44088 14804
rect 44082 14764 44088 14776
rect 44140 14804 44146 14816
rect 44634 14804 44640 14816
rect 44140 14776 44640 14804
rect 44140 14764 44146 14776
rect 44634 14764 44640 14776
rect 44692 14764 44698 14816
rect 45094 14764 45100 14816
rect 45152 14804 45158 14816
rect 47118 14804 47124 14816
rect 45152 14776 47124 14804
rect 45152 14764 45158 14776
rect 47118 14764 47124 14776
rect 47176 14764 47182 14816
rect 47210 14764 47216 14816
rect 47268 14764 47274 14816
rect 48222 14764 48228 14816
rect 48280 14764 48286 14816
rect 48407 14813 48413 14816
rect 48396 14807 48413 14813
rect 48396 14773 48408 14807
rect 48396 14767 48413 14773
rect 48407 14764 48413 14767
rect 48465 14764 48471 14816
rect 54680 14804 54708 14912
rect 54754 14900 54760 14952
rect 54812 14900 54818 14952
rect 54941 14943 54999 14949
rect 54941 14909 54953 14943
rect 54987 14940 54999 14943
rect 55030 14940 55036 14952
rect 54987 14912 55036 14940
rect 54987 14909 54999 14912
rect 54941 14903 54999 14909
rect 55030 14900 55036 14912
rect 55088 14940 55094 14952
rect 55950 14940 55956 14952
rect 55088 14912 55956 14940
rect 55088 14900 55094 14912
rect 55950 14900 55956 14912
rect 56008 14900 56014 14952
rect 56686 14804 56692 14816
rect 54680 14776 56692 14804
rect 56686 14764 56692 14776
rect 56744 14764 56750 14816
rect 1104 14714 58880 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 58880 14714
rect 1104 14640 58880 14662
rect 12894 14560 12900 14612
rect 12952 14600 12958 14612
rect 13265 14603 13323 14609
rect 13265 14600 13277 14603
rect 12952 14572 13277 14600
rect 12952 14560 12958 14572
rect 13265 14569 13277 14572
rect 13311 14569 13323 14603
rect 13265 14563 13323 14569
rect 19245 14603 19303 14609
rect 19245 14569 19257 14603
rect 19291 14600 19303 14603
rect 19702 14600 19708 14612
rect 19291 14572 19708 14600
rect 19291 14569 19303 14572
rect 19245 14563 19303 14569
rect 19702 14560 19708 14572
rect 19760 14560 19766 14612
rect 20254 14560 20260 14612
rect 20312 14600 20318 14612
rect 20312 14572 22876 14600
rect 20312 14560 20318 14572
rect 22848 14532 22876 14572
rect 22922 14560 22928 14612
rect 22980 14600 22986 14612
rect 23293 14603 23351 14609
rect 23293 14600 23305 14603
rect 22980 14572 23305 14600
rect 22980 14560 22986 14572
rect 23293 14569 23305 14572
rect 23339 14569 23351 14603
rect 23293 14563 23351 14569
rect 24489 14603 24547 14609
rect 24489 14569 24501 14603
rect 24535 14569 24547 14603
rect 24489 14563 24547 14569
rect 22848 14504 23060 14532
rect 12710 14464 12716 14476
rect 12176 14436 12716 14464
rect 1210 14356 1216 14408
rect 1268 14396 1274 14408
rect 12176 14405 12204 14436
rect 12710 14424 12716 14436
rect 12768 14424 12774 14476
rect 12989 14467 13047 14473
rect 12989 14433 13001 14467
rect 13035 14464 13047 14467
rect 13170 14464 13176 14476
rect 13035 14436 13176 14464
rect 13035 14433 13047 14436
rect 12989 14427 13047 14433
rect 13170 14424 13176 14436
rect 13228 14424 13234 14476
rect 13446 14424 13452 14476
rect 13504 14464 13510 14476
rect 13817 14467 13875 14473
rect 13817 14464 13829 14467
rect 13504 14436 13829 14464
rect 13504 14424 13510 14436
rect 13817 14433 13829 14436
rect 13863 14433 13875 14467
rect 13817 14427 13875 14433
rect 14734 14424 14740 14476
rect 14792 14424 14798 14476
rect 15105 14467 15163 14473
rect 15105 14433 15117 14467
rect 15151 14464 15163 14467
rect 15194 14464 15200 14476
rect 15151 14436 15200 14464
rect 15151 14433 15163 14436
rect 15105 14427 15163 14433
rect 15194 14424 15200 14436
rect 15252 14424 15258 14476
rect 15381 14467 15439 14473
rect 15381 14433 15393 14467
rect 15427 14464 15439 14467
rect 16945 14467 17003 14473
rect 16945 14464 16957 14467
rect 15427 14436 16957 14464
rect 15427 14433 15439 14436
rect 15381 14427 15439 14433
rect 16945 14433 16957 14436
rect 16991 14433 17003 14467
rect 16945 14427 17003 14433
rect 17221 14467 17279 14473
rect 17221 14433 17233 14467
rect 17267 14464 17279 14467
rect 17310 14464 17316 14476
rect 17267 14436 17316 14464
rect 17267 14433 17279 14436
rect 17221 14427 17279 14433
rect 17310 14424 17316 14436
rect 17368 14464 17374 14476
rect 17862 14464 17868 14476
rect 17368 14436 17868 14464
rect 17368 14424 17374 14436
rect 17862 14424 17868 14436
rect 17920 14424 17926 14476
rect 18046 14424 18052 14476
rect 18104 14464 18110 14476
rect 20622 14464 20628 14476
rect 18104 14436 20628 14464
rect 18104 14424 18110 14436
rect 20622 14424 20628 14436
rect 20680 14424 20686 14476
rect 20714 14424 20720 14476
rect 20772 14424 20778 14476
rect 21726 14424 21732 14476
rect 21784 14424 21790 14476
rect 1397 14399 1455 14405
rect 1397 14396 1409 14399
rect 1268 14368 1409 14396
rect 1268 14356 1274 14368
rect 1397 14365 1409 14368
rect 1443 14396 1455 14399
rect 1673 14399 1731 14405
rect 1673 14396 1685 14399
rect 1443 14368 1685 14396
rect 1443 14365 1455 14368
rect 1397 14359 1455 14365
rect 1673 14365 1685 14368
rect 1719 14365 1731 14399
rect 1673 14359 1731 14365
rect 12161 14399 12219 14405
rect 12161 14365 12173 14399
rect 12207 14365 12219 14399
rect 12161 14359 12219 14365
rect 12342 14356 12348 14408
rect 12400 14356 12406 14408
rect 12621 14399 12679 14405
rect 12621 14365 12633 14399
rect 12667 14365 12679 14399
rect 12621 14359 12679 14365
rect 15013 14399 15071 14405
rect 15013 14365 15025 14399
rect 15059 14396 15071 14399
rect 15286 14396 15292 14408
rect 15059 14368 15292 14396
rect 15059 14365 15071 14368
rect 15013 14359 15071 14365
rect 11698 14328 11704 14340
rect 1596 14300 11704 14328
rect 1596 14269 1624 14300
rect 11698 14288 11704 14300
rect 11756 14288 11762 14340
rect 12636 14328 12664 14359
rect 15286 14356 15292 14368
rect 15344 14356 15350 14408
rect 20993 14399 21051 14405
rect 20993 14365 21005 14399
rect 21039 14396 21051 14399
rect 21450 14396 21456 14408
rect 21039 14368 21456 14396
rect 21039 14365 21051 14368
rect 20993 14359 21051 14365
rect 21450 14356 21456 14368
rect 21508 14356 21514 14408
rect 14093 14331 14151 14337
rect 14093 14328 14105 14331
rect 12636 14300 14105 14328
rect 14093 14297 14105 14300
rect 14139 14297 14151 14331
rect 17954 14328 17960 14340
rect 16514 14300 17960 14328
rect 14093 14291 14151 14297
rect 16776 14272 16804 14300
rect 17954 14288 17960 14300
rect 18012 14288 18018 14340
rect 18509 14331 18567 14337
rect 18509 14297 18521 14331
rect 18555 14328 18567 14331
rect 18877 14331 18935 14337
rect 18877 14328 18889 14331
rect 18555 14300 18889 14328
rect 18555 14297 18567 14300
rect 18509 14291 18567 14297
rect 18877 14297 18889 14300
rect 18923 14328 18935 14331
rect 19426 14328 19432 14340
rect 18923 14300 19432 14328
rect 18923 14297 18935 14300
rect 18877 14291 18935 14297
rect 19426 14288 19432 14300
rect 19484 14288 19490 14340
rect 20438 14328 20444 14340
rect 20286 14300 20444 14328
rect 20438 14288 20444 14300
rect 20496 14328 20502 14340
rect 22002 14328 22008 14340
rect 20496 14300 22008 14328
rect 20496 14288 20502 14300
rect 22002 14288 22008 14300
rect 22060 14328 22066 14340
rect 22186 14328 22192 14340
rect 22060 14300 22192 14328
rect 22060 14288 22066 14300
rect 22186 14288 22192 14300
rect 22244 14288 22250 14340
rect 23032 14328 23060 14504
rect 23106 14492 23112 14544
rect 23164 14532 23170 14544
rect 24504 14532 24532 14563
rect 24762 14560 24768 14612
rect 24820 14560 24826 14612
rect 25240 14572 26464 14600
rect 23164 14504 24532 14532
rect 23164 14492 23170 14504
rect 24780 14464 24808 14560
rect 23860 14436 24808 14464
rect 23198 14356 23204 14408
rect 23256 14396 23262 14408
rect 23431 14399 23489 14405
rect 23431 14396 23443 14399
rect 23256 14368 23443 14396
rect 23256 14356 23262 14368
rect 23431 14365 23443 14368
rect 23477 14365 23489 14399
rect 23431 14359 23489 14365
rect 23566 14356 23572 14408
rect 23624 14356 23630 14408
rect 23860 14405 23888 14436
rect 23844 14399 23902 14405
rect 23844 14365 23856 14399
rect 23890 14365 23902 14399
rect 23844 14359 23902 14365
rect 23937 14399 23995 14405
rect 23937 14365 23949 14399
rect 23983 14365 23995 14399
rect 23937 14359 23995 14365
rect 23584 14328 23612 14356
rect 23032 14300 23612 14328
rect 23661 14331 23719 14337
rect 1581 14263 1639 14269
rect 1581 14229 1593 14263
rect 1627 14229 1639 14263
rect 1581 14223 1639 14229
rect 12250 14220 12256 14272
rect 12308 14220 12314 14272
rect 15470 14220 15476 14272
rect 15528 14220 15534 14272
rect 16758 14220 16764 14272
rect 16816 14220 16822 14272
rect 18138 14220 18144 14272
rect 18196 14260 18202 14272
rect 18693 14263 18751 14269
rect 18693 14260 18705 14263
rect 18196 14232 18705 14260
rect 18196 14220 18202 14232
rect 18693 14229 18705 14232
rect 18739 14260 18751 14263
rect 18969 14263 19027 14269
rect 18969 14260 18981 14263
rect 18739 14232 18981 14260
rect 18739 14229 18751 14232
rect 18693 14223 18751 14229
rect 18969 14229 18981 14232
rect 19015 14260 19027 14263
rect 19150 14260 19156 14272
rect 19015 14232 19156 14260
rect 19015 14229 19027 14232
rect 18969 14223 19027 14229
rect 19150 14220 19156 14232
rect 19208 14260 19214 14272
rect 19886 14260 19892 14272
rect 19208 14232 19892 14260
rect 19208 14220 19214 14232
rect 19886 14220 19892 14232
rect 19944 14220 19950 14272
rect 23216 14269 23244 14300
rect 23661 14297 23673 14331
rect 23707 14297 23719 14331
rect 23661 14291 23719 14297
rect 23201 14263 23259 14269
rect 23201 14229 23213 14263
rect 23247 14229 23259 14263
rect 23201 14223 23259 14229
rect 23474 14220 23480 14272
rect 23532 14260 23538 14272
rect 23676 14260 23704 14291
rect 23750 14288 23756 14340
rect 23808 14328 23814 14340
rect 23952 14328 23980 14359
rect 24210 14356 24216 14408
rect 24268 14356 24274 14408
rect 24670 14356 24676 14408
rect 24728 14356 24734 14408
rect 25240 14396 25268 14572
rect 26436 14532 26464 14572
rect 26694 14560 26700 14612
rect 26752 14560 26758 14612
rect 28350 14600 28356 14612
rect 27724 14572 28356 14600
rect 27724 14532 27752 14572
rect 28350 14560 28356 14572
rect 28408 14600 28414 14612
rect 30282 14600 30288 14612
rect 28408 14572 30288 14600
rect 28408 14560 28414 14572
rect 30282 14560 30288 14572
rect 30340 14560 30346 14612
rect 34330 14560 34336 14612
rect 34388 14560 34394 14612
rect 34747 14603 34805 14609
rect 34747 14569 34759 14603
rect 34793 14600 34805 14603
rect 35986 14600 35992 14612
rect 34793 14572 35992 14600
rect 34793 14569 34805 14572
rect 34747 14563 34805 14569
rect 35986 14560 35992 14572
rect 36044 14600 36050 14612
rect 36262 14600 36268 14612
rect 36044 14572 36268 14600
rect 36044 14560 36050 14572
rect 36262 14560 36268 14572
rect 36320 14560 36326 14612
rect 36906 14560 36912 14612
rect 36964 14600 36970 14612
rect 37093 14603 37151 14609
rect 37093 14600 37105 14603
rect 36964 14572 37105 14600
rect 36964 14560 36970 14572
rect 37093 14569 37105 14572
rect 37139 14569 37151 14603
rect 37093 14563 37151 14569
rect 38194 14560 38200 14612
rect 38252 14600 38258 14612
rect 41322 14600 41328 14612
rect 38252 14572 41328 14600
rect 38252 14560 38258 14572
rect 41322 14560 41328 14572
rect 41380 14600 41386 14612
rect 41380 14572 42472 14600
rect 41380 14560 41386 14572
rect 26436 14504 27752 14532
rect 30006 14492 30012 14544
rect 30064 14532 30070 14544
rect 30742 14532 30748 14544
rect 30064 14504 30748 14532
rect 30064 14492 30070 14504
rect 30742 14492 30748 14504
rect 30800 14492 30806 14544
rect 30926 14492 30932 14544
rect 30984 14532 30990 14544
rect 31662 14532 31668 14544
rect 30984 14504 31668 14532
rect 30984 14492 30990 14504
rect 31662 14492 31668 14504
rect 31720 14532 31726 14544
rect 31720 14504 32720 14532
rect 31720 14492 31726 14504
rect 26234 14424 26240 14476
rect 26292 14424 26298 14476
rect 26513 14467 26571 14473
rect 26513 14433 26525 14467
rect 26559 14464 26571 14467
rect 26970 14464 26976 14476
rect 26559 14436 26976 14464
rect 26559 14433 26571 14436
rect 26513 14427 26571 14433
rect 26970 14424 26976 14436
rect 27028 14424 27034 14476
rect 27062 14424 27068 14476
rect 27120 14464 27126 14476
rect 27341 14467 27399 14473
rect 27341 14464 27353 14467
rect 27120 14436 27353 14464
rect 27120 14424 27126 14436
rect 27341 14433 27353 14436
rect 27387 14433 27399 14467
rect 27341 14427 27399 14433
rect 28626 14424 28632 14476
rect 28684 14464 28690 14476
rect 29365 14467 29423 14473
rect 29365 14464 29377 14467
rect 28684 14436 29377 14464
rect 28684 14424 28690 14436
rect 29365 14433 29377 14436
rect 29411 14464 29423 14467
rect 30190 14464 30196 14476
rect 29411 14436 30196 14464
rect 29411 14433 29423 14436
rect 29365 14427 29423 14433
rect 30190 14424 30196 14436
rect 30248 14464 30254 14476
rect 32582 14464 32588 14476
rect 30248 14436 32588 14464
rect 30248 14424 30254 14436
rect 32582 14424 32588 14436
rect 32640 14424 32646 14476
rect 32692 14464 32720 14504
rect 36814 14492 36820 14544
rect 36872 14492 36878 14544
rect 41248 14504 42380 14532
rect 34698 14464 34704 14476
rect 32692 14436 34704 14464
rect 34698 14424 34704 14436
rect 34756 14464 34762 14476
rect 35250 14464 35256 14476
rect 34756 14436 35256 14464
rect 34756 14424 34762 14436
rect 35250 14424 35256 14436
rect 35308 14424 35314 14476
rect 36541 14467 36599 14473
rect 36541 14433 36553 14467
rect 36587 14464 36599 14467
rect 37274 14464 37280 14476
rect 36587 14436 37280 14464
rect 36587 14433 36599 14436
rect 36541 14427 36599 14433
rect 37274 14424 37280 14436
rect 37332 14424 37338 14476
rect 40402 14424 40408 14476
rect 40460 14464 40466 14476
rect 40589 14467 40647 14473
rect 40589 14464 40601 14467
rect 40460 14436 40601 14464
rect 40460 14424 40466 14436
rect 40589 14433 40601 14436
rect 40635 14464 40647 14467
rect 40635 14436 41092 14464
rect 40635 14433 40647 14436
rect 40589 14427 40647 14433
rect 24780 14368 25268 14396
rect 26881 14399 26939 14405
rect 23808 14300 23980 14328
rect 24228 14328 24256 14356
rect 24780 14328 24808 14368
rect 26881 14365 26893 14399
rect 26927 14396 26939 14399
rect 27092 14396 27120 14424
rect 26927 14368 27120 14396
rect 26927 14365 26939 14368
rect 26881 14359 26939 14365
rect 27154 14356 27160 14408
rect 27212 14356 27218 14408
rect 29733 14399 29791 14405
rect 29733 14365 29745 14399
rect 29779 14365 29791 14399
rect 29733 14359 29791 14365
rect 24228 14300 24808 14328
rect 23808 14288 23814 14300
rect 25958 14288 25964 14340
rect 26016 14328 26022 14340
rect 26326 14328 26332 14340
rect 26016 14300 26332 14328
rect 26016 14288 26022 14300
rect 26326 14288 26332 14300
rect 26384 14328 26390 14340
rect 26973 14331 27031 14337
rect 26973 14328 26985 14331
rect 26384 14300 26985 14328
rect 26384 14288 26390 14300
rect 26973 14297 26985 14300
rect 27019 14297 27031 14331
rect 26973 14291 27031 14297
rect 28350 14288 28356 14340
rect 28408 14288 28414 14340
rect 29089 14331 29147 14337
rect 29089 14297 29101 14331
rect 29135 14297 29147 14331
rect 29748 14328 29776 14359
rect 29822 14356 29828 14408
rect 29880 14356 29886 14408
rect 29914 14356 29920 14408
rect 29972 14356 29978 14408
rect 30009 14399 30067 14405
rect 30009 14365 30021 14399
rect 30055 14396 30067 14399
rect 30745 14399 30803 14405
rect 30745 14396 30757 14399
rect 30055 14368 30757 14396
rect 30055 14365 30067 14368
rect 30009 14359 30067 14365
rect 30745 14365 30757 14368
rect 30791 14365 30803 14399
rect 30745 14359 30803 14365
rect 30926 14356 30932 14408
rect 30984 14356 30990 14408
rect 31021 14399 31079 14405
rect 31021 14365 31033 14399
rect 31067 14365 31079 14399
rect 33994 14368 35388 14396
rect 31021 14359 31079 14365
rect 29748 14300 30052 14328
rect 29089 14291 29147 14297
rect 23532 14232 23704 14260
rect 24213 14263 24271 14269
rect 23532 14220 23538 14232
rect 24213 14229 24225 14263
rect 24259 14260 24271 14263
rect 24302 14260 24308 14272
rect 24259 14232 24308 14260
rect 24259 14229 24271 14232
rect 24213 14223 24271 14229
rect 24302 14220 24308 14232
rect 24360 14260 24366 14272
rect 26142 14260 26148 14272
rect 24360 14232 26148 14260
rect 24360 14220 24366 14232
rect 26142 14220 26148 14232
rect 26200 14220 26206 14272
rect 26510 14220 26516 14272
rect 26568 14260 26574 14272
rect 27617 14263 27675 14269
rect 27617 14260 27629 14263
rect 26568 14232 27629 14260
rect 26568 14220 26574 14232
rect 27617 14229 27629 14232
rect 27663 14229 27675 14263
rect 29104 14260 29132 14291
rect 30024 14272 30052 14300
rect 30282 14288 30288 14340
rect 30340 14288 30346 14340
rect 30466 14288 30472 14340
rect 30524 14328 30530 14340
rect 31036 14328 31064 14359
rect 35360 14340 35388 14368
rect 36170 14356 36176 14408
rect 36228 14356 36234 14408
rect 36446 14356 36452 14408
rect 36504 14396 36510 14408
rect 36633 14399 36691 14405
rect 36633 14396 36645 14399
rect 36504 14368 36645 14396
rect 36504 14356 36510 14368
rect 36633 14365 36645 14368
rect 36679 14365 36691 14399
rect 36633 14359 36691 14365
rect 36814 14356 36820 14408
rect 36872 14396 36878 14408
rect 37001 14399 37059 14405
rect 37001 14396 37013 14399
rect 36872 14368 37013 14396
rect 36872 14356 36878 14368
rect 37001 14365 37013 14368
rect 37047 14365 37059 14399
rect 37001 14359 37059 14365
rect 37185 14399 37243 14405
rect 37185 14365 37197 14399
rect 37231 14365 37243 14399
rect 37185 14359 37243 14365
rect 30524 14300 31064 14328
rect 30524 14288 30530 14300
rect 32858 14288 32864 14340
rect 32916 14288 32922 14340
rect 35342 14288 35348 14340
rect 35400 14288 35406 14340
rect 36906 14288 36912 14340
rect 36964 14328 36970 14340
rect 37200 14328 37228 14359
rect 40126 14356 40132 14408
rect 40184 14396 40190 14408
rect 40773 14399 40831 14405
rect 40773 14396 40785 14399
rect 40184 14368 40785 14396
rect 40184 14356 40190 14368
rect 40773 14365 40785 14368
rect 40819 14365 40831 14399
rect 40773 14359 40831 14365
rect 40954 14356 40960 14408
rect 41012 14356 41018 14408
rect 41064 14405 41092 14436
rect 41049 14399 41107 14405
rect 41049 14365 41061 14399
rect 41095 14365 41107 14399
rect 41049 14359 41107 14365
rect 41138 14356 41144 14408
rect 41196 14356 41202 14408
rect 36964 14300 37228 14328
rect 41248 14328 41276 14504
rect 41322 14424 41328 14476
rect 41380 14464 41386 14476
rect 41380 14424 41414 14464
rect 41386 14396 41414 14424
rect 42352 14405 42380 14504
rect 42444 14464 42472 14572
rect 42518 14560 42524 14612
rect 42576 14560 42582 14612
rect 42794 14560 42800 14612
rect 42852 14600 42858 14612
rect 43717 14603 43775 14609
rect 43717 14600 43729 14603
rect 42852 14572 43729 14600
rect 42852 14560 42858 14572
rect 43717 14569 43729 14572
rect 43763 14569 43775 14603
rect 43717 14563 43775 14569
rect 43806 14560 43812 14612
rect 43864 14600 43870 14612
rect 47026 14600 47032 14612
rect 43864 14572 47032 14600
rect 43864 14560 43870 14572
rect 47026 14560 47032 14572
rect 47084 14600 47090 14612
rect 47305 14603 47363 14609
rect 47305 14600 47317 14603
rect 47084 14572 47317 14600
rect 47084 14560 47090 14572
rect 47305 14569 47317 14572
rect 47351 14569 47363 14603
rect 47305 14563 47363 14569
rect 48409 14603 48467 14609
rect 48409 14569 48421 14603
rect 48455 14600 48467 14603
rect 48774 14600 48780 14612
rect 48455 14572 48780 14600
rect 48455 14569 48467 14572
rect 48409 14563 48467 14569
rect 48774 14560 48780 14572
rect 48832 14560 48838 14612
rect 49234 14560 49240 14612
rect 49292 14600 49298 14612
rect 51258 14600 51264 14612
rect 49292 14572 51264 14600
rect 49292 14560 49298 14572
rect 51258 14560 51264 14572
rect 51316 14600 51322 14612
rect 51810 14600 51816 14612
rect 51316 14572 51816 14600
rect 51316 14560 51322 14572
rect 51810 14560 51816 14572
rect 51868 14560 51874 14612
rect 42536 14532 42564 14560
rect 44450 14532 44456 14544
rect 42536 14504 43668 14532
rect 42521 14467 42579 14473
rect 42521 14464 42533 14467
rect 42444 14436 42533 14464
rect 42521 14433 42533 14436
rect 42567 14464 42579 14467
rect 43070 14464 43076 14476
rect 42567 14436 43076 14464
rect 42567 14433 42579 14436
rect 42521 14427 42579 14433
rect 43070 14424 43076 14436
rect 43128 14424 43134 14476
rect 43640 14473 43668 14504
rect 44008 14504 44456 14532
rect 43625 14467 43683 14473
rect 43625 14433 43637 14467
rect 43671 14433 43683 14467
rect 43625 14427 43683 14433
rect 41509 14399 41567 14405
rect 41509 14396 41521 14399
rect 41386 14368 41521 14396
rect 41509 14365 41521 14368
rect 41555 14365 41567 14399
rect 41509 14359 41567 14365
rect 42245 14399 42303 14405
rect 42245 14365 42257 14399
rect 42291 14365 42303 14399
rect 42245 14359 42303 14365
rect 42337 14399 42395 14405
rect 42337 14365 42349 14399
rect 42383 14365 42395 14399
rect 42337 14359 42395 14365
rect 41248 14300 41368 14328
rect 36964 14288 36970 14300
rect 29549 14263 29607 14269
rect 29549 14260 29561 14263
rect 29104 14232 29561 14260
rect 27617 14223 27675 14229
rect 29549 14229 29561 14232
rect 29595 14229 29607 14263
rect 29549 14223 29607 14229
rect 30006 14220 30012 14272
rect 30064 14220 30070 14272
rect 30374 14220 30380 14272
rect 30432 14260 30438 14272
rect 30558 14260 30564 14272
rect 30432 14232 30564 14260
rect 30432 14220 30438 14232
rect 30558 14220 30564 14232
rect 30616 14220 30622 14272
rect 35250 14220 35256 14272
rect 35308 14260 35314 14272
rect 38470 14260 38476 14272
rect 35308 14232 38476 14260
rect 35308 14220 35314 14232
rect 38470 14220 38476 14232
rect 38528 14220 38534 14272
rect 40037 14263 40095 14269
rect 40037 14229 40049 14263
rect 40083 14260 40095 14263
rect 40126 14260 40132 14272
rect 40083 14232 40132 14260
rect 40083 14229 40095 14232
rect 40037 14223 40095 14229
rect 40126 14220 40132 14232
rect 40184 14220 40190 14272
rect 41340 14269 41368 14300
rect 41325 14263 41383 14269
rect 41325 14229 41337 14263
rect 41371 14229 41383 14263
rect 41325 14223 41383 14229
rect 42058 14220 42064 14272
rect 42116 14220 42122 14272
rect 42260 14260 42288 14359
rect 42426 14356 42432 14408
rect 42484 14396 42490 14408
rect 42613 14399 42671 14405
rect 42613 14396 42625 14399
rect 42484 14368 42625 14396
rect 42484 14356 42490 14368
rect 42613 14365 42625 14368
rect 42659 14365 42671 14399
rect 42613 14359 42671 14365
rect 42628 14328 42656 14359
rect 43346 14356 43352 14408
rect 43404 14396 43410 14408
rect 43901 14399 43959 14405
rect 43901 14396 43913 14399
rect 43404 14368 43913 14396
rect 43404 14356 43410 14368
rect 43901 14365 43913 14368
rect 43947 14396 43959 14399
rect 44008 14396 44036 14504
rect 44450 14492 44456 14504
rect 44508 14492 44514 14544
rect 48958 14492 48964 14544
rect 49016 14532 49022 14544
rect 49016 14504 50568 14532
rect 49016 14492 49022 14504
rect 44082 14424 44088 14476
rect 44140 14424 44146 14476
rect 46014 14424 46020 14476
rect 46072 14464 46078 14476
rect 48222 14464 48228 14476
rect 46072 14436 48228 14464
rect 46072 14424 46078 14436
rect 48222 14424 48228 14436
rect 48280 14424 48286 14476
rect 49786 14464 49792 14476
rect 48608 14436 49792 14464
rect 43947 14368 44036 14396
rect 44100 14396 44128 14424
rect 44269 14399 44327 14405
rect 44269 14396 44281 14399
rect 44100 14368 44281 14396
rect 43947 14365 43959 14368
rect 43901 14359 43959 14365
rect 44269 14365 44281 14368
rect 44315 14365 44327 14399
rect 44269 14359 44327 14365
rect 46566 14356 46572 14408
rect 46624 14356 46630 14408
rect 46750 14356 46756 14408
rect 46808 14356 46814 14408
rect 46845 14399 46903 14405
rect 46845 14365 46857 14399
rect 46891 14396 46903 14399
rect 47578 14396 47584 14408
rect 46891 14368 47584 14396
rect 46891 14365 46903 14368
rect 46845 14359 46903 14365
rect 47578 14356 47584 14368
rect 47636 14356 47642 14408
rect 48608 14405 48636 14436
rect 48593 14399 48651 14405
rect 48593 14365 48605 14399
rect 48639 14365 48651 14399
rect 48593 14359 48651 14365
rect 48774 14356 48780 14408
rect 48832 14356 48838 14408
rect 48958 14356 48964 14408
rect 49016 14356 49022 14408
rect 49252 14405 49280 14436
rect 49786 14424 49792 14436
rect 49844 14424 49850 14476
rect 50540 14408 50568 14504
rect 51445 14467 51503 14473
rect 51445 14433 51457 14467
rect 51491 14464 51503 14467
rect 53006 14464 53012 14476
rect 51491 14436 53012 14464
rect 51491 14433 51503 14436
rect 51445 14427 51503 14433
rect 53006 14424 53012 14436
rect 53064 14424 53070 14476
rect 49237 14399 49295 14405
rect 49237 14365 49249 14399
rect 49283 14365 49295 14399
rect 49237 14359 49295 14365
rect 49329 14399 49387 14405
rect 49329 14365 49341 14399
rect 49375 14365 49387 14399
rect 49329 14359 49387 14365
rect 49421 14399 49479 14405
rect 49421 14365 49433 14399
rect 49467 14396 49479 14399
rect 49467 14368 49556 14396
rect 49467 14365 49479 14368
rect 49421 14359 49479 14365
rect 43993 14331 44051 14337
rect 43993 14328 44005 14331
rect 42628 14300 44005 14328
rect 43993 14297 44005 14300
rect 44039 14297 44051 14331
rect 43993 14291 44051 14297
rect 44085 14331 44143 14337
rect 44085 14297 44097 14331
rect 44131 14328 44143 14331
rect 44174 14328 44180 14340
rect 44131 14300 44180 14328
rect 44131 14297 44143 14300
rect 44085 14291 44143 14297
rect 44174 14288 44180 14300
rect 44232 14288 44238 14340
rect 45646 14288 45652 14340
rect 45704 14328 45710 14340
rect 46658 14328 46664 14340
rect 45704 14300 46664 14328
rect 45704 14288 45710 14300
rect 46658 14288 46664 14300
rect 46716 14288 46722 14340
rect 47026 14288 47032 14340
rect 47084 14288 47090 14340
rect 47210 14288 47216 14340
rect 47268 14288 47274 14340
rect 47394 14288 47400 14340
rect 47452 14328 47458 14340
rect 48685 14331 48743 14337
rect 48685 14328 48697 14331
rect 47452 14300 48697 14328
rect 47452 14288 47458 14300
rect 48685 14297 48697 14300
rect 48731 14297 48743 14331
rect 48685 14291 48743 14297
rect 42610 14260 42616 14272
rect 42260 14232 42616 14260
rect 42610 14220 42616 14232
rect 42668 14260 42674 14272
rect 43898 14260 43904 14272
rect 42668 14232 43904 14260
rect 42668 14220 42674 14232
rect 43898 14220 43904 14232
rect 43956 14220 43962 14272
rect 44192 14260 44220 14288
rect 46014 14260 46020 14272
rect 44192 14232 46020 14260
rect 46014 14220 46020 14232
rect 46072 14220 46078 14272
rect 46290 14220 46296 14272
rect 46348 14260 46354 14272
rect 46385 14263 46443 14269
rect 46385 14260 46397 14263
rect 46348 14232 46397 14260
rect 46348 14220 46354 14232
rect 46385 14229 46397 14232
rect 46431 14229 46443 14263
rect 47228 14260 47256 14288
rect 47581 14263 47639 14269
rect 47581 14260 47593 14263
rect 47228 14232 47593 14260
rect 46385 14223 46443 14229
rect 47581 14229 47593 14232
rect 47627 14260 47639 14263
rect 47765 14263 47823 14269
rect 47765 14260 47777 14263
rect 47627 14232 47777 14260
rect 47627 14229 47639 14232
rect 47581 14223 47639 14229
rect 47765 14229 47777 14232
rect 47811 14260 47823 14263
rect 48590 14260 48596 14272
rect 47811 14232 48596 14260
rect 47811 14229 47823 14232
rect 47765 14223 47823 14229
rect 48590 14220 48596 14232
rect 48648 14220 48654 14272
rect 49053 14263 49111 14269
rect 49053 14229 49065 14263
rect 49099 14260 49111 14263
rect 49142 14260 49148 14272
rect 49099 14232 49148 14260
rect 49099 14229 49111 14232
rect 49053 14223 49111 14229
rect 49142 14220 49148 14232
rect 49200 14220 49206 14272
rect 49344 14260 49372 14359
rect 49528 14328 49556 14368
rect 49602 14356 49608 14408
rect 49660 14356 49666 14408
rect 49970 14356 49976 14408
rect 50028 14356 50034 14408
rect 50062 14356 50068 14408
rect 50120 14396 50126 14408
rect 50249 14399 50307 14405
rect 50249 14396 50261 14399
rect 50120 14368 50261 14396
rect 50120 14356 50126 14368
rect 50249 14365 50261 14368
rect 50295 14365 50307 14399
rect 50249 14359 50307 14365
rect 50522 14356 50528 14408
rect 50580 14356 50586 14408
rect 50614 14356 50620 14408
rect 50672 14356 50678 14408
rect 50430 14328 50436 14340
rect 49528 14300 50436 14328
rect 50430 14288 50436 14300
rect 50488 14288 50494 14340
rect 49694 14260 49700 14272
rect 49344 14232 49700 14260
rect 49694 14220 49700 14232
rect 49752 14220 49758 14272
rect 49786 14220 49792 14272
rect 49844 14260 49850 14272
rect 50632 14260 50660 14356
rect 51718 14288 51724 14340
rect 51776 14288 51782 14340
rect 53742 14328 53748 14340
rect 52946 14300 53748 14328
rect 53742 14288 53748 14300
rect 53800 14288 53806 14340
rect 49844 14232 50660 14260
rect 49844 14220 49850 14232
rect 50798 14220 50804 14272
rect 50856 14220 50862 14272
rect 52546 14220 52552 14272
rect 52604 14260 52610 14272
rect 53193 14263 53251 14269
rect 53193 14260 53205 14263
rect 52604 14232 53205 14260
rect 52604 14220 52610 14232
rect 53193 14229 53205 14232
rect 53239 14229 53251 14263
rect 53193 14223 53251 14229
rect 1104 14170 58880 14192
rect 1104 14118 4874 14170
rect 4926 14118 4938 14170
rect 4990 14118 5002 14170
rect 5054 14118 5066 14170
rect 5118 14118 5130 14170
rect 5182 14118 35594 14170
rect 35646 14118 35658 14170
rect 35710 14118 35722 14170
rect 35774 14118 35786 14170
rect 35838 14118 35850 14170
rect 35902 14118 58880 14170
rect 1104 14096 58880 14118
rect 11698 14016 11704 14068
rect 11756 14056 11762 14068
rect 11756 14028 15240 14056
rect 11756 14016 11762 14028
rect 13170 13948 13176 14000
rect 13228 13948 13234 14000
rect 15212 13988 15240 14028
rect 15286 14016 15292 14068
rect 15344 14016 15350 14068
rect 18046 14016 18052 14068
rect 18104 14056 18110 14068
rect 18325 14059 18383 14065
rect 18325 14056 18337 14059
rect 18104 14028 18337 14056
rect 18104 14016 18110 14028
rect 18325 14025 18337 14028
rect 18371 14025 18383 14059
rect 18325 14019 18383 14025
rect 18969 14059 19027 14065
rect 18969 14025 18981 14059
rect 19015 14056 19027 14059
rect 19426 14056 19432 14068
rect 19015 14028 19432 14056
rect 19015 14025 19027 14028
rect 18969 14019 19027 14025
rect 19426 14016 19432 14028
rect 19484 14056 19490 14068
rect 19484 14028 20300 14056
rect 19484 14016 19490 14028
rect 19337 13991 19395 13997
rect 15212 13960 18644 13988
rect 14306 13906 15424 13920
rect 14292 13892 15424 13906
rect 12158 13812 12164 13864
rect 12216 13852 12222 13864
rect 12897 13855 12955 13861
rect 12897 13852 12909 13855
rect 12216 13824 12909 13852
rect 12216 13812 12222 13824
rect 12897 13821 12909 13824
rect 12943 13821 12955 13855
rect 12897 13815 12955 13821
rect 13630 13812 13636 13864
rect 13688 13852 13694 13864
rect 14292 13852 14320 13892
rect 13688 13824 14320 13852
rect 14645 13855 14703 13861
rect 13688 13812 13694 13824
rect 14645 13821 14657 13855
rect 14691 13852 14703 13855
rect 14734 13852 14740 13864
rect 14691 13824 14740 13852
rect 14691 13821 14703 13824
rect 14645 13815 14703 13821
rect 14734 13812 14740 13824
rect 14792 13812 14798 13864
rect 15396 13852 15424 13892
rect 15470 13880 15476 13932
rect 15528 13920 15534 13932
rect 15841 13923 15899 13929
rect 15841 13920 15853 13923
rect 15528 13892 15853 13920
rect 15528 13880 15534 13892
rect 15841 13889 15853 13892
rect 15887 13889 15899 13923
rect 15841 13883 15899 13889
rect 18138 13880 18144 13932
rect 18196 13880 18202 13932
rect 18616 13929 18644 13960
rect 18708 13960 19288 13988
rect 18417 13923 18475 13929
rect 18417 13889 18429 13923
rect 18463 13889 18475 13923
rect 18417 13883 18475 13889
rect 18601 13923 18659 13929
rect 18601 13889 18613 13923
rect 18647 13889 18659 13923
rect 18601 13883 18659 13889
rect 16758 13852 16764 13864
rect 15396 13824 16764 13852
rect 16758 13812 16764 13824
rect 16816 13812 16822 13864
rect 18432 13852 18460 13883
rect 18708 13852 18736 13960
rect 18785 13923 18843 13929
rect 18785 13889 18797 13923
rect 18831 13889 18843 13923
rect 18785 13883 18843 13889
rect 18432 13824 18736 13852
rect 18800 13852 18828 13883
rect 19150 13880 19156 13932
rect 19208 13880 19214 13932
rect 19260 13920 19288 13960
rect 19337 13957 19349 13991
rect 19383 13988 19395 13991
rect 19383 13960 19656 13988
rect 19383 13957 19395 13960
rect 19337 13951 19395 13957
rect 19628 13929 19656 13960
rect 20272 13932 20300 14028
rect 21836 14028 24164 14056
rect 19613 13923 19671 13929
rect 19260 13892 19564 13920
rect 19334 13852 19340 13864
rect 18800 13824 19340 13852
rect 19334 13812 19340 13824
rect 19392 13812 19398 13864
rect 19536 13725 19564 13892
rect 19613 13889 19625 13923
rect 19659 13889 19671 13923
rect 19613 13883 19671 13889
rect 19628 13852 19656 13883
rect 20254 13880 20260 13932
rect 20312 13880 20318 13932
rect 21450 13880 21456 13932
rect 21508 13920 21514 13932
rect 21836 13929 21864 14028
rect 24136 14000 24164 14028
rect 24578 14016 24584 14068
rect 24636 14016 24642 14068
rect 26970 14056 26976 14068
rect 25148 14028 26976 14056
rect 22094 13948 22100 14000
rect 22152 13948 22158 14000
rect 22186 13948 22192 14000
rect 22244 13988 22250 14000
rect 22244 13960 22586 13988
rect 22244 13948 22250 13960
rect 24118 13948 24124 14000
rect 24176 13988 24182 14000
rect 24596 13988 24624 14016
rect 25148 13988 25176 14028
rect 26970 14016 26976 14028
rect 27028 14016 27034 14068
rect 29914 14016 29920 14068
rect 29972 14056 29978 14068
rect 29972 14028 31156 14056
rect 29972 14016 29978 14028
rect 24176 13960 25176 13988
rect 25317 13991 25375 13997
rect 24176 13948 24182 13960
rect 21821 13923 21879 13929
rect 21821 13920 21833 13923
rect 21508 13892 21833 13920
rect 21508 13880 21514 13892
rect 21821 13889 21833 13892
rect 21867 13889 21879 13923
rect 21821 13883 21879 13889
rect 23842 13880 23848 13932
rect 23900 13880 23906 13932
rect 24210 13880 24216 13932
rect 24268 13880 24274 13932
rect 24302 13880 24308 13932
rect 24360 13880 24366 13932
rect 24394 13880 24400 13932
rect 24452 13920 24458 13932
rect 24581 13923 24639 13929
rect 24452 13892 24497 13920
rect 24452 13880 24458 13892
rect 24581 13889 24593 13923
rect 24627 13889 24639 13923
rect 24581 13883 24639 13889
rect 19889 13855 19947 13861
rect 19889 13852 19901 13855
rect 19628 13824 19901 13852
rect 19889 13821 19901 13824
rect 19935 13852 19947 13855
rect 20073 13855 20131 13861
rect 20073 13852 20085 13855
rect 19935 13824 20085 13852
rect 19935 13821 19947 13824
rect 19889 13815 19947 13821
rect 20073 13821 20085 13824
rect 20119 13852 20131 13855
rect 23860 13852 23888 13880
rect 20119 13824 23888 13852
rect 20119 13821 20131 13824
rect 20073 13815 20131 13821
rect 24486 13812 24492 13864
rect 24544 13852 24550 13864
rect 24596 13852 24624 13883
rect 24670 13880 24676 13932
rect 24728 13880 24734 13932
rect 24854 13929 24860 13932
rect 24811 13923 24860 13929
rect 24811 13889 24823 13923
rect 24857 13889 24860 13923
rect 24811 13883 24860 13889
rect 24854 13880 24860 13883
rect 24912 13880 24918 13932
rect 25056 13929 25084 13960
rect 25317 13957 25329 13991
rect 25363 13988 25375 13991
rect 25590 13988 25596 14000
rect 25363 13960 25596 13988
rect 25363 13957 25375 13960
rect 25317 13951 25375 13957
rect 25590 13948 25596 13960
rect 25648 13948 25654 14000
rect 28350 13988 28356 14000
rect 26542 13960 28356 13988
rect 28350 13948 28356 13960
rect 28408 13948 28414 14000
rect 30374 13988 30380 14000
rect 30130 13960 30380 13988
rect 30374 13948 30380 13960
rect 30432 13948 30438 14000
rect 31018 13988 31024 14000
rect 30484 13960 31024 13988
rect 25041 13923 25099 13929
rect 25041 13889 25053 13923
rect 25087 13889 25099 13923
rect 25041 13883 25099 13889
rect 28626 13880 28632 13932
rect 28684 13880 28690 13932
rect 30484 13920 30512 13960
rect 31018 13948 31024 13960
rect 31076 13948 31082 14000
rect 30392 13892 30512 13920
rect 24544 13824 24624 13852
rect 24544 13812 24550 13824
rect 26786 13812 26792 13864
rect 26844 13812 26850 13864
rect 28902 13812 28908 13864
rect 28960 13812 28966 13864
rect 23382 13744 23388 13796
rect 23440 13784 23446 13796
rect 30392 13793 30420 13892
rect 31018 13812 31024 13864
rect 31076 13812 31082 13864
rect 31128 13852 31156 14028
rect 32858 14016 32864 14068
rect 32916 14056 32922 14068
rect 33045 14059 33103 14065
rect 33045 14056 33057 14059
rect 32916 14028 33057 14056
rect 32916 14016 32922 14028
rect 33045 14025 33057 14028
rect 33091 14025 33103 14059
rect 33045 14019 33103 14025
rect 33413 14059 33471 14065
rect 33413 14025 33425 14059
rect 33459 14056 33471 14059
rect 34330 14056 34336 14068
rect 33459 14028 34336 14056
rect 33459 14025 33471 14028
rect 33413 14019 33471 14025
rect 34330 14016 34336 14028
rect 34388 14056 34394 14068
rect 34425 14059 34483 14065
rect 34425 14056 34437 14059
rect 34388 14028 34437 14056
rect 34388 14016 34394 14028
rect 34425 14025 34437 14028
rect 34471 14025 34483 14059
rect 34425 14019 34483 14025
rect 35713 14059 35771 14065
rect 35713 14025 35725 14059
rect 35759 14056 35771 14059
rect 36170 14056 36176 14068
rect 35759 14028 36176 14056
rect 35759 14025 35771 14028
rect 35713 14019 35771 14025
rect 36170 14016 36176 14028
rect 36228 14016 36234 14068
rect 40678 14056 40684 14068
rect 38672 14028 40684 14056
rect 32766 13948 32772 14000
rect 32824 13948 32830 14000
rect 34238 13988 34244 14000
rect 33336 13960 33824 13988
rect 31662 13880 31668 13932
rect 31720 13920 31726 13932
rect 32125 13923 32183 13929
rect 32125 13920 32137 13923
rect 31720 13892 32137 13920
rect 31720 13880 31726 13892
rect 32125 13889 32137 13892
rect 32171 13889 32183 13923
rect 32125 13883 32183 13889
rect 32582 13880 32588 13932
rect 32640 13880 32646 13932
rect 32953 13923 33011 13929
rect 32953 13889 32965 13923
rect 32999 13920 33011 13923
rect 33336 13920 33364 13960
rect 32999 13892 33364 13920
rect 33428 13892 33732 13920
rect 32999 13889 33011 13892
rect 32953 13883 33011 13889
rect 32217 13855 32275 13861
rect 32217 13852 32229 13855
rect 31128 13824 32229 13852
rect 32217 13821 32229 13824
rect 32263 13852 32275 13855
rect 33428 13852 33456 13892
rect 33704 13864 33732 13892
rect 32263 13824 33456 13852
rect 32263 13821 32275 13824
rect 32217 13815 32275 13821
rect 33502 13812 33508 13864
rect 33560 13812 33566 13864
rect 33686 13812 33692 13864
rect 33744 13812 33750 13864
rect 33796 13852 33824 13960
rect 33888 13960 34244 13988
rect 33888 13929 33916 13960
rect 34238 13948 34244 13960
rect 34296 13948 34302 14000
rect 35986 13948 35992 14000
rect 36044 13948 36050 14000
rect 36081 13991 36139 13997
rect 36081 13957 36093 13991
rect 36127 13988 36139 13991
rect 38562 13988 38568 14000
rect 36127 13960 38568 13988
rect 36127 13957 36139 13960
rect 36081 13951 36139 13957
rect 38562 13948 38568 13960
rect 38620 13948 38626 14000
rect 33873 13923 33931 13929
rect 33873 13889 33885 13923
rect 33919 13889 33931 13923
rect 34514 13920 34520 13932
rect 33873 13883 33931 13889
rect 33980 13892 34520 13920
rect 33980 13852 34008 13892
rect 34514 13880 34520 13892
rect 34572 13880 34578 13932
rect 35250 13880 35256 13932
rect 35308 13920 35314 13932
rect 35897 13923 35955 13929
rect 35897 13920 35909 13923
rect 35308 13892 35909 13920
rect 35308 13880 35314 13892
rect 35897 13889 35909 13892
rect 35943 13889 35955 13923
rect 35897 13883 35955 13889
rect 36262 13880 36268 13932
rect 36320 13880 36326 13932
rect 36538 13880 36544 13932
rect 36596 13920 36602 13932
rect 36633 13923 36691 13929
rect 36633 13920 36645 13923
rect 36596 13892 36645 13920
rect 36596 13880 36602 13892
rect 36633 13889 36645 13892
rect 36679 13889 36691 13923
rect 36633 13883 36691 13889
rect 36725 13923 36783 13929
rect 36725 13889 36737 13923
rect 36771 13889 36783 13923
rect 36725 13883 36783 13889
rect 36909 13923 36967 13929
rect 36909 13889 36921 13923
rect 36955 13889 36967 13923
rect 36909 13883 36967 13889
rect 33796 13824 34008 13852
rect 36354 13812 36360 13864
rect 36412 13852 36418 13864
rect 36740 13852 36768 13883
rect 36412 13824 36768 13852
rect 36924 13852 36952 13883
rect 36998 13880 37004 13932
rect 37056 13880 37062 13932
rect 37274 13880 37280 13932
rect 37332 13920 37338 13932
rect 38672 13929 38700 14028
rect 40678 14016 40684 14028
rect 40736 14056 40742 14068
rect 41322 14056 41328 14068
rect 40736 14028 41328 14056
rect 40736 14016 40742 14028
rect 41322 14016 41328 14028
rect 41380 14056 41386 14068
rect 41380 14028 42288 14056
rect 41380 14016 41386 14028
rect 40494 13988 40500 14000
rect 40158 13960 40500 13988
rect 40494 13948 40500 13960
rect 40552 13948 40558 14000
rect 41506 13948 41512 14000
rect 41564 13948 41570 14000
rect 41969 13991 42027 13997
rect 41969 13957 41981 13991
rect 42015 13988 42027 13991
rect 42058 13988 42064 14000
rect 42015 13960 42064 13988
rect 42015 13957 42027 13960
rect 41969 13951 42027 13957
rect 42058 13948 42064 13960
rect 42116 13948 42122 14000
rect 42260 13929 42288 14028
rect 44082 14016 44088 14068
rect 44140 14056 44146 14068
rect 44177 14059 44235 14065
rect 44177 14056 44189 14059
rect 44140 14028 44189 14056
rect 44140 14016 44146 14028
rect 44177 14025 44189 14028
rect 44223 14025 44235 14059
rect 44177 14019 44235 14025
rect 44266 14016 44272 14068
rect 44324 14016 44330 14068
rect 46014 14016 46020 14068
rect 46072 14056 46078 14068
rect 46109 14059 46167 14065
rect 46109 14056 46121 14059
rect 46072 14028 46121 14056
rect 46072 14016 46078 14028
rect 46109 14025 46121 14028
rect 46155 14025 46167 14059
rect 46109 14019 46167 14025
rect 46293 14059 46351 14065
rect 46293 14025 46305 14059
rect 46339 14056 46351 14059
rect 46566 14056 46572 14068
rect 46339 14028 46572 14056
rect 46339 14025 46351 14028
rect 46293 14019 46351 14025
rect 46566 14016 46572 14028
rect 46624 14016 46630 14068
rect 47121 14059 47179 14065
rect 47121 14056 47133 14059
rect 46676 14028 47133 14056
rect 46676 14000 46704 14028
rect 47121 14025 47133 14028
rect 47167 14025 47179 14059
rect 47121 14019 47179 14025
rect 47578 14016 47584 14068
rect 47636 14016 47642 14068
rect 51074 14056 51080 14068
rect 48424 14028 51080 14056
rect 42702 13948 42708 14000
rect 42760 13948 42766 14000
rect 43438 13948 43444 14000
rect 43496 13948 43502 14000
rect 46198 13948 46204 14000
rect 46256 13988 46262 14000
rect 46256 13960 46612 13988
rect 46256 13948 46262 13960
rect 46584 13932 46612 13960
rect 46658 13948 46664 14000
rect 46716 13948 46722 14000
rect 47394 13988 47400 14000
rect 46860 13960 47400 13988
rect 38657 13923 38715 13929
rect 38657 13920 38669 13923
rect 37332 13892 38669 13920
rect 37332 13880 37338 13892
rect 38657 13889 38669 13892
rect 38703 13889 38715 13923
rect 38657 13883 38715 13889
rect 42245 13923 42303 13929
rect 42245 13889 42257 13923
rect 42291 13920 42303 13923
rect 42429 13923 42487 13929
rect 42429 13920 42441 13923
rect 42291 13892 42441 13920
rect 42291 13889 42303 13892
rect 42245 13883 42303 13889
rect 42429 13889 42441 13892
rect 42475 13889 42487 13923
rect 42429 13883 42487 13889
rect 43990 13880 43996 13932
rect 44048 13920 44054 13932
rect 44450 13920 44456 13932
rect 44048 13892 44456 13920
rect 44048 13880 44054 13892
rect 44450 13880 44456 13892
rect 44508 13880 44514 13932
rect 44542 13880 44548 13932
rect 44600 13880 44606 13932
rect 44634 13880 44640 13932
rect 44692 13920 44698 13932
rect 44821 13923 44879 13929
rect 44821 13920 44833 13923
rect 44692 13892 44833 13920
rect 44692 13880 44698 13892
rect 44821 13889 44833 13892
rect 44867 13889 44879 13923
rect 44821 13883 44879 13889
rect 45646 13880 45652 13932
rect 45704 13920 45710 13932
rect 46474 13929 46480 13932
rect 45925 13923 45983 13929
rect 45925 13920 45937 13923
rect 45704 13892 45937 13920
rect 45704 13880 45710 13892
rect 45925 13889 45937 13892
rect 45971 13889 45983 13923
rect 46472 13920 46480 13929
rect 46435 13892 46480 13920
rect 45925 13883 45983 13889
rect 46472 13883 46480 13892
rect 46474 13880 46480 13883
rect 46532 13880 46538 13932
rect 46566 13880 46572 13932
rect 46624 13880 46630 13932
rect 46860 13929 46888 13960
rect 47394 13948 47400 13960
rect 47452 13948 47458 14000
rect 46844 13923 46902 13929
rect 46844 13889 46856 13923
rect 46890 13889 46902 13923
rect 46844 13883 46902 13889
rect 46937 13923 46995 13929
rect 46937 13889 46949 13923
rect 46983 13889 46995 13923
rect 46937 13883 46995 13889
rect 37734 13852 37740 13864
rect 36924 13824 37740 13852
rect 36412 13812 36418 13824
rect 37734 13812 37740 13824
rect 37792 13812 37798 13864
rect 38930 13812 38936 13864
rect 38988 13812 38994 13864
rect 40402 13812 40408 13864
rect 40460 13812 40466 13864
rect 40497 13855 40555 13861
rect 40497 13821 40509 13855
rect 40543 13852 40555 13855
rect 40586 13852 40592 13864
rect 40543 13824 40592 13852
rect 40543 13821 40555 13824
rect 40497 13815 40555 13821
rect 40586 13812 40592 13824
rect 40644 13852 40650 13864
rect 42334 13852 42340 13864
rect 40644 13824 42340 13852
rect 40644 13812 40650 13824
rect 42334 13812 42340 13824
rect 42392 13812 42398 13864
rect 43070 13812 43076 13864
rect 43128 13852 43134 13864
rect 44729 13855 44787 13861
rect 44729 13852 44741 13855
rect 43128 13824 44741 13852
rect 43128 13812 43134 13824
rect 44729 13821 44741 13824
rect 44775 13852 44787 13855
rect 46750 13852 46756 13864
rect 44775 13824 46756 13852
rect 44775 13821 44787 13824
rect 44729 13815 44787 13821
rect 46750 13812 46756 13824
rect 46808 13812 46814 13864
rect 46952 13852 46980 13883
rect 47118 13880 47124 13932
rect 47176 13920 47182 13932
rect 47305 13923 47363 13929
rect 47305 13920 47317 13923
rect 47176 13892 47317 13920
rect 47176 13880 47182 13892
rect 47305 13889 47317 13892
rect 47351 13889 47363 13923
rect 47305 13883 47363 13889
rect 48225 13923 48283 13929
rect 48225 13889 48237 13923
rect 48271 13920 48283 13923
rect 48314 13920 48320 13932
rect 48271 13892 48320 13920
rect 48271 13889 48283 13892
rect 48225 13883 48283 13889
rect 47210 13852 47216 13864
rect 46952 13824 47216 13852
rect 47210 13812 47216 13824
rect 47268 13812 47274 13864
rect 47320 13852 47348 13883
rect 48314 13880 48320 13892
rect 48372 13880 48378 13932
rect 48424 13861 48452 14028
rect 51074 14016 51080 14028
rect 51132 14016 51138 14068
rect 51166 14016 51172 14068
rect 51224 14056 51230 14068
rect 51994 14056 52000 14068
rect 51224 14028 52000 14056
rect 51224 14016 51230 14028
rect 51994 14016 52000 14028
rect 52052 14056 52058 14068
rect 53101 14059 53159 14065
rect 53101 14056 53113 14059
rect 52052 14028 52224 14056
rect 52052 14016 52058 14028
rect 50709 13991 50767 13997
rect 50709 13988 50721 13991
rect 49436 13960 50721 13988
rect 48774 13880 48780 13932
rect 48832 13920 48838 13932
rect 49050 13920 49056 13932
rect 48832 13892 49056 13920
rect 48832 13880 48838 13892
rect 49050 13880 49056 13892
rect 49108 13880 49114 13932
rect 49142 13880 49148 13932
rect 49200 13880 49206 13932
rect 49436 13929 49464 13960
rect 50709 13957 50721 13960
rect 50755 13957 50767 13991
rect 50709 13951 50767 13957
rect 50798 13948 50804 14000
rect 50856 13988 50862 14000
rect 52196 13997 52224 14028
rect 52288 14028 53113 14056
rect 52181 13991 52239 13997
rect 50856 13960 51764 13988
rect 50856 13948 50862 13960
rect 49421 13923 49479 13929
rect 49421 13889 49433 13923
rect 49467 13889 49479 13923
rect 49421 13883 49479 13889
rect 49786 13880 49792 13932
rect 49844 13880 49850 13932
rect 50522 13880 50528 13932
rect 50580 13920 50586 13932
rect 51261 13923 51319 13929
rect 51261 13920 51273 13923
rect 50580 13892 51273 13920
rect 50580 13880 50586 13892
rect 51261 13889 51273 13892
rect 51307 13889 51319 13923
rect 51261 13883 51319 13889
rect 51626 13880 51632 13932
rect 51684 13880 51690 13932
rect 51736 13929 51764 13960
rect 52181 13957 52193 13991
rect 52227 13957 52239 13991
rect 52181 13951 52239 13957
rect 51721 13923 51779 13929
rect 51721 13889 51733 13923
rect 51767 13889 51779 13923
rect 51721 13883 51779 13889
rect 51902 13880 51908 13932
rect 51960 13920 51966 13932
rect 51997 13923 52055 13929
rect 51997 13920 52009 13923
rect 51960 13892 52009 13920
rect 51960 13880 51966 13892
rect 51997 13889 52009 13892
rect 52043 13889 52055 13923
rect 51997 13883 52055 13889
rect 48409 13855 48467 13861
rect 48409 13852 48421 13855
rect 47320 13824 48421 13852
rect 48409 13821 48421 13824
rect 48455 13821 48467 13855
rect 48409 13815 48467 13821
rect 48590 13812 48596 13864
rect 48648 13852 48654 13864
rect 50982 13852 50988 13864
rect 48648 13824 50988 13852
rect 48648 13812 48654 13824
rect 50982 13812 50988 13824
rect 51040 13812 51046 13864
rect 51810 13812 51816 13864
rect 51868 13852 51874 13864
rect 52288 13852 52316 14028
rect 53101 14025 53113 14028
rect 53147 14056 53159 14059
rect 53742 14056 53748 14068
rect 53147 14028 53748 14056
rect 53147 14025 53159 14028
rect 53101 14019 53159 14025
rect 53742 14016 53748 14028
rect 53800 14016 53806 14068
rect 52362 13948 52368 14000
rect 52420 13988 52426 14000
rect 52825 13991 52883 13997
rect 52825 13988 52837 13991
rect 52420 13960 52837 13988
rect 52420 13948 52426 13960
rect 52825 13957 52837 13960
rect 52871 13988 52883 13991
rect 53285 13991 53343 13997
rect 53285 13988 53297 13991
rect 52871 13960 53297 13988
rect 52871 13957 52883 13960
rect 52825 13951 52883 13957
rect 53285 13957 53297 13960
rect 53331 13957 53343 13991
rect 53285 13951 53343 13957
rect 57606 13880 57612 13932
rect 57664 13920 57670 13932
rect 58253 13923 58311 13929
rect 58253 13920 58265 13923
rect 57664 13892 58265 13920
rect 57664 13880 57670 13892
rect 58253 13889 58265 13892
rect 58299 13889 58311 13923
rect 58253 13883 58311 13889
rect 51868 13824 52316 13852
rect 51868 13812 51874 13824
rect 23569 13787 23627 13793
rect 23569 13784 23581 13787
rect 23440 13756 23581 13784
rect 23440 13744 23446 13756
rect 23569 13753 23581 13756
rect 23615 13753 23627 13787
rect 23569 13747 23627 13753
rect 30377 13787 30435 13793
rect 30377 13753 30389 13787
rect 30423 13753 30435 13787
rect 30377 13747 30435 13753
rect 32766 13744 32772 13796
rect 32824 13784 32830 13796
rect 34057 13787 34115 13793
rect 34057 13784 34069 13787
rect 32824 13756 34069 13784
rect 32824 13744 32830 13756
rect 34057 13753 34069 13756
rect 34103 13784 34115 13787
rect 34609 13787 34667 13793
rect 34609 13784 34621 13787
rect 34103 13756 34621 13784
rect 34103 13753 34115 13756
rect 34057 13747 34115 13753
rect 34609 13753 34621 13756
rect 34655 13753 34667 13787
rect 34609 13747 34667 13753
rect 36078 13744 36084 13796
rect 36136 13784 36142 13796
rect 36538 13784 36544 13796
rect 36136 13756 36544 13784
rect 36136 13744 36142 13756
rect 36538 13744 36544 13756
rect 36596 13784 36602 13796
rect 37090 13784 37096 13796
rect 36596 13756 37096 13784
rect 36596 13744 36602 13756
rect 37090 13744 37096 13756
rect 37148 13784 37154 13796
rect 37642 13784 37648 13796
rect 37148 13756 37648 13784
rect 37148 13744 37154 13756
rect 37642 13744 37648 13756
rect 37700 13744 37706 13796
rect 51718 13784 51724 13796
rect 39960 13756 40632 13784
rect 19521 13719 19579 13725
rect 19521 13685 19533 13719
rect 19567 13716 19579 13719
rect 19978 13716 19984 13728
rect 19567 13688 19984 13716
rect 19567 13685 19579 13688
rect 19521 13679 19579 13685
rect 19978 13676 19984 13688
rect 20036 13676 20042 13728
rect 24949 13719 25007 13725
rect 24949 13685 24961 13719
rect 24995 13716 25007 13719
rect 25774 13716 25780 13728
rect 24995 13688 25780 13716
rect 24995 13685 25007 13688
rect 24949 13679 25007 13685
rect 25774 13676 25780 13688
rect 25832 13676 25838 13728
rect 30466 13676 30472 13728
rect 30524 13676 30530 13728
rect 36446 13676 36452 13728
rect 36504 13676 36510 13728
rect 36814 13676 36820 13728
rect 36872 13716 36878 13728
rect 39960 13716 39988 13756
rect 36872 13688 39988 13716
rect 40604 13716 40632 13756
rect 44100 13756 51724 13784
rect 44100 13716 44128 13756
rect 51718 13744 51724 13756
rect 51776 13744 51782 13796
rect 40604 13688 44128 13716
rect 36872 13676 36878 13688
rect 48682 13676 48688 13728
rect 48740 13676 48746 13728
rect 48869 13719 48927 13725
rect 48869 13685 48881 13719
rect 48915 13716 48927 13719
rect 49050 13716 49056 13728
rect 48915 13688 49056 13716
rect 48915 13685 48927 13688
rect 48869 13679 48927 13685
rect 49050 13676 49056 13688
rect 49108 13676 49114 13728
rect 49234 13676 49240 13728
rect 49292 13716 49298 13728
rect 49329 13719 49387 13725
rect 49329 13716 49341 13719
rect 49292 13688 49341 13716
rect 49292 13676 49298 13688
rect 49329 13685 49341 13688
rect 49375 13685 49387 13719
rect 49329 13679 49387 13685
rect 51442 13676 51448 13728
rect 51500 13676 51506 13728
rect 51920 13725 51948 13824
rect 51905 13719 51963 13725
rect 51905 13685 51917 13719
rect 51951 13685 51963 13719
rect 51905 13679 51963 13685
rect 52270 13676 52276 13728
rect 52328 13716 52334 13728
rect 52730 13716 52736 13728
rect 52328 13688 52736 13716
rect 52328 13676 52334 13688
rect 52730 13676 52736 13688
rect 52788 13716 52794 13728
rect 53469 13719 53527 13725
rect 53469 13716 53481 13719
rect 52788 13688 53481 13716
rect 52788 13676 52794 13688
rect 53469 13685 53481 13688
rect 53515 13685 53527 13719
rect 53469 13679 53527 13685
rect 58434 13676 58440 13728
rect 58492 13676 58498 13728
rect 1104 13626 58880 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 58880 13626
rect 1104 13552 58880 13574
rect 13446 13472 13452 13524
rect 13504 13512 13510 13524
rect 13725 13515 13783 13521
rect 13725 13512 13737 13515
rect 13504 13484 13737 13512
rect 13504 13472 13510 13484
rect 13725 13481 13737 13484
rect 13771 13481 13783 13515
rect 13725 13475 13783 13481
rect 12250 13336 12256 13388
rect 12308 13336 12314 13388
rect 11977 13311 12035 13317
rect 11977 13277 11989 13311
rect 12023 13277 12035 13311
rect 11977 13271 12035 13277
rect 11992 13240 12020 13271
rect 12158 13240 12164 13252
rect 11992 13212 12164 13240
rect 12158 13200 12164 13212
rect 12216 13200 12222 13252
rect 13630 13240 13636 13252
rect 13478 13212 13636 13240
rect 13630 13200 13636 13212
rect 13688 13200 13694 13252
rect 13740 13240 13768 13475
rect 15194 13472 15200 13524
rect 15252 13512 15258 13524
rect 15289 13515 15347 13521
rect 15289 13512 15301 13515
rect 15252 13484 15301 13512
rect 15252 13472 15258 13484
rect 15289 13481 15301 13484
rect 15335 13481 15347 13515
rect 15289 13475 15347 13481
rect 24029 13515 24087 13521
rect 24029 13481 24041 13515
rect 24075 13512 24087 13515
rect 24302 13512 24308 13524
rect 24075 13484 24308 13512
rect 24075 13481 24087 13484
rect 24029 13475 24087 13481
rect 24302 13472 24308 13484
rect 24360 13512 24366 13524
rect 24673 13515 24731 13521
rect 24673 13512 24685 13515
rect 24360 13484 24685 13512
rect 24360 13472 24366 13484
rect 24673 13481 24685 13484
rect 24719 13481 24731 13515
rect 24673 13475 24731 13481
rect 28902 13472 28908 13524
rect 28960 13512 28966 13524
rect 29549 13515 29607 13521
rect 29549 13512 29561 13515
rect 28960 13484 29561 13512
rect 28960 13472 28966 13484
rect 29549 13481 29561 13484
rect 29595 13481 29607 13515
rect 29549 13475 29607 13481
rect 32766 13472 32772 13524
rect 32824 13512 32830 13524
rect 33045 13515 33103 13521
rect 33045 13512 33057 13515
rect 32824 13484 33057 13512
rect 32824 13472 32830 13484
rect 33045 13481 33057 13484
rect 33091 13481 33103 13515
rect 33045 13475 33103 13481
rect 35434 13472 35440 13524
rect 35492 13512 35498 13524
rect 35989 13515 36047 13521
rect 35989 13512 36001 13515
rect 35492 13484 36001 13512
rect 35492 13472 35498 13484
rect 35989 13481 36001 13484
rect 36035 13481 36047 13515
rect 35989 13475 36047 13481
rect 36262 13472 36268 13524
rect 36320 13472 36326 13524
rect 36446 13472 36452 13524
rect 36504 13472 36510 13524
rect 36538 13472 36544 13524
rect 36596 13512 36602 13524
rect 36596 13484 37504 13512
rect 36596 13472 36602 13484
rect 27982 13404 27988 13456
rect 28040 13444 28046 13456
rect 29730 13444 29736 13456
rect 28040 13416 29736 13444
rect 28040 13404 28046 13416
rect 29730 13404 29736 13416
rect 29788 13404 29794 13456
rect 29822 13404 29828 13456
rect 29880 13444 29886 13456
rect 37182 13444 37188 13456
rect 29880 13416 32444 13444
rect 29880 13404 29886 13416
rect 14734 13336 14740 13388
rect 14792 13376 14798 13388
rect 14792 13348 15056 13376
rect 14792 13336 14798 13348
rect 14918 13268 14924 13320
rect 14976 13268 14982 13320
rect 15028 13317 15056 13348
rect 15654 13336 15660 13388
rect 15712 13376 15718 13388
rect 16393 13379 16451 13385
rect 16393 13376 16405 13379
rect 15712 13348 16405 13376
rect 15712 13336 15718 13348
rect 16393 13345 16405 13348
rect 16439 13345 16451 13379
rect 16393 13339 16451 13345
rect 16666 13336 16672 13388
rect 16724 13336 16730 13388
rect 17310 13336 17316 13388
rect 17368 13336 17374 13388
rect 17954 13336 17960 13388
rect 18012 13376 18018 13388
rect 20073 13379 20131 13385
rect 20073 13376 20085 13379
rect 18012 13348 20085 13376
rect 18012 13336 18018 13348
rect 15013 13311 15071 13317
rect 15013 13277 15025 13311
rect 15059 13277 15071 13311
rect 15013 13271 15071 13277
rect 15381 13311 15439 13317
rect 15381 13277 15393 13311
rect 15427 13308 15439 13311
rect 16574 13308 16580 13320
rect 15427 13280 16580 13308
rect 15427 13277 15439 13280
rect 15381 13271 15439 13277
rect 16574 13268 16580 13280
rect 16632 13268 16638 13320
rect 16761 13311 16819 13317
rect 16761 13277 16773 13311
rect 16807 13308 16819 13311
rect 16850 13308 16856 13320
rect 16807 13280 16856 13308
rect 16807 13277 16819 13280
rect 16761 13271 16819 13277
rect 16850 13268 16856 13280
rect 16908 13268 16914 13320
rect 17034 13268 17040 13320
rect 17092 13268 17098 13320
rect 17218 13268 17224 13320
rect 17276 13268 17282 13320
rect 18708 13294 18736 13348
rect 20073 13345 20085 13348
rect 20119 13345 20131 13379
rect 20073 13339 20131 13345
rect 23661 13379 23719 13385
rect 23661 13345 23673 13379
rect 23707 13376 23719 13379
rect 23842 13376 23848 13388
rect 23707 13348 23848 13376
rect 23707 13345 23719 13348
rect 23661 13339 23719 13345
rect 23842 13336 23848 13348
rect 23900 13376 23906 13388
rect 26418 13376 26424 13388
rect 23900 13348 26424 13376
rect 23900 13336 23906 13348
rect 26418 13336 26424 13348
rect 26476 13336 26482 13388
rect 26605 13379 26663 13385
rect 26605 13345 26617 13379
rect 26651 13376 26663 13379
rect 27154 13376 27160 13388
rect 26651 13348 27160 13376
rect 26651 13345 26663 13348
rect 26605 13339 26663 13345
rect 27154 13336 27160 13348
rect 27212 13376 27218 13388
rect 29086 13376 29092 13388
rect 27212 13348 29092 13376
rect 27212 13336 27218 13348
rect 29086 13336 29092 13348
rect 29144 13336 29150 13388
rect 30006 13336 30012 13388
rect 30064 13336 30070 13388
rect 19797 13311 19855 13317
rect 19797 13308 19809 13311
rect 19076 13280 19809 13308
rect 14737 13243 14795 13249
rect 14737 13240 14749 13243
rect 13740 13212 14749 13240
rect 14737 13209 14749 13212
rect 14783 13209 14795 13243
rect 14737 13203 14795 13209
rect 16209 13243 16267 13249
rect 16209 13209 16221 13243
rect 16255 13240 16267 13243
rect 17310 13240 17316 13252
rect 16255 13212 17316 13240
rect 16255 13209 16267 13212
rect 16209 13203 16267 13209
rect 17310 13200 17316 13212
rect 17368 13200 17374 13252
rect 17589 13243 17647 13249
rect 17589 13209 17601 13243
rect 17635 13209 17647 13243
rect 17589 13203 17647 13209
rect 15102 13132 15108 13184
rect 15160 13172 15166 13184
rect 17034 13172 17040 13184
rect 15160 13144 17040 13172
rect 15160 13132 15166 13144
rect 17034 13132 17040 13144
rect 17092 13132 17098 13184
rect 17129 13175 17187 13181
rect 17129 13141 17141 13175
rect 17175 13172 17187 13175
rect 17604 13172 17632 13203
rect 17175 13144 17632 13172
rect 17175 13141 17187 13144
rect 17129 13135 17187 13141
rect 17954 13132 17960 13184
rect 18012 13172 18018 13184
rect 19076 13181 19104 13280
rect 19797 13277 19809 13280
rect 19843 13277 19855 13311
rect 19797 13271 19855 13277
rect 20349 13311 20407 13317
rect 20349 13277 20361 13311
rect 20395 13308 20407 13311
rect 20622 13308 20628 13320
rect 20395 13280 20628 13308
rect 20395 13277 20407 13280
rect 20349 13271 20407 13277
rect 20622 13268 20628 13280
rect 20680 13268 20686 13320
rect 23934 13268 23940 13320
rect 23992 13308 23998 13320
rect 24121 13311 24179 13317
rect 24121 13308 24133 13311
rect 23992 13280 24133 13308
rect 23992 13268 23998 13280
rect 24121 13277 24133 13280
rect 24167 13277 24179 13311
rect 24121 13271 24179 13277
rect 24136 13240 24164 13271
rect 24394 13268 24400 13320
rect 24452 13308 24458 13320
rect 24857 13311 24915 13317
rect 24857 13308 24869 13311
rect 24452 13280 24869 13308
rect 24452 13268 24458 13280
rect 24857 13277 24869 13280
rect 24903 13277 24915 13311
rect 24857 13271 24915 13277
rect 26881 13311 26939 13317
rect 26881 13277 26893 13311
rect 26927 13308 26939 13311
rect 27982 13308 27988 13320
rect 26927 13280 27988 13308
rect 26927 13277 26939 13280
rect 26881 13271 26939 13277
rect 27982 13268 27988 13280
rect 28040 13268 28046 13320
rect 29730 13268 29736 13320
rect 29788 13268 29794 13320
rect 29825 13311 29883 13317
rect 29825 13277 29837 13311
rect 29871 13277 29883 13311
rect 29825 13271 29883 13277
rect 30101 13311 30159 13317
rect 30101 13277 30113 13311
rect 30147 13308 30159 13311
rect 30466 13308 30472 13320
rect 30147 13280 30472 13308
rect 30147 13277 30159 13280
rect 30101 13271 30159 13277
rect 24489 13243 24547 13249
rect 24489 13240 24501 13243
rect 24136 13212 24501 13240
rect 24489 13209 24501 13212
rect 24535 13240 24547 13243
rect 29638 13240 29644 13252
rect 24535 13212 29644 13240
rect 24535 13209 24547 13212
rect 24489 13203 24547 13209
rect 29638 13200 29644 13212
rect 29696 13200 29702 13252
rect 29840 13240 29868 13271
rect 30466 13268 30472 13280
rect 30524 13268 30530 13320
rect 30837 13311 30895 13317
rect 30837 13277 30849 13311
rect 30883 13308 30895 13311
rect 30926 13308 30932 13320
rect 30883 13280 30932 13308
rect 30883 13277 30895 13280
rect 30837 13271 30895 13277
rect 30926 13268 30932 13280
rect 30984 13268 30990 13320
rect 31110 13268 31116 13320
rect 31168 13268 31174 13320
rect 32125 13311 32183 13317
rect 32125 13277 32137 13311
rect 32171 13277 32183 13311
rect 32125 13271 32183 13277
rect 30653 13243 30711 13249
rect 30653 13240 30665 13243
rect 29840 13212 30665 13240
rect 30653 13209 30665 13212
rect 30699 13209 30711 13243
rect 32140 13240 32168 13271
rect 32306 13268 32312 13320
rect 32364 13268 32370 13320
rect 32416 13317 32444 13416
rect 35912 13416 37188 13444
rect 35912 13385 35940 13416
rect 37182 13404 37188 13416
rect 37240 13444 37246 13456
rect 37476 13444 37504 13484
rect 37642 13472 37648 13524
rect 37700 13472 37706 13524
rect 37734 13472 37740 13524
rect 37792 13472 37798 13524
rect 38930 13472 38936 13524
rect 38988 13512 38994 13524
rect 39025 13515 39083 13521
rect 39025 13512 39037 13515
rect 38988 13484 39037 13512
rect 38988 13472 38994 13484
rect 39025 13481 39037 13484
rect 39071 13481 39083 13515
rect 39025 13475 39083 13481
rect 41046 13472 41052 13524
rect 41104 13472 41110 13524
rect 41506 13472 41512 13524
rect 41564 13512 41570 13524
rect 42153 13515 42211 13521
rect 42153 13512 42165 13515
rect 41564 13484 42165 13512
rect 41564 13472 41570 13484
rect 42153 13481 42165 13484
rect 42199 13512 42211 13515
rect 42426 13512 42432 13524
rect 42199 13484 42432 13512
rect 42199 13481 42211 13484
rect 42153 13475 42211 13481
rect 42426 13472 42432 13484
rect 42484 13472 42490 13524
rect 45370 13472 45376 13524
rect 45428 13512 45434 13524
rect 45833 13515 45891 13521
rect 45833 13512 45845 13515
rect 45428 13484 45845 13512
rect 45428 13472 45434 13484
rect 45833 13481 45845 13484
rect 45879 13481 45891 13515
rect 45833 13475 45891 13481
rect 48498 13472 48504 13524
rect 48556 13472 48562 13524
rect 48774 13472 48780 13524
rect 48832 13472 48838 13524
rect 51902 13472 51908 13524
rect 51960 13472 51966 13524
rect 51994 13472 52000 13524
rect 52052 13472 52058 13524
rect 54849 13515 54907 13521
rect 54849 13481 54861 13515
rect 54895 13512 54907 13515
rect 54938 13512 54944 13524
rect 54895 13484 54944 13512
rect 54895 13481 54907 13484
rect 54849 13475 54907 13481
rect 54938 13472 54944 13484
rect 54996 13472 55002 13524
rect 37826 13444 37832 13456
rect 37240 13416 37320 13444
rect 37476 13416 37832 13444
rect 37240 13404 37246 13416
rect 35897 13379 35955 13385
rect 35897 13345 35909 13379
rect 35943 13345 35955 13379
rect 36630 13376 36636 13388
rect 35897 13339 35955 13345
rect 36188 13348 36636 13376
rect 32401 13311 32459 13317
rect 32401 13277 32413 13311
rect 32447 13308 32459 13311
rect 33318 13308 33324 13320
rect 32447 13280 33324 13308
rect 32447 13277 32459 13280
rect 32401 13271 32459 13277
rect 33318 13268 33324 13280
rect 33376 13308 33382 13320
rect 36078 13308 36084 13320
rect 33376 13280 36084 13308
rect 33376 13268 33382 13280
rect 36078 13268 36084 13280
rect 36136 13268 36142 13320
rect 36188 13317 36216 13348
rect 36630 13336 36636 13348
rect 36688 13376 36694 13388
rect 37001 13379 37059 13385
rect 37001 13376 37013 13379
rect 36688 13348 37013 13376
rect 36688 13336 36694 13348
rect 37001 13345 37013 13348
rect 37047 13345 37059 13379
rect 37001 13339 37059 13345
rect 36173 13311 36231 13317
rect 36173 13277 36185 13311
rect 36219 13277 36231 13311
rect 36173 13271 36231 13277
rect 36446 13268 36452 13320
rect 36504 13268 36510 13320
rect 36538 13268 36544 13320
rect 36596 13268 36602 13320
rect 32582 13240 32588 13252
rect 32140 13212 32588 13240
rect 30653 13203 30711 13209
rect 32582 13200 32588 13212
rect 32640 13240 32646 13252
rect 33962 13240 33968 13252
rect 32640 13212 33968 13240
rect 32640 13200 32646 13212
rect 33962 13200 33968 13212
rect 34020 13200 34026 13252
rect 36906 13200 36912 13252
rect 36964 13200 36970 13252
rect 37016 13240 37044 13339
rect 37090 13336 37096 13388
rect 37148 13336 37154 13388
rect 37292 13317 37320 13416
rect 37826 13404 37832 13416
rect 37884 13444 37890 13456
rect 37921 13447 37979 13453
rect 37921 13444 37933 13447
rect 37884 13416 37933 13444
rect 37884 13404 37890 13416
rect 37921 13413 37933 13416
rect 37967 13413 37979 13447
rect 37921 13407 37979 13413
rect 38470 13404 38476 13456
rect 38528 13444 38534 13456
rect 40034 13444 40040 13456
rect 38528 13416 40040 13444
rect 38528 13404 38534 13416
rect 40034 13404 40040 13416
rect 40092 13404 40098 13456
rect 51718 13404 51724 13456
rect 51776 13444 51782 13456
rect 54573 13447 54631 13453
rect 54573 13444 54585 13447
rect 51776 13416 54585 13444
rect 51776 13404 51782 13416
rect 54573 13413 54585 13416
rect 54619 13444 54631 13447
rect 55309 13447 55367 13453
rect 55309 13444 55321 13447
rect 54619 13416 55321 13444
rect 54619 13413 54631 13416
rect 54573 13407 54631 13413
rect 55309 13413 55321 13416
rect 55355 13444 55367 13447
rect 55355 13416 55628 13444
rect 55355 13413 55367 13416
rect 55309 13407 55367 13413
rect 37553 13379 37611 13385
rect 37553 13376 37565 13379
rect 37384 13348 37565 13376
rect 37277 13311 37335 13317
rect 37277 13277 37289 13311
rect 37323 13277 37335 13311
rect 37277 13271 37335 13277
rect 37384 13240 37412 13348
rect 37553 13345 37565 13348
rect 37599 13345 37611 13379
rect 37553 13339 37611 13345
rect 39669 13379 39727 13385
rect 39669 13345 39681 13379
rect 39715 13376 39727 13379
rect 40126 13376 40132 13388
rect 39715 13348 40132 13376
rect 39715 13345 39727 13348
rect 39669 13339 39727 13345
rect 40126 13336 40132 13348
rect 40184 13336 40190 13388
rect 40678 13336 40684 13388
rect 40736 13376 40742 13388
rect 40773 13379 40831 13385
rect 40773 13376 40785 13379
rect 40736 13348 40785 13376
rect 40736 13336 40742 13348
rect 40773 13345 40785 13348
rect 40819 13345 40831 13379
rect 40773 13339 40831 13345
rect 44910 13336 44916 13388
rect 44968 13376 44974 13388
rect 46017 13379 46075 13385
rect 46017 13376 46029 13379
rect 44968 13348 46029 13376
rect 44968 13336 44974 13348
rect 46017 13345 46029 13348
rect 46063 13345 46075 13379
rect 46017 13339 46075 13345
rect 46290 13336 46296 13388
rect 46348 13336 46354 13388
rect 46842 13336 46848 13388
rect 46900 13376 46906 13388
rect 47765 13379 47823 13385
rect 46900 13348 47532 13376
rect 46900 13336 46906 13348
rect 37642 13268 37648 13320
rect 37700 13308 37706 13320
rect 37700 13280 38056 13308
rect 37700 13268 37706 13280
rect 37016 13212 37412 13240
rect 37458 13200 37464 13252
rect 37516 13200 37522 13252
rect 37918 13200 37924 13252
rect 37976 13200 37982 13252
rect 38028 13240 38056 13280
rect 38562 13268 38568 13320
rect 38620 13308 38626 13320
rect 39150 13311 39208 13317
rect 39150 13308 39162 13311
rect 38620 13280 39162 13308
rect 38620 13268 38626 13280
rect 39150 13277 39162 13280
rect 39196 13277 39208 13311
rect 39150 13271 39208 13277
rect 39577 13311 39635 13317
rect 39577 13277 39589 13311
rect 39623 13308 39635 13311
rect 39758 13308 39764 13320
rect 39623 13280 39764 13308
rect 39623 13277 39635 13280
rect 39577 13271 39635 13277
rect 39758 13268 39764 13280
rect 39816 13268 39822 13320
rect 40037 13311 40095 13317
rect 40037 13277 40049 13311
rect 40083 13308 40095 13311
rect 41046 13308 41052 13320
rect 40083 13280 41052 13308
rect 40083 13277 40095 13280
rect 40037 13271 40095 13277
rect 41046 13268 41052 13280
rect 41104 13268 41110 13320
rect 44450 13268 44456 13320
rect 44508 13308 44514 13320
rect 45557 13311 45615 13317
rect 45557 13308 45569 13311
rect 44508 13280 45569 13308
rect 44508 13268 44514 13280
rect 45557 13277 45569 13280
rect 45603 13277 45615 13311
rect 45557 13271 45615 13277
rect 45649 13311 45707 13317
rect 45649 13277 45661 13311
rect 45695 13277 45707 13311
rect 45649 13271 45707 13277
rect 40310 13240 40316 13252
rect 38028 13212 40316 13240
rect 40310 13200 40316 13212
rect 40368 13200 40374 13252
rect 41506 13200 41512 13252
rect 41564 13240 41570 13252
rect 42061 13243 42119 13249
rect 42061 13240 42073 13243
rect 41564 13212 42073 13240
rect 41564 13200 41570 13212
rect 42061 13209 42073 13212
rect 42107 13209 42119 13243
rect 42061 13203 42119 13209
rect 19061 13175 19119 13181
rect 19061 13172 19073 13175
rect 18012 13144 19073 13172
rect 18012 13132 18018 13144
rect 19061 13141 19073 13144
rect 19107 13141 19119 13175
rect 19061 13135 19119 13141
rect 19242 13132 19248 13184
rect 19300 13132 19306 13184
rect 25501 13175 25559 13181
rect 25501 13141 25513 13175
rect 25547 13172 25559 13175
rect 26510 13172 26516 13184
rect 25547 13144 26516 13172
rect 25547 13141 25559 13144
rect 25501 13135 25559 13141
rect 26510 13132 26516 13144
rect 26568 13132 26574 13184
rect 30374 13132 30380 13184
rect 30432 13172 30438 13184
rect 31021 13175 31079 13181
rect 31021 13172 31033 13175
rect 30432 13144 31033 13172
rect 30432 13132 30438 13144
rect 31021 13141 31033 13144
rect 31067 13141 31079 13175
rect 31021 13135 31079 13141
rect 31662 13132 31668 13184
rect 31720 13172 31726 13184
rect 31941 13175 31999 13181
rect 31941 13172 31953 13175
rect 31720 13144 31953 13172
rect 31720 13132 31726 13144
rect 31941 13141 31953 13144
rect 31987 13141 31999 13175
rect 31941 13135 31999 13141
rect 36538 13132 36544 13184
rect 36596 13172 36602 13184
rect 37550 13172 37556 13184
rect 36596 13144 37556 13172
rect 36596 13132 36602 13144
rect 37550 13132 37556 13144
rect 37608 13132 37614 13184
rect 39206 13132 39212 13184
rect 39264 13132 39270 13184
rect 45373 13175 45431 13181
rect 45373 13141 45385 13175
rect 45419 13172 45431 13175
rect 45462 13172 45468 13184
rect 45419 13144 45468 13172
rect 45419 13141 45431 13144
rect 45373 13135 45431 13141
rect 45462 13132 45468 13144
rect 45520 13132 45526 13184
rect 45664 13172 45692 13271
rect 45922 13268 45928 13320
rect 45980 13268 45986 13320
rect 47504 13308 47532 13348
rect 47765 13345 47777 13379
rect 47811 13376 47823 13379
rect 48314 13376 48320 13388
rect 47811 13348 48320 13376
rect 47811 13345 47823 13348
rect 47765 13339 47823 13345
rect 48314 13336 48320 13348
rect 48372 13336 48378 13388
rect 49786 13336 49792 13388
rect 49844 13376 49850 13388
rect 50157 13379 50215 13385
rect 50157 13376 50169 13379
rect 49844 13348 50169 13376
rect 49844 13336 49850 13348
rect 50157 13345 50169 13348
rect 50203 13345 50215 13379
rect 50157 13339 50215 13345
rect 50433 13379 50491 13385
rect 50433 13345 50445 13379
rect 50479 13376 50491 13379
rect 51442 13376 51448 13388
rect 50479 13348 51448 13376
rect 50479 13345 50491 13348
rect 50433 13339 50491 13345
rect 51442 13336 51448 13348
rect 51500 13336 51506 13388
rect 48041 13311 48099 13317
rect 48041 13308 48053 13311
rect 47504 13280 48053 13308
rect 48041 13277 48053 13280
rect 48087 13277 48099 13311
rect 48041 13271 48099 13277
rect 48130 13268 48136 13320
rect 48188 13268 48194 13320
rect 48222 13268 48228 13320
rect 48280 13268 48286 13320
rect 48332 13308 48360 13336
rect 48409 13311 48467 13317
rect 48409 13308 48421 13311
rect 48332 13280 48421 13308
rect 48409 13277 48421 13280
rect 48455 13277 48467 13311
rect 48409 13271 48467 13277
rect 48682 13268 48688 13320
rect 48740 13308 48746 13320
rect 48961 13311 49019 13317
rect 48961 13308 48973 13311
rect 48740 13280 48973 13308
rect 48740 13268 48746 13280
rect 48961 13277 48973 13280
rect 49007 13308 49019 13311
rect 54588 13308 54616 13407
rect 55122 13336 55128 13388
rect 55180 13376 55186 13388
rect 55493 13379 55551 13385
rect 55493 13376 55505 13379
rect 55180 13348 55505 13376
rect 55180 13336 55186 13348
rect 55493 13345 55505 13348
rect 55539 13345 55551 13379
rect 55600 13376 55628 13416
rect 55769 13379 55827 13385
rect 55769 13376 55781 13379
rect 55600 13348 55781 13376
rect 55493 13339 55551 13345
rect 55769 13345 55781 13348
rect 55815 13345 55827 13379
rect 55769 13339 55827 13345
rect 54665 13311 54723 13317
rect 54665 13308 54677 13311
rect 49007 13280 50108 13308
rect 54588 13280 54677 13308
rect 49007 13277 49019 13280
rect 48961 13271 49019 13277
rect 47302 13200 47308 13252
rect 47360 13200 47366 13252
rect 47596 13212 47900 13240
rect 47596 13172 47624 13212
rect 47872 13181 47900 13212
rect 48498 13200 48504 13252
rect 48556 13240 48562 13252
rect 49053 13243 49111 13249
rect 49053 13240 49065 13243
rect 48556 13212 49065 13240
rect 48556 13200 48562 13212
rect 49053 13209 49065 13212
rect 49099 13209 49111 13243
rect 49053 13203 49111 13209
rect 45664 13144 47624 13172
rect 47857 13175 47915 13181
rect 47857 13141 47869 13175
rect 47903 13141 47915 13175
rect 50080 13172 50108 13280
rect 54665 13277 54677 13280
rect 54711 13277 54723 13311
rect 54665 13271 54723 13277
rect 54849 13311 54907 13317
rect 54849 13277 54861 13311
rect 54895 13277 54907 13311
rect 54849 13271 54907 13277
rect 50154 13200 50160 13252
rect 50212 13240 50218 13252
rect 54864 13240 54892 13271
rect 55674 13240 55680 13252
rect 50212 13212 50922 13240
rect 54864 13212 55680 13240
rect 50212 13200 50218 13212
rect 55674 13200 55680 13212
rect 55732 13200 55738 13252
rect 56778 13200 56784 13252
rect 56836 13200 56842 13252
rect 52270 13172 52276 13184
rect 50080 13144 52276 13172
rect 47857 13135 47915 13141
rect 52270 13132 52276 13144
rect 52328 13132 52334 13184
rect 57241 13175 57299 13181
rect 57241 13141 57253 13175
rect 57287 13172 57299 13175
rect 57422 13172 57428 13184
rect 57287 13144 57428 13172
rect 57287 13141 57299 13144
rect 57241 13135 57299 13141
rect 57422 13132 57428 13144
rect 57480 13132 57486 13184
rect 1104 13082 58880 13104
rect 1104 13030 4874 13082
rect 4926 13030 4938 13082
rect 4990 13030 5002 13082
rect 5054 13030 5066 13082
rect 5118 13030 5130 13082
rect 5182 13030 35594 13082
rect 35646 13030 35658 13082
rect 35710 13030 35722 13082
rect 35774 13030 35786 13082
rect 35838 13030 35850 13082
rect 35902 13030 58880 13082
rect 1104 13008 58880 13030
rect 16485 12971 16543 12977
rect 16485 12937 16497 12971
rect 16531 12968 16543 12971
rect 16574 12968 16580 12980
rect 16531 12940 16580 12968
rect 16531 12937 16543 12940
rect 16485 12931 16543 12937
rect 16574 12928 16580 12940
rect 16632 12928 16638 12980
rect 16850 12928 16856 12980
rect 16908 12928 16914 12980
rect 17218 12928 17224 12980
rect 17276 12968 17282 12980
rect 17589 12971 17647 12977
rect 17589 12968 17601 12971
rect 17276 12940 17601 12968
rect 17276 12928 17282 12940
rect 17589 12937 17601 12940
rect 17635 12937 17647 12971
rect 17589 12931 17647 12937
rect 23753 12971 23811 12977
rect 23753 12937 23765 12971
rect 23799 12968 23811 12971
rect 24394 12968 24400 12980
rect 23799 12940 24400 12968
rect 23799 12937 23811 12940
rect 23753 12931 23811 12937
rect 24394 12928 24400 12940
rect 24452 12928 24458 12980
rect 24578 12928 24584 12980
rect 24636 12968 24642 12980
rect 24636 12940 25544 12968
rect 24636 12928 24642 12940
rect 18414 12900 18420 12912
rect 17512 12872 18420 12900
rect 15378 12792 15384 12844
rect 15436 12832 15442 12844
rect 16025 12835 16083 12841
rect 16025 12832 16037 12835
rect 15436 12804 16037 12832
rect 15436 12792 15442 12804
rect 16025 12801 16037 12804
rect 16071 12832 16083 12835
rect 17310 12832 17316 12844
rect 16071 12804 17316 12832
rect 16071 12801 16083 12804
rect 16025 12795 16083 12801
rect 17310 12792 17316 12804
rect 17368 12792 17374 12844
rect 17512 12841 17540 12872
rect 18414 12860 18420 12872
rect 18472 12860 18478 12912
rect 18601 12903 18659 12909
rect 18601 12869 18613 12903
rect 18647 12900 18659 12903
rect 19242 12900 19248 12912
rect 18647 12872 19248 12900
rect 18647 12869 18659 12872
rect 18601 12863 18659 12869
rect 19242 12860 19248 12872
rect 19300 12860 19306 12912
rect 24210 12860 24216 12912
rect 24268 12860 24274 12912
rect 17497 12835 17555 12841
rect 17497 12801 17509 12835
rect 17543 12801 17555 12835
rect 18325 12835 18383 12841
rect 18325 12832 18337 12835
rect 17497 12795 17555 12801
rect 17880 12804 18337 12832
rect 16666 12724 16672 12776
rect 16724 12764 16730 12776
rect 17880 12764 17908 12804
rect 18325 12801 18337 12804
rect 18371 12832 18383 12835
rect 19613 12835 19671 12841
rect 19613 12832 19625 12835
rect 18371 12804 19625 12832
rect 18371 12801 18383 12804
rect 18325 12795 18383 12801
rect 19613 12801 19625 12804
rect 19659 12801 19671 12835
rect 19613 12795 19671 12801
rect 19794 12792 19800 12844
rect 19852 12792 19858 12844
rect 16724 12736 17908 12764
rect 18233 12767 18291 12773
rect 16724 12724 16730 12736
rect 18233 12733 18245 12767
rect 18279 12733 18291 12767
rect 18233 12727 18291 12733
rect 18248 12696 18276 12727
rect 21082 12724 21088 12776
rect 21140 12724 21146 12776
rect 24228 12764 24256 12860
rect 25516 12841 25544 12940
rect 25590 12928 25596 12980
rect 25648 12928 25654 12980
rect 26510 12928 26516 12980
rect 26568 12928 26574 12980
rect 27614 12928 27620 12980
rect 27672 12928 27678 12980
rect 30006 12968 30012 12980
rect 28644 12940 30012 12968
rect 26142 12860 26148 12912
rect 26200 12900 26206 12912
rect 26697 12903 26755 12909
rect 26697 12900 26709 12903
rect 26200 12872 26709 12900
rect 26200 12860 26206 12872
rect 25501 12835 25559 12841
rect 25501 12801 25513 12835
rect 25547 12801 25559 12835
rect 25501 12795 25559 12801
rect 25774 12792 25780 12844
rect 25832 12792 25838 12844
rect 25958 12792 25964 12844
rect 26016 12792 26022 12844
rect 26326 12792 26332 12844
rect 26384 12792 26390 12844
rect 26620 12841 26648 12872
rect 26697 12869 26709 12872
rect 26743 12869 26755 12903
rect 26697 12863 26755 12869
rect 26605 12835 26663 12841
rect 26605 12801 26617 12835
rect 26651 12832 26663 12835
rect 27709 12835 27767 12841
rect 26651 12804 26685 12832
rect 26651 12801 26663 12804
rect 26605 12795 26663 12801
rect 27709 12801 27721 12835
rect 27755 12832 27767 12835
rect 28537 12835 28595 12841
rect 28537 12832 28549 12835
rect 27755 12804 28549 12832
rect 27755 12801 27767 12804
rect 27709 12795 27767 12801
rect 28537 12801 28549 12804
rect 28583 12801 28595 12835
rect 28537 12795 28595 12801
rect 24762 12764 24768 12776
rect 24228 12736 24768 12764
rect 24762 12724 24768 12736
rect 24820 12724 24826 12776
rect 25225 12767 25283 12773
rect 25225 12733 25237 12767
rect 25271 12764 25283 12767
rect 26053 12767 26111 12773
rect 25271 12736 25728 12764
rect 25271 12733 25283 12736
rect 25225 12727 25283 12733
rect 18601 12699 18659 12705
rect 18601 12696 18613 12699
rect 18248 12668 18613 12696
rect 18601 12665 18613 12668
rect 18647 12665 18659 12699
rect 25700 12696 25728 12736
rect 26053 12733 26065 12767
rect 26099 12764 26111 12767
rect 26786 12764 26792 12776
rect 26099 12736 26792 12764
rect 26099 12733 26111 12736
rect 26053 12727 26111 12733
rect 26620 12708 26648 12736
rect 26786 12724 26792 12736
rect 26844 12724 26850 12776
rect 27893 12767 27951 12773
rect 27893 12733 27905 12767
rect 27939 12764 27951 12767
rect 28644 12764 28672 12940
rect 30006 12928 30012 12940
rect 30064 12928 30070 12980
rect 31110 12928 31116 12980
rect 31168 12968 31174 12980
rect 32125 12971 32183 12977
rect 32125 12968 32137 12971
rect 31168 12940 32137 12968
rect 31168 12928 31174 12940
rect 32125 12937 32137 12940
rect 32171 12937 32183 12971
rect 32125 12931 32183 12937
rect 32214 12928 32220 12980
rect 32272 12968 32278 12980
rect 32493 12971 32551 12977
rect 32493 12968 32505 12971
rect 32272 12940 32505 12968
rect 32272 12928 32278 12940
rect 32493 12937 32505 12940
rect 32539 12937 32551 12971
rect 32493 12931 32551 12937
rect 33042 12928 33048 12980
rect 33100 12968 33106 12980
rect 33321 12971 33379 12977
rect 33321 12968 33333 12971
rect 33100 12940 33333 12968
rect 33100 12928 33106 12940
rect 33321 12937 33333 12940
rect 33367 12937 33379 12971
rect 33321 12931 33379 12937
rect 33502 12928 33508 12980
rect 33560 12928 33566 12980
rect 36630 12928 36636 12980
rect 36688 12928 36694 12980
rect 37277 12971 37335 12977
rect 37277 12937 37289 12971
rect 37323 12968 37335 12971
rect 37734 12968 37740 12980
rect 37323 12940 37740 12968
rect 37323 12937 37335 12940
rect 37277 12931 37335 12937
rect 37734 12928 37740 12940
rect 37792 12928 37798 12980
rect 38562 12928 38568 12980
rect 38620 12928 38626 12980
rect 39206 12928 39212 12980
rect 39264 12968 39270 12980
rect 39301 12971 39359 12977
rect 39301 12968 39313 12971
rect 39264 12940 39313 12968
rect 39264 12928 39270 12940
rect 39301 12937 39313 12940
rect 39347 12937 39359 12971
rect 49786 12968 49792 12980
rect 39301 12931 39359 12937
rect 48792 12940 49792 12968
rect 28736 12872 32904 12900
rect 28736 12841 28764 12872
rect 28721 12835 28779 12841
rect 28721 12801 28733 12835
rect 28767 12801 28779 12835
rect 28721 12795 28779 12801
rect 28994 12792 29000 12844
rect 29052 12792 29058 12844
rect 29362 12792 29368 12844
rect 29420 12832 29426 12844
rect 29457 12835 29515 12841
rect 29457 12832 29469 12835
rect 29420 12804 29469 12832
rect 29420 12792 29426 12804
rect 29457 12801 29469 12804
rect 29503 12801 29515 12835
rect 29457 12795 29515 12801
rect 29638 12792 29644 12844
rect 29696 12792 29702 12844
rect 32309 12835 32367 12841
rect 32309 12801 32321 12835
rect 32355 12832 32367 12835
rect 32355 12804 32444 12832
rect 32355 12801 32367 12804
rect 32309 12795 32367 12801
rect 27939 12736 28672 12764
rect 28813 12767 28871 12773
rect 27939 12733 27951 12736
rect 27893 12727 27951 12733
rect 28813 12733 28825 12767
rect 28859 12764 28871 12767
rect 29178 12764 29184 12776
rect 28859 12736 29184 12764
rect 28859 12733 28871 12736
rect 28813 12727 28871 12733
rect 29178 12724 29184 12736
rect 29236 12724 29242 12776
rect 30282 12724 30288 12776
rect 30340 12764 30346 12776
rect 32416 12764 32444 12804
rect 32582 12792 32588 12844
rect 32640 12792 32646 12844
rect 32876 12773 32904 12872
rect 33410 12860 33416 12912
rect 33468 12900 33474 12912
rect 39117 12903 39175 12909
rect 33468 12872 39068 12900
rect 33468 12860 33474 12872
rect 33324 12835 33382 12841
rect 33324 12801 33336 12835
rect 33370 12832 33382 12835
rect 33502 12832 33508 12844
rect 33370 12804 33508 12832
rect 33370 12801 33382 12804
rect 33324 12795 33382 12801
rect 33502 12792 33508 12804
rect 33560 12832 33566 12844
rect 36262 12832 36268 12844
rect 33560 12804 36268 12832
rect 33560 12792 33566 12804
rect 36262 12792 36268 12804
rect 36320 12792 36326 12844
rect 36541 12835 36599 12841
rect 36541 12801 36553 12835
rect 36587 12832 36599 12835
rect 36814 12832 36820 12844
rect 36587 12804 36820 12832
rect 36587 12801 36599 12804
rect 36541 12795 36599 12801
rect 36814 12792 36820 12804
rect 36872 12792 36878 12844
rect 36998 12792 37004 12844
rect 37056 12792 37062 12844
rect 37461 12835 37519 12841
rect 37461 12801 37473 12835
rect 37507 12801 37519 12835
rect 37461 12795 37519 12801
rect 30340 12736 32444 12764
rect 30340 12724 30346 12736
rect 26145 12699 26203 12705
rect 26145 12696 26157 12699
rect 25700 12668 26157 12696
rect 18601 12659 18659 12665
rect 26145 12665 26157 12668
rect 26191 12665 26203 12699
rect 26145 12659 26203 12665
rect 26602 12656 26608 12708
rect 26660 12656 26666 12708
rect 28905 12699 28963 12705
rect 28905 12665 28917 12699
rect 28951 12696 28963 12699
rect 29546 12696 29552 12708
rect 28951 12668 29552 12696
rect 28951 12665 28963 12668
rect 28905 12659 28963 12665
rect 29546 12656 29552 12668
rect 29604 12656 29610 12708
rect 32416 12696 32444 12736
rect 32861 12767 32919 12773
rect 32861 12733 32873 12767
rect 32907 12764 32919 12767
rect 33134 12764 33140 12776
rect 32907 12736 33140 12764
rect 32907 12733 32919 12736
rect 32861 12727 32919 12733
rect 33134 12724 33140 12736
rect 33192 12724 33198 12776
rect 36832 12764 36860 12792
rect 37090 12764 37096 12776
rect 36832 12736 37096 12764
rect 37090 12724 37096 12736
rect 37148 12724 37154 12776
rect 37476 12764 37504 12795
rect 37642 12792 37648 12844
rect 37700 12792 37706 12844
rect 38470 12792 38476 12844
rect 38528 12792 38534 12844
rect 38746 12792 38752 12844
rect 38804 12792 38810 12844
rect 38838 12792 38844 12844
rect 38896 12792 38902 12844
rect 39040 12841 39068 12872
rect 39117 12869 39129 12903
rect 39163 12900 39175 12903
rect 40586 12900 40592 12912
rect 39163 12872 40592 12900
rect 39163 12869 39175 12872
rect 39117 12863 39175 12869
rect 40586 12860 40592 12872
rect 40644 12860 40650 12912
rect 45462 12860 45468 12912
rect 45520 12860 45526 12912
rect 46750 12900 46756 12912
rect 46690 12872 46756 12900
rect 46750 12860 46756 12872
rect 46808 12900 46814 12912
rect 47302 12900 47308 12912
rect 46808 12872 47308 12900
rect 46808 12860 46814 12872
rect 47302 12860 47308 12872
rect 47360 12860 47366 12912
rect 39025 12835 39083 12841
rect 39025 12801 39037 12835
rect 39071 12801 39083 12835
rect 39025 12795 39083 12801
rect 39209 12835 39267 12841
rect 39209 12801 39221 12835
rect 39255 12801 39267 12835
rect 39209 12795 39267 12801
rect 37734 12764 37740 12776
rect 37476 12736 37740 12764
rect 37734 12724 37740 12736
rect 37792 12724 37798 12776
rect 38654 12724 38660 12776
rect 38712 12764 38718 12776
rect 39114 12764 39120 12776
rect 38712 12736 39120 12764
rect 38712 12724 38718 12736
rect 39114 12724 39120 12736
rect 39172 12724 39178 12776
rect 39224 12764 39252 12795
rect 39298 12792 39304 12844
rect 39356 12832 39362 12844
rect 39393 12835 39451 12841
rect 39393 12832 39405 12835
rect 39356 12804 39405 12832
rect 39356 12792 39362 12804
rect 39393 12801 39405 12804
rect 39439 12801 39451 12835
rect 39393 12795 39451 12801
rect 39485 12835 39543 12841
rect 39485 12801 39497 12835
rect 39531 12832 39543 12835
rect 39574 12832 39580 12844
rect 39531 12804 39580 12832
rect 39531 12801 39543 12804
rect 39485 12795 39543 12801
rect 39408 12764 39436 12795
rect 39574 12792 39580 12804
rect 39632 12792 39638 12844
rect 42797 12835 42855 12841
rect 42797 12801 42809 12835
rect 42843 12832 42855 12835
rect 43625 12835 43683 12841
rect 43625 12832 43637 12835
rect 42843 12804 43637 12832
rect 42843 12801 42855 12804
rect 42797 12795 42855 12801
rect 43625 12801 43637 12804
rect 43671 12801 43683 12835
rect 43625 12795 43683 12801
rect 44910 12792 44916 12844
rect 44968 12832 44974 12844
rect 45189 12835 45247 12841
rect 45189 12832 45201 12835
rect 44968 12804 45201 12832
rect 44968 12792 44974 12804
rect 45189 12801 45201 12804
rect 45235 12801 45247 12835
rect 47320 12832 47348 12860
rect 48792 12841 48820 12940
rect 49786 12928 49792 12940
rect 49844 12928 49850 12980
rect 50522 12928 50528 12980
rect 50580 12928 50586 12980
rect 57606 12928 57612 12980
rect 57664 12928 57670 12980
rect 49050 12860 49056 12912
rect 49108 12860 49114 12912
rect 48777 12835 48835 12841
rect 47320 12804 48728 12832
rect 45189 12795 45247 12801
rect 39942 12764 39948 12776
rect 39224 12736 39344 12764
rect 39408 12736 39948 12764
rect 33042 12696 33048 12708
rect 32416 12668 33048 12696
rect 33042 12656 33048 12668
rect 33100 12656 33106 12708
rect 33686 12656 33692 12708
rect 33744 12696 33750 12708
rect 33744 12668 36032 12696
rect 33744 12656 33750 12668
rect 19610 12588 19616 12640
rect 19668 12588 19674 12640
rect 19702 12588 19708 12640
rect 19760 12628 19766 12640
rect 20441 12631 20499 12637
rect 20441 12628 20453 12631
rect 19760 12600 20453 12628
rect 19760 12588 19766 12600
rect 20441 12597 20453 12600
rect 20487 12597 20499 12631
rect 20441 12591 20499 12597
rect 27246 12588 27252 12640
rect 27304 12588 27310 12640
rect 29641 12631 29699 12637
rect 29641 12597 29653 12631
rect 29687 12628 29699 12631
rect 30466 12628 30472 12640
rect 29687 12600 30472 12628
rect 29687 12597 29699 12600
rect 29641 12591 29699 12597
rect 30466 12588 30472 12600
rect 30524 12588 30530 12640
rect 32953 12631 33011 12637
rect 32953 12597 32965 12631
rect 32999 12628 33011 12631
rect 33226 12628 33232 12640
rect 32999 12600 33232 12628
rect 32999 12597 33011 12600
rect 32953 12591 33011 12597
rect 33226 12588 33232 12600
rect 33284 12588 33290 12640
rect 36004 12628 36032 12668
rect 37918 12656 37924 12708
rect 37976 12696 37982 12708
rect 39316 12696 39344 12736
rect 39942 12724 39948 12736
rect 40000 12724 40006 12776
rect 42886 12724 42892 12776
rect 42944 12724 42950 12776
rect 42981 12767 43039 12773
rect 42981 12733 42993 12767
rect 43027 12733 43039 12767
rect 42981 12727 43039 12733
rect 37976 12668 39344 12696
rect 37976 12656 37982 12668
rect 39758 12656 39764 12708
rect 39816 12696 39822 12708
rect 42996 12696 43024 12727
rect 44266 12724 44272 12776
rect 44324 12764 44330 12776
rect 48130 12764 48136 12776
rect 44324 12736 48136 12764
rect 44324 12724 44330 12736
rect 48130 12724 48136 12736
rect 48188 12724 48194 12776
rect 48700 12764 48728 12804
rect 48777 12801 48789 12835
rect 48823 12801 48835 12835
rect 48777 12795 48835 12801
rect 50154 12792 50160 12844
rect 50212 12792 50218 12844
rect 57422 12792 57428 12844
rect 57480 12792 57486 12844
rect 50172 12764 50200 12792
rect 48700 12736 50200 12764
rect 39816 12668 43024 12696
rect 39816 12656 39822 12668
rect 39776 12628 39804 12656
rect 36004 12600 39804 12628
rect 42429 12631 42487 12637
rect 42429 12597 42441 12631
rect 42475 12628 42487 12631
rect 42794 12628 42800 12640
rect 42475 12600 42800 12628
rect 42475 12597 42487 12600
rect 42429 12591 42487 12597
rect 42794 12588 42800 12600
rect 42852 12588 42858 12640
rect 45922 12588 45928 12640
rect 45980 12628 45986 12640
rect 46566 12628 46572 12640
rect 45980 12600 46572 12628
rect 45980 12588 45986 12600
rect 46566 12588 46572 12600
rect 46624 12628 46630 12640
rect 46937 12631 46995 12637
rect 46937 12628 46949 12631
rect 46624 12600 46949 12628
rect 46624 12588 46630 12600
rect 46937 12597 46949 12600
rect 46983 12597 46995 12631
rect 46937 12591 46995 12597
rect 1104 12538 58880 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 58880 12538
rect 1104 12464 58880 12486
rect 15378 12424 15384 12436
rect 13832 12396 15384 12424
rect 12158 12248 12164 12300
rect 12216 12288 12222 12300
rect 13832 12288 13860 12396
rect 15378 12384 15384 12396
rect 15436 12384 15442 12436
rect 17034 12384 17040 12436
rect 17092 12424 17098 12436
rect 17221 12427 17279 12433
rect 17221 12424 17233 12427
rect 17092 12396 17233 12424
rect 17092 12384 17098 12396
rect 17221 12393 17233 12396
rect 17267 12393 17279 12427
rect 18325 12427 18383 12433
rect 17221 12387 17279 12393
rect 17696 12396 18276 12424
rect 13909 12359 13967 12365
rect 13909 12325 13921 12359
rect 13955 12356 13967 12359
rect 13955 12328 14780 12356
rect 13955 12325 13967 12328
rect 13909 12319 13967 12325
rect 14752 12300 14780 12328
rect 12216 12260 13860 12288
rect 12216 12248 12222 12260
rect 14734 12248 14740 12300
rect 14792 12248 14798 12300
rect 15396 12297 15424 12384
rect 15381 12291 15439 12297
rect 15381 12257 15393 12291
rect 15427 12257 15439 12291
rect 15381 12251 15439 12257
rect 15654 12248 15660 12300
rect 15712 12248 15718 12300
rect 17129 12291 17187 12297
rect 17129 12257 17141 12291
rect 17175 12288 17187 12291
rect 17696 12288 17724 12396
rect 17773 12359 17831 12365
rect 17773 12325 17785 12359
rect 17819 12356 17831 12359
rect 17954 12356 17960 12368
rect 17819 12328 17960 12356
rect 17819 12325 17831 12328
rect 17773 12319 17831 12325
rect 17954 12316 17960 12328
rect 18012 12356 18018 12368
rect 18012 12328 18184 12356
rect 18012 12316 18018 12328
rect 18156 12297 18184 12328
rect 17175 12260 17724 12288
rect 17175 12257 17187 12260
rect 17129 12251 17187 12257
rect 14826 12180 14832 12232
rect 14884 12180 14890 12232
rect 15013 12223 15071 12229
rect 15013 12189 15025 12223
rect 15059 12220 15071 12223
rect 15286 12220 15292 12232
rect 15059 12192 15292 12220
rect 15059 12189 15071 12192
rect 15013 12183 15071 12189
rect 15286 12180 15292 12192
rect 15344 12180 15350 12232
rect 16758 12180 16764 12232
rect 16816 12180 16822 12232
rect 17589 12223 17647 12229
rect 17589 12189 17601 12223
rect 17635 12220 17647 12223
rect 17696 12220 17724 12260
rect 18141 12291 18199 12297
rect 18141 12257 18153 12291
rect 18187 12257 18199 12291
rect 18141 12251 18199 12257
rect 17635 12192 17724 12220
rect 18049 12223 18107 12229
rect 17635 12189 17647 12192
rect 17589 12183 17647 12189
rect 18049 12189 18061 12223
rect 18095 12222 18107 12223
rect 18095 12194 18184 12222
rect 18095 12189 18107 12194
rect 18049 12183 18107 12189
rect 12437 12155 12495 12161
rect 12437 12121 12449 12155
rect 12483 12121 12495 12155
rect 12437 12115 12495 12121
rect 12452 12084 12480 12115
rect 13446 12112 13452 12164
rect 13504 12112 13510 12164
rect 14921 12155 14979 12161
rect 14921 12152 14933 12155
rect 13740 12124 14933 12152
rect 13740 12084 13768 12124
rect 14921 12121 14933 12124
rect 14967 12121 14979 12155
rect 14921 12115 14979 12121
rect 16942 12112 16948 12164
rect 17000 12152 17006 12164
rect 17405 12155 17463 12161
rect 17405 12152 17417 12155
rect 17000 12124 17417 12152
rect 17000 12112 17006 12124
rect 17405 12121 17417 12124
rect 17451 12152 17463 12155
rect 18156 12152 18184 12194
rect 18248 12220 18276 12396
rect 18325 12393 18337 12427
rect 18371 12393 18383 12427
rect 18325 12387 18383 12393
rect 19521 12427 19579 12433
rect 19521 12393 19533 12427
rect 19567 12424 19579 12427
rect 19794 12424 19800 12436
rect 19567 12396 19800 12424
rect 19567 12393 19579 12396
rect 19521 12387 19579 12393
rect 18340 12288 18368 12387
rect 19794 12384 19800 12396
rect 19852 12384 19858 12436
rect 24854 12384 24860 12436
rect 24912 12424 24918 12436
rect 26605 12427 26663 12433
rect 24912 12396 26556 12424
rect 24912 12384 24918 12396
rect 19242 12316 19248 12368
rect 19300 12356 19306 12368
rect 19300 12328 19932 12356
rect 19300 12316 19306 12328
rect 19904 12297 19932 12328
rect 26326 12316 26332 12368
rect 26384 12356 26390 12368
rect 26421 12359 26479 12365
rect 26421 12356 26433 12359
rect 26384 12328 26433 12356
rect 26384 12316 26390 12328
rect 26421 12325 26433 12328
rect 26467 12325 26479 12359
rect 26528 12356 26556 12396
rect 26605 12393 26617 12427
rect 26651 12424 26663 12427
rect 26786 12424 26792 12436
rect 26651 12396 26792 12424
rect 26651 12393 26663 12396
rect 26605 12387 26663 12393
rect 26786 12384 26792 12396
rect 26844 12384 26850 12436
rect 27982 12384 27988 12436
rect 28040 12384 28046 12436
rect 28994 12384 29000 12436
rect 29052 12424 29058 12436
rect 29549 12427 29607 12433
rect 29549 12424 29561 12427
rect 29052 12396 29561 12424
rect 29052 12384 29058 12396
rect 29549 12393 29561 12396
rect 29595 12393 29607 12427
rect 29549 12387 29607 12393
rect 29730 12384 29736 12436
rect 29788 12424 29794 12436
rect 30285 12427 30343 12433
rect 30285 12424 30297 12427
rect 29788 12396 30297 12424
rect 29788 12384 29794 12396
rect 30285 12393 30297 12396
rect 30331 12393 30343 12427
rect 30285 12387 30343 12393
rect 30469 12427 30527 12433
rect 30469 12393 30481 12427
rect 30515 12393 30527 12427
rect 30469 12387 30527 12393
rect 26878 12356 26884 12368
rect 26528 12328 26884 12356
rect 26421 12319 26479 12325
rect 26878 12316 26884 12328
rect 26936 12356 26942 12368
rect 26973 12359 27031 12365
rect 26973 12356 26985 12359
rect 26936 12328 26985 12356
rect 26936 12316 26942 12328
rect 26973 12325 26985 12328
rect 27019 12325 27031 12359
rect 26973 12319 27031 12325
rect 28629 12359 28687 12365
rect 28629 12325 28641 12359
rect 28675 12356 28687 12359
rect 30484 12356 30512 12387
rect 31662 12384 31668 12436
rect 31720 12384 31726 12436
rect 32582 12424 32588 12436
rect 32416 12396 32588 12424
rect 32416 12356 32444 12396
rect 32582 12384 32588 12396
rect 32640 12384 32646 12436
rect 33134 12384 33140 12436
rect 33192 12424 33198 12436
rect 33505 12427 33563 12433
rect 33505 12424 33517 12427
rect 33192 12396 33517 12424
rect 33192 12384 33198 12396
rect 33505 12393 33517 12396
rect 33551 12393 33563 12427
rect 33505 12387 33563 12393
rect 33778 12384 33784 12436
rect 33836 12424 33842 12436
rect 35710 12424 35716 12436
rect 33836 12396 35716 12424
rect 33836 12384 33842 12396
rect 35710 12384 35716 12396
rect 35768 12424 35774 12436
rect 37642 12424 37648 12436
rect 35768 12396 37648 12424
rect 35768 12384 35774 12396
rect 37642 12384 37648 12396
rect 37700 12384 37706 12436
rect 37734 12384 37740 12436
rect 37792 12424 37798 12436
rect 39666 12424 39672 12436
rect 37792 12396 39672 12424
rect 37792 12384 37798 12396
rect 39666 12384 39672 12396
rect 39724 12384 39730 12436
rect 40862 12384 40868 12436
rect 40920 12424 40926 12436
rect 43441 12427 43499 12433
rect 43441 12424 43453 12427
rect 40920 12396 43453 12424
rect 40920 12384 40926 12396
rect 43441 12393 43453 12396
rect 43487 12424 43499 12427
rect 43714 12424 43720 12436
rect 43487 12396 43720 12424
rect 43487 12393 43499 12396
rect 43441 12387 43499 12393
rect 43714 12384 43720 12396
rect 43772 12384 43778 12436
rect 46198 12384 46204 12436
rect 46256 12384 46262 12436
rect 46661 12427 46719 12433
rect 46661 12393 46673 12427
rect 46707 12424 46719 12427
rect 46750 12424 46756 12436
rect 46707 12396 46756 12424
rect 46707 12393 46719 12396
rect 46661 12387 46719 12393
rect 46750 12384 46756 12396
rect 46808 12384 46814 12436
rect 28675 12328 30512 12356
rect 30576 12328 32444 12356
rect 28675 12325 28687 12328
rect 28629 12319 28687 12325
rect 19889 12291 19947 12297
rect 18340 12260 19380 12288
rect 18325 12223 18383 12229
rect 18325 12220 18337 12223
rect 18248 12192 18337 12220
rect 18325 12189 18337 12192
rect 18371 12220 18383 12223
rect 18414 12220 18420 12232
rect 18371 12192 18420 12220
rect 18371 12189 18383 12192
rect 18325 12183 18383 12189
rect 18414 12180 18420 12192
rect 18472 12180 18478 12232
rect 18616 12229 18644 12260
rect 18601 12223 18659 12229
rect 18601 12189 18613 12223
rect 18647 12189 18659 12223
rect 18601 12183 18659 12189
rect 18785 12223 18843 12229
rect 18785 12189 18797 12223
rect 18831 12189 18843 12223
rect 18785 12183 18843 12189
rect 18800 12152 18828 12183
rect 19242 12180 19248 12232
rect 19300 12180 19306 12232
rect 19352 12229 19380 12260
rect 19889 12257 19901 12291
rect 19935 12257 19947 12291
rect 19889 12251 19947 12257
rect 20165 12291 20223 12297
rect 20165 12257 20177 12291
rect 20211 12288 20223 12291
rect 22465 12291 22523 12297
rect 22465 12288 22477 12291
rect 20211 12260 22477 12288
rect 20211 12257 20223 12260
rect 20165 12251 20223 12257
rect 22465 12257 22477 12260
rect 22511 12257 22523 12291
rect 22465 12251 22523 12257
rect 22741 12291 22799 12297
rect 22741 12257 22753 12291
rect 22787 12288 22799 12291
rect 24578 12288 24584 12300
rect 22787 12260 24584 12288
rect 22787 12257 22799 12260
rect 22741 12251 22799 12257
rect 24578 12248 24584 12260
rect 24636 12248 24642 12300
rect 24857 12291 24915 12297
rect 24857 12257 24869 12291
rect 24903 12288 24915 12291
rect 26694 12288 26700 12300
rect 24903 12260 26700 12288
rect 24903 12257 24915 12260
rect 24857 12251 24915 12257
rect 26694 12248 26700 12260
rect 26752 12248 26758 12300
rect 27338 12248 27344 12300
rect 27396 12288 27402 12300
rect 29733 12291 29791 12297
rect 29733 12288 29745 12291
rect 27396 12260 27844 12288
rect 27396 12248 27402 12260
rect 19337 12223 19395 12229
rect 19337 12189 19349 12223
rect 19383 12189 19395 12223
rect 19337 12183 19395 12189
rect 19521 12223 19579 12229
rect 19521 12189 19533 12223
rect 19567 12220 19579 12223
rect 19702 12220 19708 12232
rect 19567 12192 19708 12220
rect 19567 12189 19579 12192
rect 19521 12183 19579 12189
rect 17451 12124 18000 12152
rect 18156 12124 18828 12152
rect 19352 12152 19380 12183
rect 19702 12180 19708 12192
rect 19760 12180 19766 12232
rect 19797 12223 19855 12229
rect 19797 12189 19809 12223
rect 19843 12220 19855 12223
rect 20257 12223 20315 12229
rect 20257 12220 20269 12223
rect 19843 12192 20269 12220
rect 19843 12189 19855 12192
rect 19797 12183 19855 12189
rect 20257 12189 20269 12192
rect 20303 12189 20315 12223
rect 20257 12183 20315 12189
rect 20809 12223 20867 12229
rect 20809 12189 20821 12223
rect 20855 12189 20867 12223
rect 20809 12183 20867 12189
rect 20824 12152 20852 12183
rect 26602 12180 26608 12232
rect 26660 12220 26666 12232
rect 26660 12192 26832 12220
rect 26660 12180 26666 12192
rect 22186 12152 22192 12164
rect 19352 12124 21036 12152
rect 22034 12124 22192 12152
rect 17451 12121 17463 12124
rect 17405 12115 17463 12121
rect 12452 12056 13768 12084
rect 14090 12044 14096 12096
rect 14148 12044 14154 12096
rect 15286 12044 15292 12096
rect 15344 12084 15350 12096
rect 17494 12084 17500 12096
rect 15344 12056 17500 12084
rect 15344 12044 15350 12056
rect 17494 12044 17500 12056
rect 17552 12044 17558 12096
rect 17862 12044 17868 12096
rect 17920 12044 17926 12096
rect 17972 12084 18000 12124
rect 18417 12087 18475 12093
rect 18417 12084 18429 12087
rect 17972 12056 18429 12084
rect 18417 12053 18429 12056
rect 18463 12053 18475 12087
rect 18800 12084 18828 12124
rect 20898 12084 20904 12096
rect 18800 12056 20904 12084
rect 18417 12047 18475 12053
rect 20898 12044 20904 12056
rect 20956 12044 20962 12096
rect 21008 12093 21036 12124
rect 22186 12112 22192 12124
rect 22244 12112 22250 12164
rect 26804 12161 26832 12192
rect 27154 12180 27160 12232
rect 27212 12180 27218 12232
rect 27816 12229 27844 12260
rect 28000 12260 28948 12288
rect 28000 12229 28028 12260
rect 28920 12232 28948 12260
rect 29288 12260 29745 12288
rect 27801 12223 27859 12229
rect 27801 12189 27813 12223
rect 27847 12189 27859 12223
rect 27801 12183 27859 12189
rect 27985 12223 28043 12229
rect 27985 12189 27997 12223
rect 28031 12189 28043 12223
rect 27985 12183 28043 12189
rect 28718 12180 28724 12232
rect 28776 12220 28782 12232
rect 28813 12223 28871 12229
rect 28813 12220 28825 12223
rect 28776 12192 28825 12220
rect 28776 12180 28782 12192
rect 28813 12189 28825 12192
rect 28859 12189 28871 12223
rect 28813 12183 28871 12189
rect 28902 12180 28908 12232
rect 28960 12180 28966 12232
rect 29288 12229 29316 12260
rect 29733 12257 29745 12260
rect 29779 12288 29791 12291
rect 30576 12288 30604 12328
rect 32674 12316 32680 12368
rect 32732 12356 32738 12368
rect 37752 12356 37780 12384
rect 32732 12328 37780 12356
rect 32732 12316 32738 12328
rect 32953 12291 33011 12297
rect 32953 12288 32965 12291
rect 29779 12260 30604 12288
rect 30668 12260 32965 12288
rect 29779 12257 29791 12260
rect 29733 12251 29791 12257
rect 28997 12223 29055 12229
rect 28997 12189 29009 12223
rect 29043 12189 29055 12223
rect 28997 12183 29055 12189
rect 29089 12223 29147 12229
rect 29089 12189 29101 12223
rect 29135 12189 29147 12223
rect 29089 12183 29147 12189
rect 29273 12223 29331 12229
rect 29273 12189 29285 12223
rect 29319 12189 29331 12223
rect 29273 12183 29331 12189
rect 29825 12223 29883 12229
rect 29825 12189 29837 12223
rect 29871 12220 29883 12223
rect 30374 12220 30380 12232
rect 29871 12192 30380 12220
rect 29871 12189 29883 12192
rect 29825 12183 29883 12189
rect 26789 12155 26847 12161
rect 24964 12124 25346 12152
rect 20993 12087 21051 12093
rect 20993 12053 21005 12087
rect 21039 12053 21051 12087
rect 20993 12047 21051 12053
rect 24762 12044 24768 12096
rect 24820 12084 24826 12096
rect 24964 12084 24992 12124
rect 26789 12121 26801 12155
rect 26835 12121 26847 12155
rect 29012 12152 29040 12183
rect 26789 12115 26847 12121
rect 27632 12124 29040 12152
rect 29104 12152 29132 12183
rect 29840 12152 29868 12183
rect 30374 12180 30380 12192
rect 30432 12180 30438 12232
rect 30466 12180 30472 12232
rect 30524 12180 30530 12232
rect 30558 12180 30564 12232
rect 30616 12180 30622 12232
rect 29104 12124 29868 12152
rect 27632 12096 27660 12124
rect 29914 12112 29920 12164
rect 29972 12152 29978 12164
rect 30668 12152 30696 12260
rect 32953 12257 32965 12260
rect 32999 12257 33011 12291
rect 32953 12251 33011 12257
rect 31478 12180 31484 12232
rect 31536 12180 31542 12232
rect 31754 12180 31760 12232
rect 31812 12180 31818 12232
rect 33042 12180 33048 12232
rect 33100 12180 33106 12232
rect 33152 12229 33180 12328
rect 38654 12316 38660 12368
rect 38712 12316 38718 12368
rect 40236 12328 41828 12356
rect 34238 12288 34244 12300
rect 33244 12260 34244 12288
rect 33244 12229 33272 12260
rect 34238 12248 34244 12260
rect 34296 12248 34302 12300
rect 38672 12288 38700 12316
rect 34532 12260 38700 12288
rect 33137 12223 33195 12229
rect 33137 12189 33149 12223
rect 33183 12189 33195 12223
rect 33137 12183 33195 12189
rect 33229 12223 33287 12229
rect 33229 12189 33241 12223
rect 33275 12189 33287 12223
rect 33229 12183 33287 12189
rect 33318 12180 33324 12232
rect 33376 12220 33382 12232
rect 33413 12223 33471 12229
rect 33413 12220 33425 12223
rect 33376 12192 33425 12220
rect 33376 12180 33382 12192
rect 33413 12189 33425 12192
rect 33459 12189 33471 12223
rect 33413 12183 33471 12189
rect 33686 12180 33692 12232
rect 33744 12180 33750 12232
rect 33778 12180 33784 12232
rect 33836 12180 33842 12232
rect 33873 12223 33931 12229
rect 33873 12189 33885 12223
rect 33919 12189 33931 12223
rect 33873 12183 33931 12189
rect 29972 12124 30696 12152
rect 30745 12155 30803 12161
rect 29972 12112 29978 12124
rect 30745 12121 30757 12155
rect 30791 12121 30803 12155
rect 30745 12115 30803 12121
rect 24820 12056 24992 12084
rect 24820 12044 24826 12056
rect 26234 12044 26240 12096
rect 26292 12084 26298 12096
rect 26329 12087 26387 12093
rect 26329 12084 26341 12087
rect 26292 12056 26341 12084
rect 26292 12044 26298 12056
rect 26329 12053 26341 12056
rect 26375 12053 26387 12087
rect 26329 12047 26387 12053
rect 26589 12087 26647 12093
rect 26589 12053 26601 12087
rect 26635 12084 26647 12087
rect 26878 12084 26884 12096
rect 26635 12056 26884 12084
rect 26635 12053 26647 12056
rect 26589 12047 26647 12053
rect 26878 12044 26884 12056
rect 26936 12044 26942 12096
rect 26970 12044 26976 12096
rect 27028 12084 27034 12096
rect 27249 12087 27307 12093
rect 27249 12084 27261 12087
rect 27028 12056 27261 12084
rect 27028 12044 27034 12056
rect 27249 12053 27261 12056
rect 27295 12053 27307 12087
rect 27249 12047 27307 12053
rect 27614 12044 27620 12096
rect 27672 12044 27678 12096
rect 29454 12044 29460 12096
rect 29512 12084 29518 12096
rect 30193 12087 30251 12093
rect 30193 12084 30205 12087
rect 29512 12056 30205 12084
rect 29512 12044 29518 12056
rect 30193 12053 30205 12056
rect 30239 12084 30251 12087
rect 30282 12084 30288 12096
rect 30239 12056 30288 12084
rect 30239 12053 30251 12056
rect 30193 12047 30251 12053
rect 30282 12044 30288 12056
rect 30340 12044 30346 12096
rect 30760 12084 30788 12115
rect 31018 12112 31024 12164
rect 31076 12152 31082 12164
rect 33888 12152 33916 12183
rect 33962 12180 33968 12232
rect 34020 12220 34026 12232
rect 34422 12220 34428 12232
rect 34020 12192 34428 12220
rect 34020 12180 34026 12192
rect 34422 12180 34428 12192
rect 34480 12180 34486 12232
rect 34532 12152 34560 12260
rect 34882 12180 34888 12232
rect 34940 12180 34946 12232
rect 34977 12223 35035 12229
rect 34977 12189 34989 12223
rect 35023 12189 35035 12223
rect 34977 12183 35035 12189
rect 31076 12124 34560 12152
rect 34992 12152 35020 12183
rect 35158 12180 35164 12232
rect 35216 12180 35222 12232
rect 35253 12223 35311 12229
rect 35253 12189 35265 12223
rect 35299 12220 35311 12223
rect 35434 12220 35440 12232
rect 35299 12192 35440 12220
rect 35299 12189 35311 12192
rect 35253 12183 35311 12189
rect 35434 12180 35440 12192
rect 35492 12180 35498 12232
rect 35710 12229 35716 12232
rect 35708 12220 35716 12229
rect 35671 12192 35716 12220
rect 35708 12183 35716 12192
rect 35710 12180 35716 12183
rect 35768 12180 35774 12232
rect 35805 12223 35863 12229
rect 35805 12189 35817 12223
rect 35851 12220 35863 12223
rect 35986 12220 35992 12232
rect 35851 12192 35992 12220
rect 35851 12189 35863 12192
rect 35805 12183 35863 12189
rect 35986 12180 35992 12192
rect 36044 12180 36050 12232
rect 36080 12223 36138 12229
rect 36080 12189 36092 12223
rect 36126 12189 36138 12223
rect 36080 12183 36138 12189
rect 36173 12223 36231 12229
rect 36173 12189 36185 12223
rect 36219 12220 36231 12223
rect 36219 12192 37412 12220
rect 36219 12189 36231 12192
rect 36173 12183 36231 12189
rect 35897 12155 35955 12161
rect 34992 12124 35572 12152
rect 31076 12112 31082 12124
rect 31205 12087 31263 12093
rect 31205 12084 31217 12087
rect 30760 12056 31217 12084
rect 31205 12053 31217 12056
rect 31251 12053 31263 12087
rect 31205 12047 31263 12053
rect 32582 12044 32588 12096
rect 32640 12084 32646 12096
rect 32677 12087 32735 12093
rect 32677 12084 32689 12087
rect 32640 12056 32689 12084
rect 32640 12044 32646 12056
rect 32677 12053 32689 12056
rect 32723 12053 32735 12087
rect 32677 12047 32735 12053
rect 35342 12044 35348 12096
rect 35400 12084 35406 12096
rect 35544 12093 35572 12124
rect 35897 12121 35909 12155
rect 35943 12152 35955 12155
rect 36095 12152 36123 12183
rect 36262 12152 36268 12164
rect 35943 12124 36032 12152
rect 36095 12124 36268 12152
rect 35943 12121 35955 12124
rect 35897 12115 35955 12121
rect 36004 12096 36032 12124
rect 36262 12112 36268 12124
rect 36320 12112 36326 12164
rect 37384 12152 37412 12192
rect 37826 12180 37832 12232
rect 37884 12220 37890 12232
rect 38657 12223 38715 12229
rect 38657 12220 38669 12223
rect 37884 12192 38669 12220
rect 37884 12180 37890 12192
rect 38657 12189 38669 12192
rect 38703 12189 38715 12223
rect 38657 12183 38715 12189
rect 38746 12180 38752 12232
rect 38804 12220 38810 12232
rect 39025 12223 39083 12229
rect 39025 12220 39037 12223
rect 38804 12192 39037 12220
rect 38804 12180 38810 12192
rect 39025 12189 39037 12192
rect 39071 12189 39083 12223
rect 39025 12183 39083 12189
rect 39206 12180 39212 12232
rect 39264 12180 39270 12232
rect 39482 12180 39488 12232
rect 39540 12220 39546 12232
rect 39853 12223 39911 12229
rect 39853 12220 39865 12223
rect 39540 12192 39865 12220
rect 39540 12180 39546 12192
rect 39853 12189 39865 12192
rect 39899 12189 39911 12223
rect 39853 12183 39911 12189
rect 39942 12180 39948 12232
rect 40000 12180 40006 12232
rect 40236 12229 40264 12328
rect 41322 12288 41328 12300
rect 41064 12260 41328 12288
rect 40221 12223 40279 12229
rect 40221 12189 40233 12223
rect 40267 12189 40279 12223
rect 40221 12183 40279 12189
rect 40310 12180 40316 12232
rect 40368 12229 40374 12232
rect 40368 12220 40376 12229
rect 40368 12192 40413 12220
rect 40368 12183 40376 12192
rect 40368 12180 40374 12183
rect 40586 12180 40592 12232
rect 40644 12180 40650 12232
rect 40862 12180 40868 12232
rect 40920 12180 40926 12232
rect 40954 12180 40960 12232
rect 41012 12180 41018 12232
rect 37384 12124 39528 12152
rect 35437 12087 35495 12093
rect 35437 12084 35449 12087
rect 35400 12056 35449 12084
rect 35400 12044 35406 12056
rect 35437 12053 35449 12056
rect 35483 12053 35495 12087
rect 35437 12047 35495 12053
rect 35529 12087 35587 12093
rect 35529 12053 35541 12087
rect 35575 12053 35587 12087
rect 35529 12047 35587 12053
rect 35986 12044 35992 12096
rect 36044 12044 36050 12096
rect 36446 12044 36452 12096
rect 36504 12084 36510 12096
rect 37734 12084 37740 12096
rect 36504 12056 37740 12084
rect 36504 12044 36510 12056
rect 37734 12044 37740 12056
rect 37792 12084 37798 12096
rect 38654 12084 38660 12096
rect 37792 12056 38660 12084
rect 37792 12044 37798 12056
rect 38654 12044 38660 12056
rect 38712 12044 38718 12096
rect 38838 12044 38844 12096
rect 38896 12044 38902 12096
rect 39117 12087 39175 12093
rect 39117 12053 39129 12087
rect 39163 12084 39175 12087
rect 39390 12084 39396 12096
rect 39163 12056 39396 12084
rect 39163 12053 39175 12056
rect 39117 12047 39175 12053
rect 39390 12044 39396 12056
rect 39448 12044 39454 12096
rect 39500 12084 39528 12124
rect 39666 12112 39672 12164
rect 39724 12152 39730 12164
rect 40129 12155 40187 12161
rect 40129 12152 40141 12155
rect 39724 12124 40141 12152
rect 39724 12112 39730 12124
rect 40129 12121 40141 12124
rect 40175 12121 40187 12155
rect 40129 12115 40187 12121
rect 40770 12112 40776 12164
rect 40828 12112 40834 12164
rect 40497 12087 40555 12093
rect 40497 12084 40509 12087
rect 39500 12056 40509 12084
rect 40497 12053 40509 12056
rect 40543 12053 40555 12087
rect 40497 12047 40555 12053
rect 40678 12044 40684 12096
rect 40736 12084 40742 12096
rect 41064 12084 41092 12260
rect 41322 12248 41328 12260
rect 41380 12288 41386 12300
rect 41693 12291 41751 12297
rect 41693 12288 41705 12291
rect 41380 12260 41705 12288
rect 41380 12248 41386 12260
rect 41693 12257 41705 12260
rect 41739 12257 41751 12291
rect 41800 12288 41828 12328
rect 45922 12288 45928 12300
rect 41800 12260 45928 12288
rect 41693 12251 41751 12257
rect 45922 12248 45928 12260
rect 45980 12248 45986 12300
rect 46198 12180 46204 12232
rect 46256 12220 46262 12232
rect 46753 12223 46811 12229
rect 46753 12220 46765 12223
rect 46256 12192 46765 12220
rect 46256 12180 46262 12192
rect 46753 12189 46765 12192
rect 46799 12189 46811 12223
rect 46753 12183 46811 12189
rect 41969 12155 42027 12161
rect 41969 12121 41981 12155
rect 42015 12121 42027 12155
rect 41969 12115 42027 12121
rect 40736 12056 41092 12084
rect 41141 12087 41199 12093
rect 40736 12044 40742 12056
rect 41141 12053 41153 12087
rect 41187 12084 41199 12087
rect 41984 12084 42012 12115
rect 42426 12112 42432 12164
rect 42484 12112 42490 12164
rect 41187 12056 42012 12084
rect 41187 12053 41199 12056
rect 41141 12047 41199 12053
rect 1104 11994 58880 12016
rect 1104 11942 4874 11994
rect 4926 11942 4938 11994
rect 4990 11942 5002 11994
rect 5054 11942 5066 11994
rect 5118 11942 5130 11994
rect 5182 11942 35594 11994
rect 35646 11942 35658 11994
rect 35710 11942 35722 11994
rect 35774 11942 35786 11994
rect 35838 11942 35850 11994
rect 35902 11942 58880 11994
rect 1104 11920 58880 11942
rect 17494 11840 17500 11892
rect 17552 11880 17558 11892
rect 19242 11880 19248 11892
rect 17552 11852 19248 11880
rect 17552 11840 17558 11852
rect 19242 11840 19248 11852
rect 19300 11840 19306 11892
rect 26694 11840 26700 11892
rect 26752 11880 26758 11892
rect 27246 11880 27252 11892
rect 26752 11852 27252 11880
rect 26752 11840 26758 11852
rect 27246 11840 27252 11852
rect 27304 11840 27310 11892
rect 29546 11840 29552 11892
rect 29604 11840 29610 11892
rect 32401 11883 32459 11889
rect 29840 11852 30972 11880
rect 13446 11772 13452 11824
rect 13504 11772 13510 11824
rect 19610 11772 19616 11824
rect 19668 11812 19674 11824
rect 19705 11815 19763 11821
rect 19705 11812 19717 11815
rect 19668 11784 19717 11812
rect 19668 11772 19674 11784
rect 19705 11781 19717 11784
rect 19751 11781 19763 11815
rect 22186 11812 22192 11824
rect 20930 11784 22192 11812
rect 19705 11775 19763 11781
rect 22186 11772 22192 11784
rect 22244 11772 22250 11824
rect 29840 11821 29868 11852
rect 29825 11815 29883 11821
rect 29825 11812 29837 11815
rect 29564 11784 29837 11812
rect 29564 11756 29592 11784
rect 29825 11781 29837 11784
rect 29871 11781 29883 11815
rect 29825 11775 29883 11781
rect 29917 11815 29975 11821
rect 29917 11781 29929 11815
rect 29963 11812 29975 11815
rect 30374 11812 30380 11824
rect 29963 11784 30380 11812
rect 29963 11781 29975 11784
rect 29917 11775 29975 11781
rect 12158 11704 12164 11756
rect 12216 11704 12222 11756
rect 14734 11704 14740 11756
rect 14792 11704 14798 11756
rect 14921 11747 14979 11753
rect 14921 11713 14933 11747
rect 14967 11713 14979 11747
rect 14921 11707 14979 11713
rect 12434 11636 12440 11688
rect 12492 11636 12498 11688
rect 13909 11679 13967 11685
rect 13909 11645 13921 11679
rect 13955 11676 13967 11679
rect 14274 11676 14280 11688
rect 13955 11648 14280 11676
rect 13955 11645 13967 11648
rect 13909 11639 13967 11645
rect 14274 11636 14280 11648
rect 14332 11676 14338 11688
rect 14553 11679 14611 11685
rect 14553 11676 14565 11679
rect 14332 11648 14565 11676
rect 14332 11636 14338 11648
rect 14553 11645 14565 11648
rect 14599 11676 14611 11679
rect 14936 11676 14964 11707
rect 17310 11704 17316 11756
rect 17368 11744 17374 11756
rect 19429 11747 19487 11753
rect 19429 11744 19441 11747
rect 17368 11716 19441 11744
rect 17368 11704 17374 11716
rect 19429 11713 19441 11716
rect 19475 11713 19487 11747
rect 19429 11707 19487 11713
rect 26694 11704 26700 11756
rect 26752 11744 26758 11756
rect 26973 11747 27031 11753
rect 26973 11744 26985 11747
rect 26752 11716 26985 11744
rect 26752 11704 26758 11716
rect 26973 11713 26985 11716
rect 27019 11713 27031 11747
rect 26973 11707 27031 11713
rect 27341 11747 27399 11753
rect 27341 11713 27353 11747
rect 27387 11744 27399 11747
rect 28350 11744 28356 11756
rect 27387 11716 28356 11744
rect 27387 11713 27399 11716
rect 27341 11707 27399 11713
rect 14599 11648 14964 11676
rect 14599 11645 14611 11648
rect 14553 11639 14611 11645
rect 21082 11636 21088 11688
rect 21140 11676 21146 11688
rect 21177 11679 21235 11685
rect 21177 11676 21189 11679
rect 21140 11648 21189 11676
rect 21140 11636 21146 11648
rect 21177 11645 21189 11648
rect 21223 11645 21235 11679
rect 21177 11639 21235 11645
rect 22462 11636 22468 11688
rect 22520 11676 22526 11688
rect 22833 11679 22891 11685
rect 22833 11676 22845 11679
rect 22520 11648 22845 11676
rect 22520 11636 22526 11648
rect 22833 11645 22845 11648
rect 22879 11645 22891 11679
rect 22833 11639 22891 11645
rect 27157 11611 27215 11617
rect 27157 11577 27169 11611
rect 27203 11608 27215 11611
rect 27356 11608 27384 11707
rect 28350 11704 28356 11716
rect 28408 11704 28414 11756
rect 28810 11704 28816 11756
rect 28868 11704 28874 11756
rect 29365 11747 29423 11753
rect 29365 11713 29377 11747
rect 29411 11713 29423 11747
rect 29365 11707 29423 11713
rect 29089 11679 29147 11685
rect 29089 11645 29101 11679
rect 29135 11645 29147 11679
rect 29089 11639 29147 11645
rect 29181 11679 29239 11685
rect 29181 11645 29193 11679
rect 29227 11676 29239 11679
rect 29270 11676 29276 11688
rect 29227 11648 29276 11676
rect 29227 11645 29239 11648
rect 29181 11639 29239 11645
rect 27203 11580 27384 11608
rect 29104 11608 29132 11639
rect 29270 11636 29276 11648
rect 29328 11636 29334 11688
rect 29380 11676 29408 11707
rect 29546 11704 29552 11756
rect 29604 11704 29610 11756
rect 29730 11753 29736 11756
rect 29728 11707 29736 11753
rect 29730 11704 29736 11707
rect 29788 11704 29794 11756
rect 29932 11676 29960 11775
rect 30374 11772 30380 11784
rect 30432 11772 30438 11824
rect 30100 11747 30158 11753
rect 30100 11713 30112 11747
rect 30146 11713 30158 11747
rect 30100 11707 30158 11713
rect 29380 11648 29960 11676
rect 29638 11608 29644 11620
rect 29104 11580 29644 11608
rect 27203 11577 27215 11580
rect 27157 11571 27215 11577
rect 29638 11568 29644 11580
rect 29696 11568 29702 11620
rect 30116 11608 30144 11707
rect 30190 11704 30196 11756
rect 30248 11704 30254 11756
rect 30944 11753 30972 11852
rect 32401 11849 32413 11883
rect 32447 11880 32459 11883
rect 32490 11880 32496 11892
rect 32447 11852 32496 11880
rect 32447 11849 32459 11852
rect 32401 11843 32459 11849
rect 31018 11772 31024 11824
rect 31076 11772 31082 11824
rect 31110 11772 31116 11824
rect 31168 11821 31174 11824
rect 31168 11815 31197 11821
rect 31185 11781 31197 11815
rect 32416 11812 32444 11843
rect 32490 11840 32496 11852
rect 32548 11840 32554 11892
rect 33226 11840 33232 11892
rect 33284 11840 33290 11892
rect 33318 11840 33324 11892
rect 33376 11840 33382 11892
rect 34882 11840 34888 11892
rect 34940 11880 34946 11892
rect 34977 11883 35035 11889
rect 34977 11880 34989 11883
rect 34940 11852 34989 11880
rect 34940 11840 34946 11852
rect 34977 11849 34989 11852
rect 35023 11849 35035 11883
rect 34977 11843 35035 11849
rect 35066 11840 35072 11892
rect 35124 11880 35130 11892
rect 35161 11883 35219 11889
rect 35161 11880 35173 11883
rect 35124 11852 35173 11880
rect 35124 11840 35130 11852
rect 35161 11849 35173 11852
rect 35207 11849 35219 11883
rect 35161 11843 35219 11849
rect 35250 11840 35256 11892
rect 35308 11880 35314 11892
rect 36633 11883 36691 11889
rect 36633 11880 36645 11883
rect 35308 11852 36645 11880
rect 35308 11840 35314 11852
rect 36633 11849 36645 11852
rect 36679 11849 36691 11883
rect 36633 11843 36691 11849
rect 37550 11840 37556 11892
rect 37608 11880 37614 11892
rect 37645 11883 37703 11889
rect 37645 11880 37657 11883
rect 37608 11852 37657 11880
rect 37608 11840 37614 11852
rect 37645 11849 37657 11852
rect 37691 11849 37703 11883
rect 37645 11843 37703 11849
rect 38378 11840 38384 11892
rect 38436 11880 38442 11892
rect 38473 11883 38531 11889
rect 38473 11880 38485 11883
rect 38436 11852 38485 11880
rect 38436 11840 38442 11852
rect 38473 11849 38485 11852
rect 38519 11849 38531 11883
rect 38473 11843 38531 11849
rect 39390 11840 39396 11892
rect 39448 11840 39454 11892
rect 39761 11883 39819 11889
rect 39761 11849 39773 11883
rect 39807 11880 39819 11883
rect 40770 11880 40776 11892
rect 39807 11852 40776 11880
rect 39807 11849 39819 11852
rect 39761 11843 39819 11849
rect 40770 11840 40776 11852
rect 40828 11840 40834 11892
rect 42426 11840 42432 11892
rect 42484 11880 42490 11892
rect 42484 11852 42932 11880
rect 42484 11840 42490 11852
rect 31168 11775 31197 11781
rect 32140 11784 32444 11812
rect 32953 11815 33011 11821
rect 31168 11772 31174 11775
rect 30837 11747 30895 11753
rect 30837 11713 30849 11747
rect 30883 11713 30895 11747
rect 30837 11707 30895 11713
rect 30929 11747 30987 11753
rect 30929 11713 30941 11747
rect 30975 11713 30987 11747
rect 32140 11744 32168 11784
rect 32953 11781 32965 11815
rect 32999 11812 33011 11815
rect 33689 11815 33747 11821
rect 33689 11812 33701 11815
rect 32999 11784 33701 11812
rect 32999 11781 33011 11784
rect 32953 11775 33011 11781
rect 33689 11781 33701 11784
rect 33735 11812 33747 11815
rect 35986 11812 35992 11824
rect 33735 11784 35992 11812
rect 33735 11781 33747 11784
rect 33689 11775 33747 11781
rect 35986 11772 35992 11784
rect 36044 11772 36050 11824
rect 36078 11772 36084 11824
rect 36136 11812 36142 11824
rect 36357 11815 36415 11821
rect 36357 11812 36369 11815
rect 36136 11784 36369 11812
rect 36136 11772 36142 11784
rect 36357 11781 36369 11784
rect 36403 11781 36415 11815
rect 36357 11775 36415 11781
rect 37844 11784 38424 11812
rect 30929 11707 30987 11713
rect 31220 11716 32168 11744
rect 32217 11747 32275 11753
rect 30742 11636 30748 11688
rect 30800 11676 30806 11688
rect 30852 11676 30880 11707
rect 31220 11676 31248 11716
rect 32217 11713 32229 11747
rect 32263 11744 32275 11747
rect 32306 11744 32312 11756
rect 32263 11716 32312 11744
rect 32263 11713 32275 11716
rect 32217 11707 32275 11713
rect 32306 11704 32312 11716
rect 32364 11704 32370 11756
rect 32493 11747 32551 11753
rect 32493 11713 32505 11747
rect 32539 11713 32551 11747
rect 32493 11707 32551 11713
rect 30800 11648 31248 11676
rect 31297 11679 31355 11685
rect 30800 11636 30806 11648
rect 31297 11645 31309 11679
rect 31343 11676 31355 11679
rect 32508 11676 32536 11707
rect 32582 11704 32588 11756
rect 32640 11704 32646 11756
rect 32766 11753 32772 11756
rect 32733 11747 32772 11753
rect 32733 11713 32745 11747
rect 32733 11707 32772 11713
rect 32766 11704 32772 11707
rect 32824 11704 32830 11756
rect 32858 11704 32864 11756
rect 32916 11704 32922 11756
rect 33042 11704 33048 11756
rect 33100 11753 33106 11756
rect 33100 11744 33108 11753
rect 33100 11716 33145 11744
rect 33100 11707 33108 11716
rect 33100 11704 33106 11707
rect 33318 11704 33324 11756
rect 33376 11704 33382 11756
rect 33505 11747 33563 11753
rect 33505 11713 33517 11747
rect 33551 11713 33563 11747
rect 33505 11707 33563 11713
rect 33520 11676 33548 11707
rect 33594 11704 33600 11756
rect 33652 11704 33658 11756
rect 33778 11704 33784 11756
rect 33836 11704 33842 11756
rect 34606 11704 34612 11756
rect 34664 11744 34670 11756
rect 35102 11747 35160 11753
rect 35102 11744 35114 11747
rect 34664 11742 34928 11744
rect 34992 11742 35114 11744
rect 34664 11716 35114 11742
rect 34664 11704 34670 11716
rect 34900 11714 35020 11716
rect 35102 11713 35114 11716
rect 35148 11713 35160 11747
rect 35102 11707 35160 11713
rect 35250 11704 35256 11756
rect 35308 11744 35314 11756
rect 35805 11747 35863 11753
rect 35805 11744 35817 11747
rect 35308 11716 35817 11744
rect 35308 11704 35314 11716
rect 35805 11713 35817 11716
rect 35851 11713 35863 11747
rect 35805 11707 35863 11713
rect 31343 11648 32444 11676
rect 32508 11648 33548 11676
rect 31343 11645 31355 11648
rect 31297 11639 31355 11645
rect 31312 11608 31340 11639
rect 30116 11580 31340 11608
rect 31478 11568 31484 11620
rect 31536 11608 31542 11620
rect 32217 11611 32275 11617
rect 32217 11608 32229 11611
rect 31536 11580 32229 11608
rect 31536 11568 31542 11580
rect 32217 11577 32229 11580
rect 32263 11577 32275 11611
rect 32416 11608 32444 11648
rect 32674 11608 32680 11620
rect 32416 11580 32680 11608
rect 32217 11571 32275 11577
rect 32674 11568 32680 11580
rect 32732 11568 32738 11620
rect 33520 11608 33548 11648
rect 35342 11636 35348 11688
rect 35400 11676 35406 11688
rect 35621 11679 35679 11685
rect 35621 11676 35633 11679
rect 35400 11648 35633 11676
rect 35400 11636 35406 11648
rect 35621 11645 35633 11648
rect 35667 11676 35679 11679
rect 36096 11676 36124 11772
rect 36262 11704 36268 11756
rect 36320 11704 36326 11756
rect 36449 11747 36507 11753
rect 36449 11713 36461 11747
rect 36495 11744 36507 11747
rect 36538 11744 36544 11756
rect 36495 11716 36544 11744
rect 36495 11713 36507 11716
rect 36449 11707 36507 11713
rect 36538 11704 36544 11716
rect 36596 11704 36602 11756
rect 36630 11704 36636 11756
rect 36688 11744 36694 11756
rect 36725 11747 36783 11753
rect 36725 11744 36737 11747
rect 36688 11716 36737 11744
rect 36688 11704 36694 11716
rect 36725 11713 36737 11716
rect 36771 11713 36783 11747
rect 36725 11707 36783 11713
rect 37734 11704 37740 11756
rect 37792 11744 37798 11756
rect 37844 11753 37872 11784
rect 37829 11747 37887 11753
rect 37829 11744 37841 11747
rect 37792 11716 37841 11744
rect 37792 11704 37798 11716
rect 37829 11713 37841 11716
rect 37875 11713 37887 11747
rect 37829 11707 37887 11713
rect 37918 11704 37924 11756
rect 37976 11744 37982 11756
rect 38105 11747 38163 11753
rect 38105 11744 38117 11747
rect 37976 11716 38117 11744
rect 37976 11704 37982 11716
rect 38105 11713 38117 11716
rect 38151 11713 38163 11747
rect 38105 11707 38163 11713
rect 38286 11704 38292 11756
rect 38344 11704 38350 11756
rect 38396 11753 38424 11784
rect 40034 11772 40040 11824
rect 40092 11812 40098 11824
rect 40129 11815 40187 11821
rect 40129 11812 40141 11815
rect 40092 11784 40141 11812
rect 40092 11772 40098 11784
rect 40129 11781 40141 11784
rect 40175 11812 40187 11815
rect 40954 11812 40960 11824
rect 40175 11784 40960 11812
rect 40175 11781 40187 11784
rect 40129 11775 40187 11781
rect 40954 11772 40960 11784
rect 41012 11772 41018 11824
rect 42794 11772 42800 11824
rect 42852 11772 42858 11824
rect 42904 11812 42932 11852
rect 44266 11840 44272 11892
rect 44324 11840 44330 11892
rect 42904 11784 43286 11812
rect 38381 11747 38439 11753
rect 38381 11713 38393 11747
rect 38427 11713 38439 11747
rect 38381 11707 38439 11713
rect 38470 11704 38476 11756
rect 38528 11742 38534 11756
rect 38565 11745 38623 11751
rect 38565 11742 38577 11745
rect 38528 11714 38577 11742
rect 38528 11704 38534 11714
rect 38565 11711 38577 11714
rect 38611 11711 38623 11745
rect 38565 11705 38623 11711
rect 38746 11704 38752 11756
rect 38804 11734 38810 11756
rect 38841 11747 38899 11753
rect 38841 11734 38853 11747
rect 38804 11713 38853 11734
rect 38887 11713 38899 11747
rect 38804 11707 38899 11713
rect 38804 11706 38884 11707
rect 38804 11704 38810 11706
rect 38930 11704 38936 11756
rect 38988 11704 38994 11756
rect 39301 11747 39359 11753
rect 39301 11713 39313 11747
rect 39347 11713 39359 11747
rect 39301 11707 39359 11713
rect 39577 11747 39635 11753
rect 39577 11713 39589 11747
rect 39623 11744 39635 11747
rect 39623 11716 39804 11744
rect 39623 11713 39635 11716
rect 39577 11707 39635 11713
rect 35667 11648 36124 11676
rect 36173 11679 36231 11685
rect 35667 11645 35679 11648
rect 35621 11639 35679 11645
rect 36173 11645 36185 11679
rect 36219 11676 36231 11679
rect 38013 11679 38071 11685
rect 38013 11676 38025 11679
rect 36219 11648 38025 11676
rect 36219 11645 36231 11648
rect 36173 11639 36231 11645
rect 38013 11645 38025 11648
rect 38059 11645 38071 11679
rect 38013 11639 38071 11645
rect 38657 11679 38715 11685
rect 38657 11645 38669 11679
rect 38703 11645 38715 11679
rect 38657 11639 38715 11645
rect 35529 11611 35587 11617
rect 35529 11608 35541 11611
rect 33520 11580 35541 11608
rect 35529 11577 35541 11580
rect 35575 11577 35587 11611
rect 35529 11571 35587 11577
rect 13998 11500 14004 11552
rect 14056 11500 14062 11552
rect 15105 11543 15163 11549
rect 15105 11509 15117 11543
rect 15151 11540 15163 11543
rect 15470 11540 15476 11552
rect 15151 11512 15476 11540
rect 15151 11509 15163 11512
rect 15105 11503 15163 11509
rect 15470 11500 15476 11512
rect 15528 11500 15534 11552
rect 16390 11500 16396 11552
rect 16448 11540 16454 11552
rect 20162 11540 20168 11552
rect 16448 11512 20168 11540
rect 16448 11500 16454 11512
rect 20162 11500 20168 11512
rect 20220 11500 20226 11552
rect 22002 11500 22008 11552
rect 22060 11540 22066 11552
rect 22281 11543 22339 11549
rect 22281 11540 22293 11543
rect 22060 11512 22293 11540
rect 22060 11500 22066 11512
rect 22281 11509 22293 11512
rect 22327 11509 22339 11543
rect 22281 11503 22339 11509
rect 27433 11543 27491 11549
rect 27433 11509 27445 11543
rect 27479 11540 27491 11543
rect 27614 11540 27620 11552
rect 27479 11512 27620 11540
rect 27479 11509 27491 11512
rect 27433 11503 27491 11509
rect 27614 11500 27620 11512
rect 27672 11500 27678 11552
rect 27982 11500 27988 11552
rect 28040 11540 28046 11552
rect 28718 11540 28724 11552
rect 28040 11512 28724 11540
rect 28040 11500 28046 11512
rect 28718 11500 28724 11512
rect 28776 11540 28782 11552
rect 28997 11543 29055 11549
rect 28997 11540 29009 11543
rect 28776 11512 29009 11540
rect 28776 11500 28782 11512
rect 28997 11509 29009 11512
rect 29043 11509 29055 11543
rect 28997 11503 29055 11509
rect 29178 11500 29184 11552
rect 29236 11500 29242 11552
rect 30466 11500 30472 11552
rect 30524 11540 30530 11552
rect 30653 11543 30711 11549
rect 30653 11540 30665 11543
rect 30524 11512 30665 11540
rect 30524 11500 30530 11512
rect 30653 11509 30665 11512
rect 30699 11509 30711 11543
rect 30653 11503 30711 11509
rect 30926 11500 30932 11552
rect 30984 11540 30990 11552
rect 33410 11540 33416 11552
rect 30984 11512 33416 11540
rect 30984 11500 30990 11512
rect 33410 11500 33416 11512
rect 33468 11500 33474 11552
rect 34330 11500 34336 11552
rect 34388 11540 34394 11552
rect 35342 11540 35348 11552
rect 34388 11512 35348 11540
rect 34388 11500 34394 11512
rect 35342 11500 35348 11512
rect 35400 11500 35406 11552
rect 35544 11540 35572 11571
rect 36262 11568 36268 11620
rect 36320 11608 36326 11620
rect 37921 11611 37979 11617
rect 37921 11608 37933 11611
rect 36320 11580 37933 11608
rect 36320 11568 36326 11580
rect 37921 11577 37933 11580
rect 37967 11577 37979 11611
rect 38672 11608 38700 11639
rect 39022 11636 39028 11688
rect 39080 11636 39086 11688
rect 39114 11636 39120 11688
rect 39172 11636 39178 11688
rect 39316 11676 39344 11707
rect 39666 11676 39672 11688
rect 39316 11648 39672 11676
rect 39666 11636 39672 11648
rect 39724 11636 39730 11688
rect 39776 11608 39804 11716
rect 39850 11704 39856 11756
rect 39908 11704 39914 11756
rect 39942 11704 39948 11756
rect 40000 11704 40006 11756
rect 41322 11704 41328 11756
rect 41380 11744 41386 11756
rect 42521 11747 42579 11753
rect 42521 11744 42533 11747
rect 41380 11716 42533 11744
rect 41380 11704 41386 11716
rect 42521 11713 42533 11716
rect 42567 11713 42579 11747
rect 42521 11707 42579 11713
rect 38672 11580 39804 11608
rect 40129 11611 40187 11617
rect 37921 11571 37979 11577
rect 40129 11577 40141 11611
rect 40175 11608 40187 11611
rect 40586 11608 40592 11620
rect 40175 11580 40592 11608
rect 40175 11577 40187 11580
rect 40129 11571 40187 11577
rect 36630 11540 36636 11552
rect 35544 11512 36636 11540
rect 36630 11500 36636 11512
rect 36688 11540 36694 11552
rect 37826 11540 37832 11552
rect 36688 11512 37832 11540
rect 36688 11500 36694 11512
rect 37826 11500 37832 11512
rect 37884 11500 37890 11552
rect 37936 11540 37964 11571
rect 40586 11568 40592 11580
rect 40644 11568 40650 11620
rect 39022 11540 39028 11552
rect 37936 11512 39028 11540
rect 39022 11500 39028 11512
rect 39080 11540 39086 11552
rect 39206 11540 39212 11552
rect 39080 11512 39212 11540
rect 39080 11500 39086 11512
rect 39206 11500 39212 11512
rect 39264 11500 39270 11552
rect 1104 11450 58880 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 58880 11450
rect 1104 11376 58880 11398
rect 12253 11339 12311 11345
rect 12253 11305 12265 11339
rect 12299 11336 12311 11339
rect 12434 11336 12440 11348
rect 12299 11308 12440 11336
rect 12299 11305 12311 11308
rect 12253 11299 12311 11305
rect 12434 11296 12440 11308
rect 12492 11296 12498 11348
rect 14826 11296 14832 11348
rect 14884 11296 14890 11348
rect 15013 11339 15071 11345
rect 15013 11305 15025 11339
rect 15059 11336 15071 11339
rect 15654 11336 15660 11348
rect 15059 11308 15660 11336
rect 15059 11305 15071 11308
rect 15013 11299 15071 11305
rect 15654 11296 15660 11308
rect 15712 11296 15718 11348
rect 16390 11296 16396 11348
rect 16448 11296 16454 11348
rect 16666 11296 16672 11348
rect 16724 11336 16730 11348
rect 16761 11339 16819 11345
rect 16761 11336 16773 11339
rect 16724 11308 16773 11336
rect 16724 11296 16730 11308
rect 16761 11305 16773 11308
rect 16807 11305 16819 11339
rect 16761 11299 16819 11305
rect 22462 11296 22468 11348
rect 22520 11296 22526 11348
rect 27985 11339 28043 11345
rect 27985 11305 27997 11339
rect 28031 11336 28043 11339
rect 28031 11308 28856 11336
rect 28031 11305 28043 11308
rect 27985 11299 28043 11305
rect 14093 11271 14151 11277
rect 14093 11237 14105 11271
rect 14139 11268 14151 11271
rect 14844 11268 14872 11296
rect 14139 11240 14872 11268
rect 15197 11271 15255 11277
rect 14139 11237 14151 11240
rect 14093 11231 14151 11237
rect 15197 11237 15209 11271
rect 15243 11237 15255 11271
rect 15197 11231 15255 11237
rect 12713 11203 12771 11209
rect 12713 11169 12725 11203
rect 12759 11200 12771 11203
rect 13538 11200 13544 11212
rect 12759 11172 13544 11200
rect 12759 11169 12771 11172
rect 12713 11163 12771 11169
rect 13538 11160 13544 11172
rect 13596 11200 13602 11212
rect 13596 11172 14412 11200
rect 13596 11160 13602 11172
rect 12621 11135 12679 11141
rect 12621 11101 12633 11135
rect 12667 11132 12679 11135
rect 13998 11132 14004 11144
rect 12667 11104 14004 11132
rect 12667 11101 12679 11104
rect 12621 11095 12679 11101
rect 13998 11092 14004 11104
rect 14056 11092 14062 11144
rect 14090 11092 14096 11144
rect 14148 11092 14154 11144
rect 14274 11092 14280 11144
rect 14332 11092 14338 11144
rect 14384 11141 14412 11172
rect 14734 11160 14740 11212
rect 14792 11200 14798 11212
rect 14829 11203 14887 11209
rect 14829 11200 14841 11203
rect 14792 11172 14841 11200
rect 14792 11160 14798 11172
rect 14829 11169 14841 11172
rect 14875 11169 14887 11203
rect 15212 11200 15240 11231
rect 15286 11228 15292 11280
rect 15344 11228 15350 11280
rect 16577 11271 16635 11277
rect 16577 11237 16589 11271
rect 16623 11268 16635 11271
rect 17218 11268 17224 11280
rect 16623 11240 17224 11268
rect 16623 11237 16635 11240
rect 16577 11231 16635 11237
rect 17218 11228 17224 11240
rect 17276 11228 17282 11280
rect 18230 11228 18236 11280
rect 18288 11268 18294 11280
rect 18785 11271 18843 11277
rect 18785 11268 18797 11271
rect 18288 11240 18797 11268
rect 18288 11228 18294 11240
rect 18785 11237 18797 11240
rect 18831 11237 18843 11271
rect 22554 11268 22560 11280
rect 18785 11231 18843 11237
rect 18892 11240 22560 11268
rect 16301 11203 16359 11209
rect 15212 11172 16252 11200
rect 14829 11163 14887 11169
rect 14369 11135 14427 11141
rect 14369 11101 14381 11135
rect 14415 11101 14427 11135
rect 14369 11095 14427 11101
rect 15013 11135 15071 11141
rect 15013 11101 15025 11135
rect 15059 11101 15071 11135
rect 15013 11095 15071 11101
rect 14292 11064 14320 11092
rect 14737 11067 14795 11073
rect 14737 11064 14749 11067
rect 14292 11036 14749 11064
rect 14737 11033 14749 11036
rect 14783 11033 14795 11067
rect 15028 11064 15056 11095
rect 15470 11092 15476 11144
rect 15528 11132 15534 11144
rect 15528 11104 15976 11132
rect 15528 11092 15534 11104
rect 15838 11064 15844 11076
rect 15028 11036 15844 11064
rect 14737 11027 14795 11033
rect 15838 11024 15844 11036
rect 15896 11024 15902 11076
rect 15948 11064 15976 11104
rect 16022 11092 16028 11144
rect 16080 11132 16086 11144
rect 16117 11135 16175 11141
rect 16117 11132 16129 11135
rect 16080 11104 16129 11132
rect 16080 11092 16086 11104
rect 16117 11101 16129 11104
rect 16163 11101 16175 11135
rect 16224 11132 16252 11172
rect 16301 11169 16313 11203
rect 16347 11200 16359 11203
rect 17862 11200 17868 11212
rect 16347 11172 17868 11200
rect 16347 11169 16359 11172
rect 16301 11163 16359 11169
rect 17862 11160 17868 11172
rect 17920 11160 17926 11212
rect 16393 11135 16451 11141
rect 16393 11132 16405 11135
rect 16224 11104 16405 11132
rect 16117 11095 16175 11101
rect 16393 11101 16405 11104
rect 16439 11101 16451 11135
rect 16393 11095 16451 11101
rect 16942 11092 16948 11144
rect 17000 11092 17006 11144
rect 17310 11092 17316 11144
rect 17368 11132 17374 11144
rect 18509 11135 18567 11141
rect 18509 11132 18521 11135
rect 17368 11104 18521 11132
rect 17368 11092 17374 11104
rect 18509 11101 18521 11104
rect 18555 11132 18567 11135
rect 18892 11132 18920 11240
rect 22554 11228 22560 11240
rect 22612 11228 22618 11280
rect 28534 11228 28540 11280
rect 28592 11228 28598 11280
rect 28828 11268 28856 11308
rect 28902 11296 28908 11348
rect 28960 11336 28966 11348
rect 29822 11336 29828 11348
rect 28960 11308 29828 11336
rect 28960 11296 28966 11308
rect 29822 11296 29828 11308
rect 29880 11296 29886 11348
rect 30285 11339 30343 11345
rect 30285 11305 30297 11339
rect 30331 11336 30343 11339
rect 30558 11336 30564 11348
rect 30331 11308 30564 11336
rect 30331 11305 30343 11308
rect 30285 11299 30343 11305
rect 30558 11296 30564 11308
rect 30616 11296 30622 11348
rect 33318 11296 33324 11348
rect 33376 11336 33382 11348
rect 36446 11336 36452 11348
rect 33376 11308 36452 11336
rect 33376 11296 33382 11308
rect 36446 11296 36452 11308
rect 36504 11296 36510 11348
rect 37918 11296 37924 11348
rect 37976 11336 37982 11348
rect 38381 11339 38439 11345
rect 38381 11336 38393 11339
rect 37976 11308 38393 11336
rect 37976 11296 37982 11308
rect 38381 11305 38393 11308
rect 38427 11305 38439 11339
rect 38381 11299 38439 11305
rect 38654 11296 38660 11348
rect 38712 11336 38718 11348
rect 38749 11339 38807 11345
rect 38749 11336 38761 11339
rect 38712 11308 38761 11336
rect 38712 11296 38718 11308
rect 38749 11305 38761 11308
rect 38795 11305 38807 11339
rect 38749 11299 38807 11305
rect 39114 11296 39120 11348
rect 39172 11296 39178 11348
rect 39206 11296 39212 11348
rect 39264 11336 39270 11348
rect 39301 11339 39359 11345
rect 39301 11336 39313 11339
rect 39264 11308 39313 11336
rect 39264 11296 39270 11308
rect 39301 11305 39313 11308
rect 39347 11305 39359 11339
rect 39850 11336 39856 11348
rect 39301 11299 39359 11305
rect 39408 11308 39856 11336
rect 29914 11268 29920 11280
rect 28828 11240 29920 11268
rect 29914 11228 29920 11240
rect 29972 11228 29978 11280
rect 30374 11228 30380 11280
rect 30432 11268 30438 11280
rect 32493 11271 32551 11277
rect 32493 11268 32505 11271
rect 30432 11240 32505 11268
rect 30432 11228 30438 11240
rect 32493 11237 32505 11240
rect 32539 11268 32551 11271
rect 32858 11268 32864 11280
rect 32539 11240 32864 11268
rect 32539 11237 32551 11240
rect 32493 11231 32551 11237
rect 32858 11228 32864 11240
rect 32916 11228 32922 11280
rect 35434 11228 35440 11280
rect 35492 11228 35498 11280
rect 37826 11228 37832 11280
rect 37884 11268 37890 11280
rect 39408 11268 39436 11308
rect 39850 11296 39856 11308
rect 39908 11296 39914 11348
rect 40497 11271 40555 11277
rect 40497 11268 40509 11271
rect 37884 11240 39436 11268
rect 39500 11240 40509 11268
rect 37884 11228 37890 11240
rect 21358 11160 21364 11212
rect 21416 11200 21422 11212
rect 21913 11203 21971 11209
rect 21913 11200 21925 11203
rect 21416 11172 21925 11200
rect 21416 11160 21422 11172
rect 21913 11169 21925 11172
rect 21959 11169 21971 11203
rect 21913 11163 21971 11169
rect 22373 11203 22431 11209
rect 22373 11169 22385 11203
rect 22419 11200 22431 11203
rect 23937 11203 23995 11209
rect 23937 11200 23949 11203
rect 22419 11172 23949 11200
rect 22419 11169 22431 11172
rect 22373 11163 22431 11169
rect 23937 11169 23949 11172
rect 23983 11169 23995 11203
rect 23937 11163 23995 11169
rect 28445 11203 28503 11209
rect 28445 11169 28457 11203
rect 28491 11200 28503 11203
rect 28552 11200 28580 11228
rect 29270 11200 29276 11212
rect 28491 11172 29276 11200
rect 28491 11169 28503 11172
rect 28445 11163 28503 11169
rect 29270 11160 29276 11172
rect 29328 11200 29334 11212
rect 29328 11172 30696 11200
rect 29328 11160 29334 11172
rect 18555 11104 18920 11132
rect 18555 11101 18567 11104
rect 18509 11095 18567 11101
rect 19886 11092 19892 11144
rect 19944 11092 19950 11144
rect 20257 11135 20315 11141
rect 20257 11132 20269 11135
rect 19996 11104 20269 11132
rect 17037 11067 17095 11073
rect 17037 11064 17049 11067
rect 15948 11036 17049 11064
rect 17037 11033 17049 11036
rect 17083 11033 17095 11067
rect 17037 11027 17095 11033
rect 18785 11067 18843 11073
rect 18785 11033 18797 11067
rect 18831 11064 18843 11067
rect 19337 11067 19395 11073
rect 19337 11064 19349 11067
rect 18831 11036 19349 11064
rect 18831 11033 18843 11036
rect 18785 11027 18843 11033
rect 19337 11033 19349 11036
rect 19383 11033 19395 11067
rect 19337 11027 19395 11033
rect 15562 10956 15568 11008
rect 15620 10956 15626 11008
rect 15654 10956 15660 11008
rect 15712 10956 15718 11008
rect 17126 10956 17132 11008
rect 17184 10956 17190 11008
rect 17954 10956 17960 11008
rect 18012 10996 18018 11008
rect 18601 10999 18659 11005
rect 18601 10996 18613 10999
rect 18012 10968 18613 10996
rect 18012 10956 18018 10968
rect 18601 10965 18613 10968
rect 18647 10996 18659 10999
rect 19242 10996 19248 11008
rect 18647 10968 19248 10996
rect 18647 10965 18659 10968
rect 18601 10959 18659 10965
rect 19242 10956 19248 10968
rect 19300 10996 19306 11008
rect 19996 10996 20024 11104
rect 20257 11101 20269 11104
rect 20303 11101 20315 11135
rect 20257 11095 20315 11101
rect 20441 11135 20499 11141
rect 20441 11101 20453 11135
rect 20487 11132 20499 11135
rect 20714 11132 20720 11144
rect 20487 11104 20720 11132
rect 20487 11101 20499 11104
rect 20441 11095 20499 11101
rect 20714 11092 20720 11104
rect 20772 11092 20778 11144
rect 22002 11092 22008 11144
rect 22060 11092 22066 11144
rect 24213 11135 24271 11141
rect 24213 11101 24225 11135
rect 24259 11132 24271 11135
rect 24946 11132 24952 11144
rect 24259 11104 24952 11132
rect 24259 11101 24271 11104
rect 24213 11095 24271 11101
rect 24946 11092 24952 11104
rect 25004 11092 25010 11144
rect 27525 11135 27583 11141
rect 27525 11101 27537 11135
rect 27571 11132 27583 11135
rect 28169 11135 28227 11141
rect 28169 11132 28181 11135
rect 27571 11104 28181 11132
rect 27571 11101 27583 11104
rect 27525 11095 27583 11101
rect 28169 11101 28181 11104
rect 28215 11101 28227 11135
rect 28169 11095 28227 11101
rect 28261 11135 28319 11141
rect 28261 11101 28273 11135
rect 28307 11101 28319 11135
rect 28261 11095 28319 11101
rect 22922 11024 22928 11076
rect 22980 11024 22986 11076
rect 27614 11024 27620 11076
rect 27672 11064 27678 11076
rect 27709 11067 27767 11073
rect 27709 11064 27721 11067
rect 27672 11036 27721 11064
rect 27672 11024 27678 11036
rect 27709 11033 27721 11036
rect 27755 11033 27767 11067
rect 27709 11027 27767 11033
rect 27890 11024 27896 11076
rect 27948 11024 27954 11076
rect 28276 11064 28304 11095
rect 28350 11092 28356 11144
rect 28408 11132 28414 11144
rect 28537 11135 28595 11141
rect 28537 11132 28549 11135
rect 28408 11104 28549 11132
rect 28408 11092 28414 11104
rect 28537 11101 28549 11104
rect 28583 11132 28595 11135
rect 28994 11132 29000 11144
rect 28583 11104 29000 11132
rect 28583 11101 28595 11104
rect 28537 11095 28595 11101
rect 28994 11092 29000 11104
rect 29052 11092 29058 11144
rect 29086 11092 29092 11144
rect 29144 11092 29150 11144
rect 30466 11092 30472 11144
rect 30524 11092 30530 11144
rect 30668 11141 30696 11172
rect 31110 11160 31116 11212
rect 31168 11200 31174 11212
rect 31168 11172 32168 11200
rect 31168 11160 31174 11172
rect 32140 11141 32168 11172
rect 32306 11160 32312 11212
rect 32364 11160 32370 11212
rect 33502 11200 33508 11212
rect 32416 11172 33508 11200
rect 30653 11135 30711 11141
rect 30653 11101 30665 11135
rect 30699 11101 30711 11135
rect 30653 11095 30711 11101
rect 30745 11135 30803 11141
rect 30745 11101 30757 11135
rect 30791 11132 30803 11135
rect 32125 11135 32183 11141
rect 30791 11104 32076 11132
rect 30791 11101 30803 11104
rect 30745 11095 30803 11101
rect 29546 11064 29552 11076
rect 28276 11036 29552 11064
rect 29546 11024 29552 11036
rect 29604 11024 29610 11076
rect 30668 11064 30696 11095
rect 32048 11064 32076 11104
rect 32125 11101 32137 11135
rect 32171 11132 32183 11135
rect 32416 11132 32444 11172
rect 33502 11160 33508 11172
rect 33560 11160 33566 11212
rect 36538 11200 36544 11212
rect 35544 11172 36544 11200
rect 32171 11104 32444 11132
rect 32171 11101 32183 11104
rect 32125 11095 32183 11101
rect 32490 11092 32496 11144
rect 32548 11132 32554 11144
rect 33318 11132 33324 11144
rect 32548 11104 33324 11132
rect 32548 11092 32554 11104
rect 33318 11092 33324 11104
rect 33376 11092 33382 11144
rect 34790 11092 34796 11144
rect 34848 11092 34854 11144
rect 34882 11092 34888 11144
rect 34940 11092 34946 11144
rect 35161 11135 35219 11141
rect 35161 11132 35173 11135
rect 34992 11104 35173 11132
rect 34330 11064 34336 11076
rect 30668 11036 31754 11064
rect 32048 11036 34336 11064
rect 19300 10968 20024 10996
rect 19300 10956 19306 10968
rect 20070 10956 20076 11008
rect 20128 10956 20134 11008
rect 31726 10996 31754 11036
rect 34330 11024 34336 11036
rect 34388 11024 34394 11076
rect 34992 11064 35020 11104
rect 35161 11101 35173 11104
rect 35207 11101 35219 11135
rect 35161 11095 35219 11101
rect 35253 11135 35311 11141
rect 35253 11101 35265 11135
rect 35299 11132 35311 11135
rect 35434 11132 35440 11144
rect 35299 11104 35440 11132
rect 35299 11101 35311 11104
rect 35253 11095 35311 11101
rect 35434 11092 35440 11104
rect 35492 11132 35498 11144
rect 35544 11132 35572 11172
rect 36538 11160 36544 11172
rect 36596 11200 36602 11212
rect 39500 11209 39528 11240
rect 40497 11237 40509 11240
rect 40543 11237 40555 11271
rect 40497 11231 40555 11237
rect 39485 11203 39543 11209
rect 36596 11172 38608 11200
rect 36596 11160 36602 11172
rect 38580 11144 38608 11172
rect 39485 11169 39497 11203
rect 39531 11169 39543 11203
rect 39485 11163 39543 11169
rect 40310 11160 40316 11212
rect 40368 11160 40374 11212
rect 35492 11104 35572 11132
rect 35492 11092 35498 11104
rect 38286 11092 38292 11144
rect 38344 11092 38350 11144
rect 38473 11135 38531 11141
rect 38473 11101 38485 11135
rect 38519 11101 38531 11135
rect 38473 11095 38531 11101
rect 34440 11036 35020 11064
rect 35069 11067 35127 11073
rect 34440 11008 34468 11036
rect 35069 11033 35081 11067
rect 35115 11064 35127 11067
rect 35342 11064 35348 11076
rect 35115 11036 35348 11064
rect 35115 11033 35127 11036
rect 35069 11027 35127 11033
rect 35342 11024 35348 11036
rect 35400 11024 35406 11076
rect 38102 11024 38108 11076
rect 38160 11064 38166 11076
rect 38488 11064 38516 11095
rect 38562 11092 38568 11144
rect 38620 11092 38626 11144
rect 39206 11092 39212 11144
rect 39264 11132 39270 11144
rect 39301 11135 39359 11141
rect 39301 11132 39313 11135
rect 39264 11104 39313 11132
rect 39264 11092 39270 11104
rect 39301 11101 39313 11104
rect 39347 11101 39359 11135
rect 39853 11135 39911 11141
rect 39853 11132 39865 11135
rect 39301 11095 39359 11101
rect 39408 11104 39865 11132
rect 39408 11064 39436 11104
rect 39853 11101 39865 11104
rect 39899 11101 39911 11135
rect 39853 11095 39911 11101
rect 40221 11135 40279 11141
rect 40221 11101 40233 11135
rect 40267 11132 40279 11135
rect 40267 11104 41414 11132
rect 40267 11101 40279 11104
rect 40221 11095 40279 11101
rect 38160 11036 39436 11064
rect 38160 11024 38166 11036
rect 39574 11024 39580 11076
rect 39632 11024 39638 11076
rect 41386 11064 41414 11104
rect 41690 11064 41696 11076
rect 41386 11036 41696 11064
rect 41690 11024 41696 11036
rect 41748 11024 41754 11076
rect 34422 10996 34428 11008
rect 31726 10968 34428 10996
rect 34422 10956 34428 10968
rect 34480 10956 34486 11008
rect 34514 10956 34520 11008
rect 34572 10996 34578 11008
rect 37366 10996 37372 11008
rect 34572 10968 37372 10996
rect 34572 10956 34578 10968
rect 37366 10956 37372 10968
rect 37424 10996 37430 11008
rect 39206 10996 39212 11008
rect 37424 10968 39212 10996
rect 37424 10956 37430 10968
rect 39206 10956 39212 10968
rect 39264 10996 39270 11008
rect 39482 10996 39488 11008
rect 39264 10968 39488 10996
rect 39264 10956 39270 10968
rect 39482 10956 39488 10968
rect 39540 10956 39546 11008
rect 1104 10906 58880 10928
rect 1104 10854 4874 10906
rect 4926 10854 4938 10906
rect 4990 10854 5002 10906
rect 5054 10854 5066 10906
rect 5118 10854 5130 10906
rect 5182 10854 35594 10906
rect 35646 10854 35658 10906
rect 35710 10854 35722 10906
rect 35774 10854 35786 10906
rect 35838 10854 35850 10906
rect 35902 10854 58880 10906
rect 1104 10832 58880 10854
rect 13538 10752 13544 10804
rect 13596 10752 13602 10804
rect 16669 10795 16727 10801
rect 16669 10761 16681 10795
rect 16715 10792 16727 10795
rect 17126 10792 17132 10804
rect 16715 10764 17132 10792
rect 16715 10761 16727 10764
rect 16669 10755 16727 10761
rect 17126 10752 17132 10764
rect 17184 10752 17190 10804
rect 20162 10752 20168 10804
rect 20220 10752 20226 10804
rect 22462 10792 22468 10804
rect 22066 10764 22468 10792
rect 22066 10736 22094 10764
rect 22462 10752 22468 10764
rect 22520 10752 22526 10804
rect 26694 10752 26700 10804
rect 26752 10752 26758 10804
rect 27157 10795 27215 10801
rect 27157 10761 27169 10795
rect 27203 10761 27215 10795
rect 27157 10755 27215 10761
rect 13693 10727 13751 10733
rect 13693 10724 13705 10727
rect 13004 10696 13705 10724
rect 13004 10588 13032 10696
rect 13693 10693 13705 10696
rect 13739 10693 13751 10727
rect 13693 10687 13751 10693
rect 13906 10684 13912 10736
rect 13964 10724 13970 10736
rect 15838 10724 15844 10736
rect 13964 10696 15844 10724
rect 13964 10684 13970 10696
rect 15838 10684 15844 10696
rect 15896 10724 15902 10736
rect 16945 10727 17003 10733
rect 16945 10724 16957 10727
rect 15896 10696 16957 10724
rect 15896 10684 15902 10696
rect 16945 10693 16957 10696
rect 16991 10693 17003 10727
rect 17954 10724 17960 10736
rect 16945 10687 17003 10693
rect 17052 10696 17960 10724
rect 13081 10659 13139 10665
rect 13081 10625 13093 10659
rect 13127 10656 13139 10659
rect 14001 10659 14059 10665
rect 14001 10656 14013 10659
rect 13127 10628 14013 10656
rect 13127 10625 13139 10628
rect 13081 10619 13139 10625
rect 14001 10625 14013 10628
rect 14047 10625 14059 10659
rect 14001 10619 14059 10625
rect 14645 10659 14703 10665
rect 14645 10625 14657 10659
rect 14691 10656 14703 10659
rect 14826 10656 14832 10668
rect 14691 10628 14832 10656
rect 14691 10625 14703 10628
rect 14645 10619 14703 10625
rect 14826 10616 14832 10628
rect 14884 10656 14890 10668
rect 15654 10656 15660 10668
rect 14884 10628 15660 10656
rect 14884 10616 14890 10628
rect 15654 10616 15660 10628
rect 15712 10656 15718 10668
rect 17052 10665 17080 10696
rect 17954 10684 17960 10696
rect 18012 10684 18018 10736
rect 18141 10727 18199 10733
rect 18141 10693 18153 10727
rect 18187 10724 18199 10727
rect 18601 10727 18659 10733
rect 18601 10724 18613 10727
rect 18187 10696 18613 10724
rect 18187 10693 18199 10696
rect 18141 10687 18199 10693
rect 18601 10693 18613 10696
rect 18647 10693 18659 10727
rect 19978 10724 19984 10736
rect 19826 10696 19984 10724
rect 18601 10687 18659 10693
rect 19978 10684 19984 10696
rect 20036 10684 20042 10736
rect 21453 10727 21511 10733
rect 21453 10724 21465 10727
rect 20364 10696 21465 10724
rect 16853 10659 16911 10665
rect 16853 10656 16865 10659
rect 15712 10628 16865 10656
rect 15712 10616 15718 10628
rect 16853 10625 16865 10628
rect 16899 10625 16911 10659
rect 16853 10619 16911 10625
rect 17037 10659 17095 10665
rect 17037 10625 17049 10659
rect 17083 10625 17095 10659
rect 18046 10656 18052 10668
rect 17037 10619 17095 10625
rect 17144 10628 18052 10656
rect 13173 10591 13231 10597
rect 13173 10588 13185 10591
rect 13004 10560 13185 10588
rect 13173 10557 13185 10560
rect 13219 10557 13231 10591
rect 13173 10551 13231 10557
rect 13188 10520 13216 10551
rect 16114 10548 16120 10600
rect 16172 10588 16178 10600
rect 17052 10588 17080 10619
rect 16172 10560 17080 10588
rect 16172 10548 16178 10560
rect 14090 10520 14096 10532
rect 13188 10492 14096 10520
rect 14090 10480 14096 10492
rect 14148 10520 14154 10532
rect 15562 10520 15568 10532
rect 14148 10492 15568 10520
rect 14148 10480 14154 10492
rect 15562 10480 15568 10492
rect 15620 10520 15626 10532
rect 17144 10520 17172 10628
rect 18046 10616 18052 10628
rect 18104 10616 18110 10668
rect 18230 10616 18236 10668
rect 18288 10616 18294 10668
rect 20364 10665 20392 10696
rect 21453 10693 21465 10696
rect 21499 10724 21511 10727
rect 22066 10724 22100 10736
rect 21499 10696 22100 10724
rect 21499 10693 21511 10696
rect 21453 10687 21511 10693
rect 22094 10684 22100 10696
rect 22152 10684 22158 10736
rect 22922 10684 22928 10736
rect 22980 10684 22986 10736
rect 26602 10724 26608 10736
rect 26450 10696 26608 10724
rect 26602 10684 26608 10696
rect 26660 10724 26666 10736
rect 27172 10724 27200 10755
rect 27890 10752 27896 10804
rect 27948 10752 27954 10804
rect 28442 10752 28448 10804
rect 28500 10752 28506 10804
rect 28905 10795 28963 10801
rect 28905 10761 28917 10795
rect 28951 10761 28963 10795
rect 28905 10755 28963 10761
rect 29089 10795 29147 10801
rect 29089 10761 29101 10795
rect 29135 10792 29147 10795
rect 29546 10792 29552 10804
rect 29135 10764 29552 10792
rect 29135 10761 29147 10764
rect 29089 10755 29147 10761
rect 26660 10696 27200 10724
rect 27908 10724 27936 10752
rect 28460 10724 28488 10752
rect 28629 10727 28687 10733
rect 28629 10724 28641 10727
rect 27908 10696 28304 10724
rect 28460 10696 28641 10724
rect 26660 10684 26666 10696
rect 20349 10659 20407 10665
rect 20349 10625 20361 10659
rect 20395 10625 20407 10659
rect 20349 10619 20407 10625
rect 20714 10616 20720 10668
rect 20772 10656 20778 10668
rect 20772 10628 21312 10656
rect 20772 10616 20778 10628
rect 18322 10548 18328 10600
rect 18380 10548 18386 10600
rect 19242 10548 19248 10600
rect 19300 10588 19306 10600
rect 20809 10591 20867 10597
rect 20809 10588 20821 10591
rect 19300 10560 20821 10588
rect 19300 10548 19306 10560
rect 20809 10557 20821 10560
rect 20855 10557 20867 10591
rect 21284 10588 21312 10628
rect 21358 10616 21364 10668
rect 21416 10616 21422 10668
rect 21637 10659 21695 10665
rect 21637 10625 21649 10659
rect 21683 10625 21695 10659
rect 21637 10619 21695 10625
rect 21652 10588 21680 10619
rect 26510 10616 26516 10668
rect 26568 10656 26574 10668
rect 27065 10659 27123 10665
rect 27065 10656 27077 10659
rect 26568 10628 27077 10656
rect 26568 10616 26574 10628
rect 27065 10625 27077 10628
rect 27111 10656 27123 10659
rect 27246 10656 27252 10668
rect 27111 10628 27252 10656
rect 27111 10625 27123 10628
rect 27065 10619 27123 10625
rect 27246 10616 27252 10628
rect 27304 10616 27310 10668
rect 27801 10659 27859 10665
rect 27801 10625 27813 10659
rect 27847 10625 27859 10659
rect 27801 10619 27859 10625
rect 21284 10560 21680 10588
rect 20809 10551 20867 10557
rect 15620 10492 17172 10520
rect 17221 10523 17279 10529
rect 15620 10480 15626 10492
rect 17221 10489 17233 10523
rect 17267 10489 17279 10523
rect 20254 10520 20260 10532
rect 17221 10483 17279 10489
rect 20088 10492 20260 10520
rect 13446 10412 13452 10464
rect 13504 10412 13510 10464
rect 13725 10455 13783 10461
rect 13725 10421 13737 10455
rect 13771 10452 13783 10455
rect 14826 10452 14832 10464
rect 13771 10424 14832 10452
rect 13771 10421 13783 10424
rect 13725 10415 13783 10421
rect 14826 10412 14832 10424
rect 14884 10412 14890 10464
rect 17236 10452 17264 10483
rect 19886 10452 19892 10464
rect 17236 10424 19892 10452
rect 19886 10412 19892 10424
rect 19944 10452 19950 10464
rect 20088 10461 20116 10492
rect 20254 10480 20260 10492
rect 20312 10520 20318 10532
rect 21652 10520 21680 10560
rect 22830 10548 22836 10600
rect 22888 10588 22894 10600
rect 23477 10591 23535 10597
rect 23477 10588 23489 10591
rect 22888 10560 23489 10588
rect 22888 10548 22894 10560
rect 23477 10557 23489 10560
rect 23523 10557 23535 10591
rect 23477 10551 23535 10557
rect 23753 10591 23811 10597
rect 23753 10557 23765 10591
rect 23799 10588 23811 10591
rect 23934 10588 23940 10600
rect 23799 10560 23940 10588
rect 23799 10557 23811 10560
rect 23753 10551 23811 10557
rect 23934 10548 23940 10560
rect 23992 10548 23998 10600
rect 24946 10548 24952 10600
rect 25004 10548 25010 10600
rect 25225 10591 25283 10597
rect 25225 10557 25237 10591
rect 25271 10588 25283 10591
rect 25866 10588 25872 10600
rect 25271 10560 25872 10588
rect 25271 10557 25283 10560
rect 25225 10551 25283 10557
rect 25866 10548 25872 10560
rect 25924 10548 25930 10600
rect 27816 10588 27844 10619
rect 27982 10616 27988 10668
rect 28040 10616 28046 10668
rect 28276 10665 28304 10696
rect 28629 10693 28641 10696
rect 28675 10693 28687 10727
rect 28920 10724 28948 10755
rect 29546 10752 29552 10764
rect 29604 10752 29610 10804
rect 29641 10795 29699 10801
rect 29641 10761 29653 10795
rect 29687 10792 29699 10795
rect 30190 10792 30196 10804
rect 29687 10764 30196 10792
rect 29687 10761 29699 10764
rect 29641 10755 29699 10761
rect 30190 10752 30196 10764
rect 30248 10752 30254 10804
rect 31389 10795 31447 10801
rect 31389 10761 31401 10795
rect 31435 10792 31447 10795
rect 31754 10792 31760 10804
rect 31435 10764 31760 10792
rect 31435 10761 31447 10764
rect 31389 10755 31447 10761
rect 31754 10752 31760 10764
rect 31812 10752 31818 10804
rect 32674 10752 32680 10804
rect 32732 10752 32738 10804
rect 32766 10752 32772 10804
rect 32824 10792 32830 10804
rect 32953 10795 33011 10801
rect 32953 10792 32965 10795
rect 32824 10764 32965 10792
rect 32824 10752 32830 10764
rect 32953 10761 32965 10764
rect 32999 10761 33011 10795
rect 32953 10755 33011 10761
rect 34790 10752 34796 10804
rect 34848 10792 34854 10804
rect 35345 10795 35403 10801
rect 35345 10792 35357 10795
rect 34848 10764 35357 10792
rect 34848 10752 34854 10764
rect 35345 10761 35357 10764
rect 35391 10761 35403 10795
rect 35345 10755 35403 10761
rect 36170 10752 36176 10804
rect 36228 10752 36234 10804
rect 37090 10752 37096 10804
rect 37148 10752 37154 10804
rect 37366 10752 37372 10804
rect 37424 10752 37430 10804
rect 37987 10795 38045 10801
rect 37987 10792 37999 10795
rect 37568 10764 37999 10792
rect 28920 10696 29316 10724
rect 28629 10687 28687 10693
rect 28261 10659 28319 10665
rect 28261 10625 28273 10659
rect 28307 10625 28319 10659
rect 28261 10619 28319 10625
rect 28350 10616 28356 10668
rect 28408 10656 28414 10668
rect 28408 10628 28453 10656
rect 28408 10616 28414 10628
rect 28534 10616 28540 10668
rect 28592 10616 28598 10668
rect 28767 10659 28825 10665
rect 28767 10625 28779 10659
rect 28813 10656 28825 10659
rect 28902 10656 28908 10668
rect 28813 10628 28908 10656
rect 28813 10625 28825 10628
rect 28767 10619 28825 10625
rect 28902 10616 28908 10628
rect 28960 10616 28966 10668
rect 28997 10659 29055 10665
rect 28997 10625 29009 10659
rect 29043 10625 29055 10659
rect 28997 10619 29055 10625
rect 29012 10588 29040 10619
rect 29178 10616 29184 10668
rect 29236 10616 29242 10668
rect 29288 10665 29316 10696
rect 30742 10684 30748 10736
rect 30800 10684 30806 10736
rect 30837 10727 30895 10733
rect 30837 10693 30849 10727
rect 30883 10724 30895 10727
rect 31018 10724 31024 10736
rect 30883 10696 31024 10724
rect 30883 10693 30895 10696
rect 30837 10687 30895 10693
rect 31018 10684 31024 10696
rect 31076 10684 31082 10736
rect 34882 10724 34888 10736
rect 32600 10696 32904 10724
rect 32600 10668 32628 10696
rect 29273 10659 29331 10665
rect 29273 10625 29285 10659
rect 29319 10625 29331 10659
rect 29273 10619 29331 10625
rect 29454 10616 29460 10668
rect 29512 10616 29518 10668
rect 30374 10616 30380 10668
rect 30432 10656 30438 10668
rect 31113 10659 31171 10665
rect 31113 10656 31125 10659
rect 30432 10628 31125 10656
rect 30432 10616 30438 10628
rect 31113 10625 31125 10628
rect 31159 10656 31171 10659
rect 31159 10628 32536 10656
rect 31159 10625 31171 10628
rect 31113 10619 31171 10625
rect 29086 10588 29092 10600
rect 27816 10560 29092 10588
rect 29086 10548 29092 10560
rect 29144 10588 29150 10600
rect 31018 10588 31024 10600
rect 29144 10560 31024 10588
rect 29144 10548 29150 10560
rect 31018 10548 31024 10560
rect 31076 10548 31082 10600
rect 31202 10548 31208 10600
rect 31260 10548 31266 10600
rect 32508 10588 32536 10628
rect 32582 10616 32588 10668
rect 32640 10616 32646 10668
rect 32766 10616 32772 10668
rect 32824 10616 32830 10668
rect 32876 10665 32904 10696
rect 32968 10696 34888 10724
rect 32861 10659 32919 10665
rect 32861 10625 32873 10659
rect 32907 10625 32919 10659
rect 32861 10619 32919 10625
rect 32968 10588 32996 10696
rect 34882 10684 34888 10696
rect 34940 10684 34946 10736
rect 35066 10684 35072 10736
rect 35124 10684 35130 10736
rect 36078 10724 36084 10736
rect 35544 10696 36084 10724
rect 33042 10616 33048 10668
rect 33100 10616 33106 10668
rect 34422 10616 34428 10668
rect 34480 10616 34486 10668
rect 35342 10616 35348 10668
rect 35400 10656 35406 10668
rect 35544 10665 35572 10696
rect 36078 10684 36084 10696
rect 36136 10684 36142 10736
rect 36188 10724 36216 10752
rect 36188 10696 36584 10724
rect 35529 10659 35587 10665
rect 35529 10656 35541 10659
rect 35400 10628 35541 10656
rect 35400 10616 35406 10628
rect 35529 10625 35541 10628
rect 35575 10625 35587 10659
rect 35529 10619 35587 10625
rect 35618 10616 35624 10668
rect 35676 10616 35682 10668
rect 35894 10616 35900 10668
rect 35952 10616 35958 10668
rect 36173 10659 36231 10665
rect 36173 10625 36185 10659
rect 36219 10625 36231 10659
rect 36173 10619 36231 10625
rect 36265 10659 36323 10665
rect 36265 10625 36277 10659
rect 36311 10625 36323 10659
rect 36265 10619 36323 10625
rect 32508 10560 32996 10588
rect 34517 10591 34575 10597
rect 34517 10557 34529 10591
rect 34563 10588 34575 10591
rect 36188 10588 36216 10619
rect 34563 10560 36216 10588
rect 36280 10588 36308 10619
rect 36446 10616 36452 10668
rect 36504 10616 36510 10668
rect 36556 10665 36584 10696
rect 36541 10659 36599 10665
rect 36541 10625 36553 10659
rect 36587 10625 36599 10659
rect 36541 10619 36599 10625
rect 36630 10616 36636 10668
rect 36688 10656 36694 10668
rect 37108 10656 37136 10752
rect 37182 10684 37188 10736
rect 37240 10724 37246 10736
rect 37568 10733 37596 10764
rect 37987 10761 37999 10764
rect 38033 10761 38045 10795
rect 37987 10755 38045 10761
rect 39025 10795 39083 10801
rect 39025 10761 39037 10795
rect 39071 10792 39083 10795
rect 39574 10792 39580 10804
rect 39071 10764 39580 10792
rect 39071 10761 39083 10764
rect 39025 10755 39083 10761
rect 39574 10752 39580 10764
rect 39632 10752 39638 10804
rect 37553 10727 37611 10733
rect 37553 10724 37565 10727
rect 37240 10696 37565 10724
rect 37240 10684 37246 10696
rect 37553 10693 37565 10696
rect 37599 10693 37611 10727
rect 37553 10687 37611 10693
rect 37737 10727 37795 10733
rect 37737 10693 37749 10727
rect 37783 10693 37795 10727
rect 37737 10687 37795 10693
rect 37752 10656 37780 10687
rect 38194 10684 38200 10736
rect 38252 10684 38258 10736
rect 38378 10684 38384 10736
rect 38436 10724 38442 10736
rect 39393 10727 39451 10733
rect 39393 10724 39405 10727
rect 38436 10696 39405 10724
rect 38436 10684 38442 10696
rect 39393 10693 39405 10696
rect 39439 10693 39451 10727
rect 39393 10687 39451 10693
rect 36688 10628 37780 10656
rect 38212 10656 38240 10684
rect 38470 10656 38476 10668
rect 38212 10628 38476 10656
rect 36688 10616 36694 10628
rect 38470 10616 38476 10628
rect 38528 10656 38534 10668
rect 38933 10659 38991 10665
rect 38933 10656 38945 10659
rect 38528 10628 38945 10656
rect 38528 10616 38534 10628
rect 38933 10625 38945 10628
rect 38979 10625 38991 10659
rect 38933 10619 38991 10625
rect 39117 10659 39175 10665
rect 39117 10625 39129 10659
rect 39163 10625 39175 10659
rect 39117 10619 39175 10625
rect 38286 10588 38292 10600
rect 36280 10560 38292 10588
rect 34563 10557 34575 10560
rect 34517 10551 34575 10557
rect 22002 10520 22008 10532
rect 20312 10492 20392 10520
rect 21652 10492 22008 10520
rect 20312 10480 20318 10492
rect 20364 10461 20392 10492
rect 22002 10480 22008 10492
rect 22060 10480 22066 10532
rect 20073 10455 20131 10461
rect 20073 10452 20085 10455
rect 19944 10424 20085 10452
rect 19944 10412 19950 10424
rect 20073 10421 20085 10424
rect 20119 10421 20131 10455
rect 20073 10415 20131 10421
rect 20349 10455 20407 10461
rect 20349 10421 20361 10455
rect 20395 10421 20407 10455
rect 20349 10415 20407 10421
rect 21634 10412 21640 10464
rect 21692 10412 21698 10464
rect 24964 10452 24992 10548
rect 28718 10520 28724 10532
rect 26252 10492 28724 10520
rect 26252 10452 26280 10492
rect 28718 10480 28724 10492
rect 28776 10480 28782 10532
rect 31754 10520 31760 10532
rect 28828 10492 31760 10520
rect 24964 10424 26280 10452
rect 27246 10412 27252 10464
rect 27304 10452 27310 10464
rect 27617 10455 27675 10461
rect 27617 10452 27629 10455
rect 27304 10424 27629 10452
rect 27304 10412 27310 10424
rect 27617 10421 27629 10424
rect 27663 10452 27675 10455
rect 28828 10452 28856 10492
rect 31754 10480 31760 10492
rect 31812 10480 31818 10532
rect 34698 10480 34704 10532
rect 34756 10520 34762 10532
rect 35618 10520 35624 10532
rect 34756 10492 35624 10520
rect 34756 10480 34762 10492
rect 35618 10480 35624 10492
rect 35676 10480 35682 10532
rect 36280 10520 36308 10560
rect 38286 10548 38292 10560
rect 38344 10588 38350 10600
rect 39132 10588 39160 10619
rect 39298 10616 39304 10668
rect 39356 10616 39362 10668
rect 39485 10659 39543 10665
rect 39485 10625 39497 10659
rect 39531 10656 39543 10659
rect 40586 10656 40592 10668
rect 39531 10628 40592 10656
rect 39531 10625 39543 10628
rect 39485 10619 39543 10625
rect 40586 10616 40592 10628
rect 40644 10616 40650 10668
rect 38344 10560 39160 10588
rect 38344 10548 38350 10560
rect 35728 10492 36308 10520
rect 37568 10492 38056 10520
rect 27663 10424 28856 10452
rect 27663 10421 27675 10424
rect 27617 10415 27675 10421
rect 29454 10412 29460 10464
rect 29512 10412 29518 10464
rect 30466 10412 30472 10464
rect 30524 10452 30530 10464
rect 32306 10452 32312 10464
rect 30524 10424 32312 10452
rect 30524 10412 30530 10424
rect 32306 10412 32312 10424
rect 32364 10412 32370 10464
rect 34606 10412 34612 10464
rect 34664 10452 34670 10464
rect 35069 10455 35127 10461
rect 35069 10452 35081 10455
rect 34664 10424 35081 10452
rect 34664 10412 34670 10424
rect 35069 10421 35081 10424
rect 35115 10421 35127 10455
rect 35069 10415 35127 10421
rect 35253 10455 35311 10461
rect 35253 10421 35265 10455
rect 35299 10452 35311 10455
rect 35728 10452 35756 10492
rect 37568 10464 37596 10492
rect 35299 10424 35756 10452
rect 35299 10421 35311 10424
rect 35253 10415 35311 10421
rect 35802 10412 35808 10464
rect 35860 10412 35866 10464
rect 35894 10412 35900 10464
rect 35952 10452 35958 10464
rect 35989 10455 36047 10461
rect 35989 10452 36001 10455
rect 35952 10424 36001 10452
rect 35952 10412 35958 10424
rect 35989 10421 36001 10424
rect 36035 10421 36047 10455
rect 35989 10415 36047 10421
rect 36078 10412 36084 10464
rect 36136 10452 36142 10464
rect 37458 10452 37464 10464
rect 36136 10424 37464 10452
rect 36136 10412 36142 10424
rect 37458 10412 37464 10424
rect 37516 10412 37522 10464
rect 37550 10412 37556 10464
rect 37608 10412 37614 10464
rect 37826 10412 37832 10464
rect 37884 10412 37890 10464
rect 38028 10461 38056 10492
rect 38013 10455 38071 10461
rect 38013 10421 38025 10455
rect 38059 10421 38071 10455
rect 38013 10415 38071 10421
rect 1104 10362 58880 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 58880 10362
rect 1104 10288 58880 10310
rect 14461 10251 14519 10257
rect 14461 10248 14473 10251
rect 13464 10220 14473 10248
rect 12437 10115 12495 10121
rect 12437 10081 12449 10115
rect 12483 10112 12495 10115
rect 13464 10112 13492 10220
rect 14461 10217 14473 10220
rect 14507 10217 14519 10251
rect 17310 10248 17316 10260
rect 14461 10211 14519 10217
rect 16500 10220 17316 10248
rect 13538 10140 13544 10192
rect 13596 10140 13602 10192
rect 13906 10140 13912 10192
rect 13964 10140 13970 10192
rect 14369 10183 14427 10189
rect 14369 10149 14381 10183
rect 14415 10149 14427 10183
rect 14369 10143 14427 10149
rect 12483 10084 13492 10112
rect 13556 10112 13584 10140
rect 14384 10112 14412 10143
rect 16209 10115 16267 10121
rect 13556 10084 14228 10112
rect 14384 10084 14688 10112
rect 12483 10081 12495 10084
rect 12437 10075 12495 10081
rect 12161 10047 12219 10053
rect 12161 10013 12173 10047
rect 12207 10013 12219 10047
rect 12161 10007 12219 10013
rect 12176 9976 12204 10007
rect 14090 10004 14096 10056
rect 14148 10004 14154 10056
rect 14200 10044 14228 10084
rect 14660 10053 14688 10084
rect 16209 10081 16221 10115
rect 16255 10112 16267 10115
rect 16500 10112 16528 10220
rect 17310 10208 17316 10220
rect 17368 10208 17374 10260
rect 17954 10208 17960 10260
rect 18012 10248 18018 10260
rect 18325 10251 18383 10257
rect 18325 10248 18337 10251
rect 18012 10220 18337 10248
rect 18012 10208 18018 10220
rect 18325 10217 18337 10220
rect 18371 10217 18383 10251
rect 18325 10211 18383 10217
rect 22002 10208 22008 10260
rect 22060 10248 22066 10260
rect 22373 10251 22431 10257
rect 22373 10248 22385 10251
rect 22060 10220 22385 10248
rect 22060 10208 22066 10220
rect 22373 10217 22385 10220
rect 22419 10217 22431 10251
rect 22373 10211 22431 10217
rect 22554 10208 22560 10260
rect 22612 10208 22618 10260
rect 22830 10208 22836 10260
rect 22888 10208 22894 10260
rect 25866 10208 25872 10260
rect 25924 10208 25930 10260
rect 27706 10208 27712 10260
rect 27764 10208 27770 10260
rect 29273 10251 29331 10257
rect 29273 10217 29285 10251
rect 29319 10248 29331 10251
rect 29362 10248 29368 10260
rect 29319 10220 29368 10248
rect 29319 10217 29331 10220
rect 29273 10211 29331 10217
rect 29362 10208 29368 10220
rect 29420 10208 29426 10260
rect 29454 10208 29460 10260
rect 29512 10248 29518 10260
rect 29917 10251 29975 10257
rect 29917 10248 29929 10251
rect 29512 10220 29929 10248
rect 29512 10208 29518 10220
rect 29917 10217 29929 10220
rect 29963 10217 29975 10251
rect 30466 10248 30472 10260
rect 29917 10211 29975 10217
rect 30397 10220 30472 10248
rect 18046 10140 18052 10192
rect 18104 10180 18110 10192
rect 19889 10183 19947 10189
rect 19889 10180 19901 10183
rect 18104 10152 19901 10180
rect 18104 10140 18110 10152
rect 19889 10149 19901 10152
rect 19935 10149 19947 10183
rect 19889 10143 19947 10149
rect 21634 10140 21640 10192
rect 21692 10180 21698 10192
rect 22741 10183 22799 10189
rect 22741 10180 22753 10183
rect 21692 10152 22753 10180
rect 21692 10140 21698 10152
rect 22741 10149 22753 10152
rect 22787 10149 22799 10183
rect 27614 10180 27620 10192
rect 22741 10143 22799 10149
rect 26160 10152 27620 10180
rect 16255 10084 16528 10112
rect 16577 10115 16635 10121
rect 16255 10081 16267 10084
rect 16209 10075 16267 10081
rect 16577 10081 16589 10115
rect 16623 10112 16635 10115
rect 18322 10112 18328 10124
rect 16623 10084 18328 10112
rect 16623 10081 16635 10084
rect 16577 10075 16635 10081
rect 18322 10072 18328 10084
rect 18380 10072 18386 10124
rect 22925 10115 22983 10121
rect 22925 10081 22937 10115
rect 22971 10112 22983 10115
rect 23106 10112 23112 10124
rect 22971 10084 23112 10112
rect 22971 10081 22983 10084
rect 22925 10075 22983 10081
rect 23106 10072 23112 10084
rect 23164 10072 23170 10124
rect 14461 10047 14519 10053
rect 14461 10044 14473 10047
rect 14200 10016 14473 10044
rect 14461 10013 14473 10016
rect 14507 10013 14519 10047
rect 14461 10007 14519 10013
rect 14645 10047 14703 10053
rect 14645 10013 14657 10047
rect 14691 10013 14703 10047
rect 14645 10007 14703 10013
rect 16114 10004 16120 10056
rect 16172 10004 16178 10056
rect 18785 10047 18843 10053
rect 18785 10013 18797 10047
rect 18831 10044 18843 10047
rect 19978 10044 19984 10056
rect 18831 10016 19984 10044
rect 18831 10013 18843 10016
rect 18785 10007 18843 10013
rect 19978 10004 19984 10016
rect 20036 10004 20042 10056
rect 20070 10004 20076 10056
rect 20128 10044 20134 10056
rect 20165 10047 20223 10053
rect 20165 10044 20177 10047
rect 20128 10016 20177 10044
rect 20128 10004 20134 10016
rect 20165 10013 20177 10016
rect 20211 10013 20223 10047
rect 20165 10007 20223 10013
rect 20254 10004 20260 10056
rect 20312 10004 20318 10056
rect 22554 10004 22560 10056
rect 22612 10044 22618 10056
rect 22649 10047 22707 10053
rect 22649 10044 22661 10047
rect 22612 10016 22661 10044
rect 22612 10004 22618 10016
rect 22649 10013 22661 10016
rect 22695 10013 22707 10047
rect 22649 10007 22707 10013
rect 23014 10004 23020 10056
rect 23072 10004 23078 10056
rect 26160 10053 26188 10152
rect 27614 10140 27620 10152
rect 27672 10140 27678 10192
rect 30397 10180 30425 10220
rect 30466 10208 30472 10220
rect 30524 10208 30530 10260
rect 30926 10208 30932 10260
rect 30984 10248 30990 10260
rect 31021 10251 31079 10257
rect 31021 10248 31033 10251
rect 30984 10220 31033 10248
rect 30984 10208 30990 10220
rect 31021 10217 31033 10220
rect 31067 10217 31079 10251
rect 31021 10211 31079 10217
rect 31113 10251 31171 10257
rect 31113 10217 31125 10251
rect 31159 10248 31171 10251
rect 31202 10248 31208 10260
rect 31159 10220 31208 10248
rect 31159 10217 31171 10220
rect 31113 10211 31171 10217
rect 31128 10180 31156 10211
rect 31202 10208 31208 10220
rect 31260 10208 31266 10260
rect 32033 10251 32091 10257
rect 32033 10217 32045 10251
rect 32079 10248 32091 10251
rect 32214 10248 32220 10260
rect 32079 10220 32220 10248
rect 32079 10217 32091 10220
rect 32033 10211 32091 10217
rect 32214 10208 32220 10220
rect 32272 10208 32278 10260
rect 32950 10208 32956 10260
rect 33008 10248 33014 10260
rect 35342 10248 35348 10260
rect 33008 10220 35348 10248
rect 33008 10208 33014 10220
rect 28966 10152 30425 10180
rect 30760 10152 31156 10180
rect 26237 10115 26295 10121
rect 26237 10081 26249 10115
rect 26283 10112 26295 10115
rect 27249 10115 27307 10121
rect 27249 10112 27261 10115
rect 26283 10084 27261 10112
rect 26283 10081 26295 10084
rect 26237 10075 26295 10081
rect 27249 10081 27261 10084
rect 27295 10081 27307 10115
rect 27632 10112 27660 10140
rect 28966 10112 28994 10152
rect 27632 10084 28994 10112
rect 27249 10075 27307 10081
rect 30374 10072 30380 10124
rect 30432 10072 30438 10124
rect 30466 10072 30472 10124
rect 30524 10112 30530 10124
rect 30561 10115 30619 10121
rect 30561 10112 30573 10115
rect 30524 10084 30573 10112
rect 30524 10072 30530 10084
rect 30561 10081 30573 10084
rect 30607 10081 30619 10115
rect 30561 10075 30619 10081
rect 23201 10047 23259 10053
rect 23201 10013 23213 10047
rect 23247 10013 23259 10047
rect 23201 10007 23259 10013
rect 26145 10047 26203 10053
rect 26145 10013 26157 10047
rect 26191 10013 26203 10047
rect 26145 10007 26203 10013
rect 27157 10047 27215 10053
rect 27157 10013 27169 10047
rect 27203 10013 27215 10047
rect 27157 10007 27215 10013
rect 12342 9976 12348 9988
rect 12176 9948 12348 9976
rect 12342 9936 12348 9948
rect 12400 9936 12406 9988
rect 13722 9976 13728 9988
rect 13662 9948 13728 9976
rect 13722 9936 13728 9948
rect 13780 9936 13786 9988
rect 13906 9936 13912 9988
rect 13964 9976 13970 9988
rect 14369 9979 14427 9985
rect 14369 9976 14381 9979
rect 13964 9948 14381 9976
rect 13964 9936 13970 9948
rect 14369 9945 14381 9948
rect 14415 9945 14427 9979
rect 14369 9939 14427 9945
rect 16850 9936 16856 9988
rect 16908 9936 16914 9988
rect 18417 9979 18475 9985
rect 18417 9976 18429 9979
rect 18078 9948 18429 9976
rect 14185 9911 14243 9917
rect 14185 9877 14197 9911
rect 14231 9908 14243 9911
rect 14826 9908 14832 9920
rect 14231 9880 14832 9908
rect 14231 9877 14243 9880
rect 14185 9871 14243 9877
rect 14826 9868 14832 9880
rect 14884 9868 14890 9920
rect 16485 9911 16543 9917
rect 16485 9877 16497 9911
rect 16531 9908 16543 9911
rect 16758 9908 16764 9920
rect 16531 9880 16764 9908
rect 16531 9877 16543 9880
rect 16485 9871 16543 9877
rect 16758 9868 16764 9880
rect 16816 9868 16822 9920
rect 17678 9868 17684 9920
rect 17736 9908 17742 9920
rect 18156 9908 18184 9948
rect 18417 9945 18429 9948
rect 18463 9945 18475 9979
rect 18417 9939 18475 9945
rect 20441 9979 20499 9985
rect 20441 9945 20453 9979
rect 20487 9976 20499 9979
rect 22094 9976 22100 9988
rect 20487 9948 22100 9976
rect 20487 9945 20499 9948
rect 20441 9939 20499 9945
rect 22094 9936 22100 9948
rect 22152 9976 22158 9988
rect 22189 9979 22247 9985
rect 22189 9976 22201 9979
rect 22152 9948 22201 9976
rect 22152 9936 22158 9948
rect 22189 9945 22201 9948
rect 22235 9945 22247 9979
rect 23216 9976 23244 10007
rect 22189 9939 22247 9945
rect 23032 9948 23244 9976
rect 17736 9880 18184 9908
rect 20073 9911 20131 9917
rect 17736 9868 17742 9880
rect 20073 9877 20085 9911
rect 20119 9908 20131 9911
rect 21358 9908 21364 9920
rect 20119 9880 21364 9908
rect 20119 9877 20131 9880
rect 20073 9871 20131 9877
rect 21358 9868 21364 9880
rect 21416 9868 21422 9920
rect 22370 9868 22376 9920
rect 22428 9917 22434 9920
rect 22428 9911 22447 9917
rect 22435 9908 22447 9911
rect 23032 9908 23060 9948
rect 22435 9880 23060 9908
rect 23109 9911 23167 9917
rect 22435 9877 22447 9880
rect 22428 9871 22447 9877
rect 23109 9877 23121 9911
rect 23155 9908 23167 9911
rect 23658 9908 23664 9920
rect 23155 9880 23664 9908
rect 23155 9877 23167 9880
rect 23109 9871 23167 9877
rect 22428 9868 22434 9871
rect 23658 9868 23664 9880
rect 23716 9868 23722 9920
rect 27172 9908 27200 10007
rect 27338 10004 27344 10056
rect 27396 10004 27402 10056
rect 27706 10004 27712 10056
rect 27764 10044 27770 10056
rect 27801 10047 27859 10053
rect 27801 10044 27813 10047
rect 27764 10016 27813 10044
rect 27764 10004 27770 10016
rect 27801 10013 27813 10016
rect 27847 10013 27859 10047
rect 30285 10047 30343 10053
rect 27801 10007 27859 10013
rect 28552 10016 30236 10044
rect 27356 9976 27384 10004
rect 28552 9976 28580 10016
rect 27356 9948 28580 9976
rect 28629 9979 28687 9985
rect 28629 9945 28641 9979
rect 28675 9976 28687 9979
rect 28718 9976 28724 9988
rect 28675 9948 28724 9976
rect 28675 9945 28687 9948
rect 28629 9939 28687 9945
rect 28718 9936 28724 9948
rect 28776 9936 28782 9988
rect 28905 9979 28963 9985
rect 28905 9945 28917 9979
rect 28951 9976 28963 9979
rect 28994 9976 29000 9988
rect 28951 9948 29000 9976
rect 28951 9945 28963 9948
rect 28905 9939 28963 9945
rect 28994 9936 29000 9948
rect 29052 9936 29058 9988
rect 29086 9936 29092 9988
rect 29144 9936 29150 9988
rect 30208 9976 30236 10016
rect 30285 10013 30297 10047
rect 30331 10044 30343 10047
rect 30760 10044 30788 10152
rect 31294 10140 31300 10192
rect 31352 10180 31358 10192
rect 32122 10180 32128 10192
rect 31352 10152 32128 10180
rect 31352 10140 31358 10152
rect 32122 10140 32128 10152
rect 32180 10140 32186 10192
rect 32232 10152 32996 10180
rect 31478 10112 31484 10124
rect 31036 10084 31484 10112
rect 31036 10053 31064 10084
rect 30331 10016 30788 10044
rect 30837 10047 30895 10053
rect 30331 10013 30343 10016
rect 30285 10007 30343 10013
rect 30837 10013 30849 10047
rect 30883 10013 30895 10047
rect 30837 10007 30895 10013
rect 31021 10047 31079 10053
rect 31021 10013 31033 10047
rect 31067 10013 31079 10047
rect 31021 10007 31079 10013
rect 31113 10047 31171 10053
rect 31113 10013 31125 10047
rect 31159 10044 31171 10047
rect 31202 10044 31208 10056
rect 31159 10016 31208 10044
rect 31159 10013 31171 10016
rect 31113 10007 31171 10013
rect 30852 9976 30880 10007
rect 31202 10004 31208 10016
rect 31260 10004 31266 10056
rect 31312 10053 31340 10084
rect 31478 10072 31484 10084
rect 31536 10112 31542 10124
rect 32232 10112 32260 10152
rect 31536 10084 32260 10112
rect 31536 10072 31542 10084
rect 32306 10072 32312 10124
rect 32364 10112 32370 10124
rect 32401 10115 32459 10121
rect 32401 10112 32413 10115
rect 32364 10084 32413 10112
rect 32364 10072 32370 10084
rect 32401 10081 32413 10084
rect 32447 10081 32459 10115
rect 32401 10075 32459 10081
rect 32674 10072 32680 10124
rect 32732 10072 32738 10124
rect 32968 10121 32996 10152
rect 32953 10115 33011 10121
rect 32953 10081 32965 10115
rect 32999 10081 33011 10115
rect 32953 10075 33011 10081
rect 31297 10047 31355 10053
rect 31297 10013 31309 10047
rect 31343 10013 31355 10047
rect 31297 10007 31355 10013
rect 31938 10004 31944 10056
rect 31996 10044 32002 10056
rect 32033 10047 32091 10053
rect 32033 10044 32045 10047
rect 31996 10016 32045 10044
rect 31996 10004 32002 10016
rect 32033 10013 32045 10016
rect 32079 10013 32091 10047
rect 32033 10007 32091 10013
rect 32217 10047 32275 10053
rect 32217 10013 32229 10047
rect 32263 10013 32275 10047
rect 32217 10007 32275 10013
rect 32493 10047 32551 10053
rect 32493 10013 32505 10047
rect 32539 10013 32551 10047
rect 32493 10007 32551 10013
rect 30208 9948 31754 9976
rect 29104 9908 29132 9936
rect 27172 9880 29132 9908
rect 31726 9908 31754 9948
rect 32030 9908 32036 9920
rect 31726 9880 32036 9908
rect 32030 9868 32036 9880
rect 32088 9868 32094 9920
rect 32232 9908 32260 10007
rect 32306 9936 32312 9988
rect 32364 9976 32370 9988
rect 32508 9976 32536 10007
rect 32582 10004 32588 10056
rect 32640 10044 32646 10056
rect 33244 10053 33272 10220
rect 35342 10208 35348 10220
rect 35400 10208 35406 10260
rect 35802 10208 35808 10260
rect 35860 10248 35866 10260
rect 38102 10248 38108 10260
rect 35860 10220 38108 10248
rect 35860 10208 35866 10220
rect 38102 10208 38108 10220
rect 38160 10208 38166 10260
rect 38289 10251 38347 10257
rect 38289 10217 38301 10251
rect 38335 10248 38347 10251
rect 38562 10248 38568 10260
rect 38335 10220 38568 10248
rect 38335 10217 38347 10220
rect 38289 10211 38347 10217
rect 38562 10208 38568 10220
rect 38620 10208 38626 10260
rect 34790 10140 34796 10192
rect 34848 10180 34854 10192
rect 34848 10152 35572 10180
rect 34848 10140 34854 10152
rect 35544 10121 35572 10152
rect 36170 10140 36176 10192
rect 36228 10140 36234 10192
rect 36262 10140 36268 10192
rect 36320 10180 36326 10192
rect 36725 10183 36783 10189
rect 36725 10180 36737 10183
rect 36320 10152 36737 10180
rect 36320 10140 36326 10152
rect 36725 10149 36737 10152
rect 36771 10149 36783 10183
rect 36725 10143 36783 10149
rect 33413 10115 33471 10121
rect 33413 10081 33425 10115
rect 33459 10112 33471 10115
rect 35437 10115 35495 10121
rect 35437 10112 35449 10115
rect 33459 10084 35449 10112
rect 33459 10081 33471 10084
rect 33413 10075 33471 10081
rect 35437 10081 35449 10084
rect 35483 10081 35495 10115
rect 35437 10075 35495 10081
rect 35529 10115 35587 10121
rect 35529 10081 35541 10115
rect 35575 10081 35587 10115
rect 35529 10075 35587 10081
rect 35894 10072 35900 10124
rect 35952 10072 35958 10124
rect 37108 10084 38148 10112
rect 33045 10047 33103 10053
rect 33045 10044 33057 10047
rect 32640 10016 33057 10044
rect 32640 10004 32646 10016
rect 33045 10013 33057 10016
rect 33091 10013 33103 10047
rect 33045 10007 33103 10013
rect 33229 10047 33287 10053
rect 33229 10013 33241 10047
rect 33275 10013 33287 10047
rect 33778 10044 33784 10056
rect 33229 10007 33287 10013
rect 33428 10016 33784 10044
rect 33428 9976 33456 10016
rect 33778 10004 33784 10016
rect 33836 10004 33842 10056
rect 35345 10047 35403 10053
rect 35345 10013 35357 10047
rect 35391 10044 35403 10047
rect 35391 10016 36308 10044
rect 35391 10013 35403 10016
rect 35345 10007 35403 10013
rect 32364 9948 33456 9976
rect 32364 9936 32370 9948
rect 33686 9936 33692 9988
rect 33744 9976 33750 9988
rect 36170 9976 36176 9988
rect 33744 9948 36176 9976
rect 33744 9936 33750 9948
rect 36170 9936 36176 9948
rect 36228 9936 36234 9988
rect 36280 9976 36308 10016
rect 36354 10004 36360 10056
rect 36412 10044 36418 10056
rect 36541 10047 36599 10053
rect 36412 10016 36457 10044
rect 36412 10004 36418 10016
rect 36541 10013 36553 10047
rect 36587 10044 36599 10047
rect 36909 10047 36967 10053
rect 36909 10044 36921 10047
rect 36587 10016 36921 10044
rect 36587 10013 36599 10016
rect 36541 10007 36599 10013
rect 36909 10013 36921 10016
rect 36955 10013 36967 10047
rect 36909 10007 36967 10013
rect 36446 9976 36452 9988
rect 36280 9948 36452 9976
rect 36446 9936 36452 9948
rect 36504 9936 36510 9988
rect 36633 9979 36691 9985
rect 36633 9945 36645 9979
rect 36679 9976 36691 9979
rect 36924 9976 36952 10007
rect 36998 10004 37004 10056
rect 37056 10044 37062 10056
rect 37108 10053 37136 10084
rect 37093 10047 37151 10053
rect 37093 10044 37105 10047
rect 37056 10016 37105 10044
rect 37056 10004 37062 10016
rect 37093 10013 37105 10016
rect 37139 10013 37151 10047
rect 37093 10007 37151 10013
rect 37182 10004 37188 10056
rect 37240 10004 37246 10056
rect 38120 10053 38148 10084
rect 39206 10072 39212 10124
rect 39264 10072 39270 10124
rect 40126 10112 40132 10124
rect 39316 10084 40132 10112
rect 39316 10053 39344 10084
rect 40126 10072 40132 10084
rect 40184 10072 40190 10124
rect 40586 10072 40592 10124
rect 40644 10112 40650 10124
rect 41230 10112 41236 10124
rect 40644 10084 41236 10112
rect 40644 10072 40650 10084
rect 41230 10072 41236 10084
rect 41288 10112 41294 10124
rect 41969 10115 42027 10121
rect 41969 10112 41981 10115
rect 41288 10084 41981 10112
rect 41288 10072 41294 10084
rect 41969 10081 41981 10084
rect 42015 10081 42027 10115
rect 41969 10075 42027 10081
rect 37921 10047 37979 10053
rect 37921 10013 37933 10047
rect 37967 10013 37979 10047
rect 37921 10007 37979 10013
rect 38105 10047 38163 10053
rect 38105 10013 38117 10047
rect 38151 10013 38163 10047
rect 38105 10007 38163 10013
rect 39301 10047 39359 10053
rect 39301 10013 39313 10047
rect 39347 10013 39359 10047
rect 39301 10007 39359 10013
rect 37274 9976 37280 9988
rect 36679 9948 36860 9976
rect 36924 9948 37280 9976
rect 36679 9945 36691 9948
rect 36633 9939 36691 9945
rect 32766 9908 32772 9920
rect 32232 9880 32772 9908
rect 32766 9868 32772 9880
rect 32824 9868 32830 9920
rect 32861 9911 32919 9917
rect 32861 9877 32873 9911
rect 32907 9908 32919 9911
rect 35802 9908 35808 9920
rect 32907 9880 35808 9908
rect 32907 9877 32919 9880
rect 32861 9871 32919 9877
rect 35802 9868 35808 9880
rect 35860 9868 35866 9920
rect 36078 9868 36084 9920
rect 36136 9908 36142 9920
rect 36648 9908 36676 9939
rect 36136 9880 36676 9908
rect 36832 9908 36860 9948
rect 37274 9936 37280 9948
rect 37332 9976 37338 9988
rect 37550 9976 37556 9988
rect 37332 9948 37556 9976
rect 37332 9936 37338 9948
rect 37550 9936 37556 9948
rect 37608 9976 37614 9988
rect 37936 9976 37964 10007
rect 40034 10004 40040 10056
rect 40092 10044 40098 10056
rect 40221 10047 40279 10053
rect 40221 10044 40233 10047
rect 40092 10016 40233 10044
rect 40092 10004 40098 10016
rect 40221 10013 40233 10016
rect 40267 10013 40279 10047
rect 40221 10007 40279 10013
rect 40497 9979 40555 9985
rect 40497 9976 40509 9979
rect 37608 9948 37964 9976
rect 39684 9948 40509 9976
rect 37608 9936 37614 9948
rect 37090 9908 37096 9920
rect 36832 9880 37096 9908
rect 36136 9868 36142 9880
rect 37090 9868 37096 9880
rect 37148 9868 37154 9920
rect 39684 9917 39712 9948
rect 40497 9945 40509 9948
rect 40543 9945 40555 9979
rect 40497 9939 40555 9945
rect 41506 9936 41512 9988
rect 41564 9936 41570 9988
rect 39669 9911 39727 9917
rect 39669 9877 39681 9911
rect 39715 9877 39727 9911
rect 39669 9871 39727 9877
rect 1104 9818 58880 9840
rect 1104 9766 4874 9818
rect 4926 9766 4938 9818
rect 4990 9766 5002 9818
rect 5054 9766 5066 9818
rect 5118 9766 5130 9818
rect 5182 9766 35594 9818
rect 35646 9766 35658 9818
rect 35710 9766 35722 9818
rect 35774 9766 35786 9818
rect 35838 9766 35850 9818
rect 35902 9766 58880 9818
rect 1104 9744 58880 9766
rect 14826 9664 14832 9716
rect 14884 9664 14890 9716
rect 16850 9664 16856 9716
rect 16908 9664 16914 9716
rect 23290 9664 23296 9716
rect 23348 9704 23354 9716
rect 27706 9704 27712 9716
rect 23348 9676 27712 9704
rect 23348 9664 23354 9676
rect 27706 9664 27712 9676
rect 27764 9664 27770 9716
rect 29270 9664 29276 9716
rect 29328 9664 29334 9716
rect 30285 9707 30343 9713
rect 30285 9673 30297 9707
rect 30331 9704 30343 9707
rect 30374 9704 30380 9716
rect 30331 9676 30380 9704
rect 30331 9673 30343 9676
rect 30285 9667 30343 9673
rect 30374 9664 30380 9676
rect 30432 9664 30438 9716
rect 32582 9704 32588 9716
rect 31726 9676 32588 9704
rect 13357 9639 13415 9645
rect 13357 9605 13369 9639
rect 13403 9636 13415 9639
rect 13446 9636 13452 9648
rect 13403 9608 13452 9636
rect 13403 9605 13415 9608
rect 13357 9599 13415 9605
rect 13446 9596 13452 9608
rect 13504 9596 13510 9648
rect 15470 9636 15476 9648
rect 14582 9622 15476 9636
rect 14568 9608 15476 9622
rect 12342 9460 12348 9512
rect 12400 9500 12406 9512
rect 12434 9500 12440 9512
rect 12400 9472 12440 9500
rect 12400 9460 12406 9472
rect 12434 9460 12440 9472
rect 12492 9500 12498 9512
rect 13081 9503 13139 9509
rect 13081 9500 13093 9503
rect 12492 9472 13093 9500
rect 12492 9460 12498 9472
rect 13081 9469 13093 9472
rect 13127 9469 13139 9503
rect 13081 9463 13139 9469
rect 13722 9460 13728 9512
rect 13780 9500 13786 9512
rect 14568 9500 14596 9608
rect 15470 9596 15476 9608
rect 15528 9596 15534 9648
rect 21928 9608 23520 9636
rect 21928 9580 21956 9608
rect 16758 9528 16764 9580
rect 16816 9528 16822 9580
rect 16942 9528 16948 9580
rect 17000 9528 17006 9580
rect 21818 9528 21824 9580
rect 21876 9528 21882 9580
rect 21910 9528 21916 9580
rect 21968 9528 21974 9580
rect 22097 9571 22155 9577
rect 22097 9537 22109 9571
rect 22143 9568 22155 9571
rect 22189 9571 22247 9577
rect 22189 9568 22201 9571
rect 22143 9540 22201 9568
rect 22143 9537 22155 9540
rect 22097 9531 22155 9537
rect 22189 9537 22201 9540
rect 22235 9537 22247 9571
rect 22189 9531 22247 9537
rect 23492 9512 23520 9608
rect 28994 9596 29000 9648
rect 29052 9636 29058 9648
rect 31726 9636 31754 9676
rect 32582 9664 32588 9676
rect 32640 9664 32646 9716
rect 32950 9664 32956 9716
rect 33008 9704 33014 9716
rect 33008 9676 33180 9704
rect 33008 9664 33014 9676
rect 29052 9608 31754 9636
rect 29052 9596 29058 9608
rect 28718 9528 28724 9580
rect 28776 9528 28782 9580
rect 29086 9528 29092 9580
rect 29144 9528 29150 9580
rect 30392 9577 30420 9608
rect 32030 9596 32036 9648
rect 32088 9636 32094 9648
rect 33152 9636 33180 9676
rect 36464 9676 37044 9704
rect 33965 9639 34023 9645
rect 33965 9636 33977 9639
rect 32088 9608 33088 9636
rect 33152 9608 33977 9636
rect 32088 9596 32094 9608
rect 29365 9571 29423 9577
rect 29365 9537 29377 9571
rect 29411 9568 29423 9571
rect 30193 9571 30251 9577
rect 30193 9568 30205 9571
rect 29411 9540 30205 9568
rect 29411 9537 29423 9540
rect 29365 9531 29423 9537
rect 30193 9537 30205 9540
rect 30239 9537 30251 9571
rect 30193 9531 30251 9537
rect 30377 9571 30435 9577
rect 30377 9537 30389 9571
rect 30423 9537 30435 9571
rect 30377 9531 30435 9537
rect 13780 9472 14596 9500
rect 13780 9460 13786 9472
rect 21726 9460 21732 9512
rect 21784 9500 21790 9512
rect 22741 9503 22799 9509
rect 22741 9500 22753 9503
rect 21784 9472 22753 9500
rect 21784 9460 21790 9472
rect 22741 9469 22753 9472
rect 22787 9469 22799 9503
rect 22741 9463 22799 9469
rect 23474 9460 23480 9512
rect 23532 9460 23538 9512
rect 28810 9460 28816 9512
rect 28868 9500 28874 9512
rect 29380 9500 29408 9531
rect 28868 9472 29408 9500
rect 28868 9460 28874 9472
rect 22097 9435 22155 9441
rect 22097 9401 22109 9435
rect 22143 9432 22155 9435
rect 23014 9432 23020 9444
rect 22143 9404 23020 9432
rect 22143 9401 22155 9404
rect 22097 9395 22155 9401
rect 23014 9392 23020 9404
rect 23072 9392 23078 9444
rect 30208 9432 30236 9531
rect 32122 9528 32128 9580
rect 32180 9568 32186 9580
rect 32217 9571 32275 9577
rect 32217 9568 32229 9571
rect 32180 9540 32229 9568
rect 32180 9528 32186 9540
rect 32217 9537 32229 9540
rect 32263 9537 32275 9571
rect 32217 9531 32275 9537
rect 32493 9571 32551 9577
rect 32493 9537 32505 9571
rect 32539 9537 32551 9571
rect 32493 9531 32551 9537
rect 31478 9460 31484 9512
rect 31536 9500 31542 9512
rect 32508 9500 32536 9531
rect 32582 9528 32588 9580
rect 32640 9528 32646 9580
rect 32950 9528 32956 9580
rect 33008 9528 33014 9580
rect 33060 9577 33088 9608
rect 33965 9605 33977 9608
rect 34011 9605 34023 9639
rect 33965 9599 34023 9605
rect 34149 9639 34207 9645
rect 34149 9605 34161 9639
rect 34195 9636 34207 9639
rect 36464 9636 36492 9676
rect 34195 9608 36492 9636
rect 36541 9639 36599 9645
rect 34195 9605 34207 9608
rect 34149 9599 34207 9605
rect 36541 9605 36553 9639
rect 36587 9636 36599 9639
rect 36906 9636 36912 9648
rect 36587 9608 36912 9636
rect 36587 9605 36599 9608
rect 36541 9599 36599 9605
rect 36906 9596 36912 9608
rect 36964 9596 36970 9648
rect 37016 9636 37044 9676
rect 40126 9664 40132 9716
rect 40184 9704 40190 9716
rect 40681 9707 40739 9713
rect 40681 9704 40693 9707
rect 40184 9676 40693 9704
rect 40184 9664 40190 9676
rect 40681 9673 40693 9676
rect 40727 9673 40739 9707
rect 40681 9667 40739 9673
rect 39206 9636 39212 9648
rect 37016 9608 39212 9636
rect 39206 9596 39212 9608
rect 39264 9596 39270 9648
rect 33045 9571 33103 9577
rect 33045 9537 33057 9571
rect 33091 9537 33103 9571
rect 33045 9531 33103 9537
rect 33226 9528 33232 9580
rect 33284 9528 33290 9580
rect 33321 9571 33379 9577
rect 33321 9537 33333 9571
rect 33367 9537 33379 9571
rect 33321 9531 33379 9537
rect 33336 9500 33364 9531
rect 33778 9528 33784 9580
rect 33836 9528 33842 9580
rect 36449 9571 36507 9577
rect 36449 9537 36461 9571
rect 36495 9568 36507 9571
rect 36630 9568 36636 9580
rect 36495 9540 36636 9568
rect 36495 9537 36507 9540
rect 36449 9531 36507 9537
rect 31536 9472 33364 9500
rect 31536 9460 31542 9472
rect 33410 9460 33416 9512
rect 33468 9500 33474 9512
rect 36556 9509 36584 9540
rect 36630 9528 36636 9540
rect 36688 9528 36694 9580
rect 36817 9571 36875 9577
rect 36817 9537 36829 9571
rect 36863 9537 36875 9571
rect 36817 9531 36875 9537
rect 33505 9503 33563 9509
rect 33505 9500 33517 9503
rect 33468 9472 33517 9500
rect 33468 9460 33474 9472
rect 33505 9469 33517 9472
rect 33551 9469 33563 9503
rect 33505 9463 33563 9469
rect 36541 9503 36599 9509
rect 36541 9469 36553 9503
rect 36587 9500 36599 9503
rect 36832 9500 36860 9531
rect 37090 9528 37096 9580
rect 37148 9528 37154 9580
rect 37274 9528 37280 9580
rect 37332 9568 37338 9580
rect 37553 9571 37611 9577
rect 37553 9568 37565 9571
rect 37332 9540 37565 9568
rect 37332 9528 37338 9540
rect 37553 9537 37565 9540
rect 37599 9537 37611 9571
rect 37553 9531 37611 9537
rect 41230 9528 41236 9580
rect 41288 9528 41294 9580
rect 36587 9472 36621 9500
rect 36832 9472 37688 9500
rect 36587 9469 36599 9472
rect 36541 9463 36599 9469
rect 31846 9432 31852 9444
rect 30208 9404 31852 9432
rect 31846 9392 31852 9404
rect 31904 9392 31910 9444
rect 31938 9392 31944 9444
rect 31996 9432 32002 9444
rect 32582 9432 32588 9444
rect 31996 9404 32588 9432
rect 31996 9392 32002 9404
rect 32582 9392 32588 9404
rect 32640 9432 32646 9444
rect 33689 9435 33747 9441
rect 33689 9432 33701 9435
rect 32640 9404 33701 9432
rect 32640 9392 32646 9404
rect 33689 9401 33701 9404
rect 33735 9401 33747 9435
rect 34698 9432 34704 9444
rect 33689 9395 33747 9401
rect 34072 9404 34704 9432
rect 22462 9324 22468 9376
rect 22520 9364 22526 9376
rect 22925 9367 22983 9373
rect 22925 9364 22937 9367
rect 22520 9336 22937 9364
rect 22520 9324 22526 9336
rect 22925 9333 22937 9336
rect 22971 9333 22983 9367
rect 22925 9327 22983 9333
rect 27982 9324 27988 9376
rect 28040 9364 28046 9376
rect 28810 9364 28816 9376
rect 28040 9336 28816 9364
rect 28040 9324 28046 9336
rect 28810 9324 28816 9336
rect 28868 9364 28874 9376
rect 31202 9364 31208 9376
rect 28868 9336 31208 9364
rect 28868 9324 28874 9336
rect 31202 9324 31208 9336
rect 31260 9364 31266 9376
rect 32306 9364 32312 9376
rect 31260 9336 32312 9364
rect 31260 9324 31266 9336
rect 32306 9324 32312 9336
rect 32364 9324 32370 9376
rect 32398 9324 32404 9376
rect 32456 9364 32462 9376
rect 32769 9367 32827 9373
rect 32769 9364 32781 9367
rect 32456 9336 32781 9364
rect 32456 9324 32462 9336
rect 32769 9333 32781 9336
rect 32815 9333 32827 9367
rect 32769 9327 32827 9333
rect 33410 9324 33416 9376
rect 33468 9324 33474 9376
rect 33505 9367 33563 9373
rect 33505 9333 33517 9367
rect 33551 9364 33563 9367
rect 34072 9364 34100 9404
rect 34698 9392 34704 9404
rect 34756 9392 34762 9444
rect 33551 9336 34100 9364
rect 36725 9367 36783 9373
rect 33551 9333 33563 9336
rect 33505 9327 33563 9333
rect 36725 9333 36737 9367
rect 36771 9364 36783 9367
rect 36814 9364 36820 9376
rect 36771 9336 36820 9364
rect 36771 9333 36783 9336
rect 36725 9327 36783 9333
rect 36814 9324 36820 9336
rect 36872 9364 36878 9376
rect 37660 9373 37688 9472
rect 37001 9367 37059 9373
rect 37001 9364 37013 9367
rect 36872 9336 37013 9364
rect 36872 9324 36878 9336
rect 37001 9333 37013 9336
rect 37047 9333 37059 9367
rect 37001 9327 37059 9333
rect 37645 9367 37703 9373
rect 37645 9333 37657 9367
rect 37691 9364 37703 9367
rect 39390 9364 39396 9376
rect 37691 9336 39396 9364
rect 37691 9333 37703 9336
rect 37645 9327 37703 9333
rect 39390 9324 39396 9336
rect 39448 9324 39454 9376
rect 1104 9274 58880 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 58880 9274
rect 1104 9200 58880 9222
rect 20993 9163 21051 9169
rect 20993 9129 21005 9163
rect 21039 9160 21051 9163
rect 21174 9160 21180 9172
rect 21039 9132 21180 9160
rect 21039 9129 21051 9132
rect 20993 9123 21051 9129
rect 21174 9120 21180 9132
rect 21232 9120 21238 9172
rect 21910 9160 21916 9172
rect 21284 9132 21916 9160
rect 16666 8916 16672 8968
rect 16724 8956 16730 8968
rect 21284 8965 21312 9132
rect 21910 9120 21916 9132
rect 21968 9120 21974 9172
rect 22189 9163 22247 9169
rect 22189 9160 22201 9163
rect 22020 9132 22201 9160
rect 21726 9052 21732 9104
rect 21784 9092 21790 9104
rect 22020 9092 22048 9132
rect 22189 9129 22201 9132
rect 22235 9129 22247 9163
rect 22189 9123 22247 9129
rect 27709 9163 27767 9169
rect 27709 9129 27721 9163
rect 27755 9160 27767 9163
rect 28074 9160 28080 9172
rect 27755 9132 28080 9160
rect 27755 9129 27767 9132
rect 27709 9123 27767 9129
rect 28074 9120 28080 9132
rect 28132 9160 28138 9172
rect 28445 9163 28503 9169
rect 28445 9160 28457 9163
rect 28132 9132 28457 9160
rect 28132 9120 28138 9132
rect 28445 9129 28457 9132
rect 28491 9129 28503 9163
rect 28445 9123 28503 9129
rect 28810 9120 28816 9172
rect 28868 9120 28874 9172
rect 29086 9120 29092 9172
rect 29144 9160 29150 9172
rect 31938 9160 31944 9172
rect 29144 9132 31944 9160
rect 29144 9120 29150 9132
rect 31938 9120 31944 9132
rect 31996 9120 32002 9172
rect 32214 9120 32220 9172
rect 32272 9120 32278 9172
rect 33226 9120 33232 9172
rect 33284 9160 33290 9172
rect 33413 9163 33471 9169
rect 33413 9160 33425 9163
rect 33284 9132 33425 9160
rect 33284 9120 33290 9132
rect 33413 9129 33425 9132
rect 33459 9160 33471 9163
rect 36630 9160 36636 9172
rect 33459 9132 36636 9160
rect 33459 9129 33471 9132
rect 33413 9123 33471 9129
rect 36630 9120 36636 9132
rect 36688 9120 36694 9172
rect 36722 9120 36728 9172
rect 36780 9160 36786 9172
rect 38010 9160 38016 9172
rect 36780 9132 38016 9160
rect 36780 9120 36786 9132
rect 38010 9120 38016 9132
rect 38068 9120 38074 9172
rect 21784 9064 22048 9092
rect 22097 9095 22155 9101
rect 21784 9052 21790 9064
rect 22097 9061 22109 9095
rect 22143 9092 22155 9095
rect 22370 9092 22376 9104
rect 22143 9064 22376 9092
rect 22143 9061 22155 9064
rect 22097 9055 22155 9061
rect 22370 9052 22376 9064
rect 22428 9052 22434 9104
rect 27798 9052 27804 9104
rect 27856 9092 27862 9104
rect 28353 9095 28411 9101
rect 28353 9092 28365 9095
rect 27856 9064 28365 9092
rect 27856 9052 27862 9064
rect 28353 9061 28365 9064
rect 28399 9061 28411 9095
rect 28353 9055 28411 9061
rect 32122 9052 32128 9104
rect 32180 9092 32186 9104
rect 33042 9092 33048 9104
rect 32180 9064 33048 9092
rect 32180 9052 32186 9064
rect 33042 9052 33048 9064
rect 33100 9052 33106 9104
rect 23658 8984 23664 9036
rect 23716 8984 23722 9036
rect 28534 8984 28540 9036
rect 28592 8984 28598 9036
rect 36722 9024 36728 9036
rect 35728 8996 36728 9024
rect 17405 8959 17463 8965
rect 17405 8956 17417 8959
rect 16724 8928 17417 8956
rect 16724 8916 16730 8928
rect 17405 8925 17417 8928
rect 17451 8925 17463 8959
rect 17405 8919 17463 8925
rect 21269 8959 21327 8965
rect 21269 8925 21281 8959
rect 21315 8925 21327 8959
rect 21269 8919 21327 8925
rect 21376 8928 22586 8956
rect 19978 8848 19984 8900
rect 20036 8888 20042 8900
rect 20441 8891 20499 8897
rect 20441 8888 20453 8891
rect 20036 8860 20453 8888
rect 20036 8848 20042 8860
rect 20441 8857 20453 8860
rect 20487 8888 20499 8891
rect 21376 8888 21404 8928
rect 23934 8916 23940 8968
rect 23992 8916 23998 8968
rect 27249 8959 27307 8965
rect 27249 8925 27261 8959
rect 27295 8925 27307 8959
rect 27249 8919 27307 8925
rect 20487 8860 21404 8888
rect 20487 8857 20499 8860
rect 20441 8851 20499 8857
rect 21542 8848 21548 8900
rect 21600 8848 21606 8900
rect 21726 8848 21732 8900
rect 21784 8848 21790 8900
rect 21818 8848 21824 8900
rect 21876 8888 21882 8900
rect 21929 8891 21987 8897
rect 21929 8888 21941 8891
rect 21876 8860 21941 8888
rect 21876 8848 21882 8860
rect 21929 8857 21941 8860
rect 21975 8857 21987 8891
rect 27264 8888 27292 8919
rect 27614 8916 27620 8968
rect 27672 8916 27678 8968
rect 27893 8959 27951 8965
rect 27893 8925 27905 8959
rect 27939 8956 27951 8959
rect 27985 8959 28043 8965
rect 27985 8956 27997 8959
rect 27939 8928 27997 8956
rect 27939 8925 27951 8928
rect 27893 8919 27951 8925
rect 27985 8925 27997 8928
rect 28031 8956 28043 8959
rect 28626 8956 28632 8968
rect 28031 8928 28632 8956
rect 28031 8925 28043 8928
rect 27985 8919 28043 8925
rect 28626 8916 28632 8928
rect 28684 8916 28690 8968
rect 31754 8916 31760 8968
rect 31812 8956 31818 8968
rect 32033 8959 32091 8965
rect 32033 8956 32045 8959
rect 31812 8928 32045 8956
rect 31812 8916 31818 8928
rect 32033 8925 32045 8928
rect 32079 8925 32091 8959
rect 32033 8919 32091 8925
rect 32306 8916 32312 8968
rect 32364 8916 32370 8968
rect 32490 8916 32496 8968
rect 32548 8956 32554 8968
rect 32677 8959 32735 8965
rect 32677 8956 32689 8959
rect 32548 8928 32689 8956
rect 32548 8916 32554 8928
rect 32677 8925 32689 8928
rect 32723 8925 32735 8959
rect 35728 8942 35756 8996
rect 36722 8984 36728 8996
rect 36780 8984 36786 9036
rect 36814 8984 36820 9036
rect 36872 8984 36878 9036
rect 39669 9027 39727 9033
rect 39669 9024 39681 9027
rect 37108 8996 39681 9024
rect 37108 8968 37136 8996
rect 39669 8993 39681 8996
rect 39715 9024 39727 9027
rect 40034 9024 40040 9036
rect 39715 8996 40040 9024
rect 39715 8993 39727 8996
rect 39669 8987 39727 8993
rect 40034 8984 40040 8996
rect 40092 8984 40098 9036
rect 32677 8919 32735 8925
rect 37090 8916 37096 8968
rect 37148 8916 37154 8968
rect 37185 8959 37243 8965
rect 37185 8925 37197 8959
rect 37231 8925 37243 8959
rect 37185 8919 37243 8925
rect 37369 8959 37427 8965
rect 37369 8925 37381 8959
rect 37415 8956 37427 8959
rect 37415 8928 37964 8956
rect 37415 8925 37427 8928
rect 37369 8919 37427 8925
rect 27798 8888 27804 8900
rect 27264 8860 27804 8888
rect 21929 8851 21987 8857
rect 27798 8848 27804 8860
rect 27856 8848 27862 8900
rect 36538 8848 36544 8900
rect 36596 8888 36602 8900
rect 37200 8888 37228 8919
rect 36596 8860 37228 8888
rect 36596 8848 36602 8860
rect 18049 8823 18107 8829
rect 18049 8789 18061 8823
rect 18095 8820 18107 8823
rect 18138 8820 18144 8832
rect 18095 8792 18144 8820
rect 18095 8789 18107 8792
rect 18049 8783 18107 8789
rect 18138 8780 18144 8792
rect 18196 8780 18202 8832
rect 20714 8780 20720 8832
rect 20772 8780 20778 8832
rect 21082 8780 21088 8832
rect 21140 8820 21146 8832
rect 21177 8823 21235 8829
rect 21177 8820 21189 8823
rect 21140 8792 21189 8820
rect 21140 8780 21146 8792
rect 21177 8789 21189 8792
rect 21223 8789 21235 8823
rect 21177 8783 21235 8789
rect 21358 8780 21364 8832
rect 21416 8820 21422 8832
rect 21744 8820 21772 8848
rect 21416 8792 21772 8820
rect 21416 8780 21422 8792
rect 27338 8780 27344 8832
rect 27396 8820 27402 8832
rect 27433 8823 27491 8829
rect 27433 8820 27445 8823
rect 27396 8792 27445 8820
rect 27396 8780 27402 8792
rect 27433 8789 27445 8792
rect 27479 8789 27491 8823
rect 27433 8783 27491 8789
rect 32493 8823 32551 8829
rect 32493 8789 32505 8823
rect 32539 8820 32551 8823
rect 32950 8820 32956 8832
rect 32539 8792 32956 8820
rect 32539 8789 32551 8792
rect 32493 8783 32551 8789
rect 32950 8780 32956 8792
rect 33008 8780 33014 8832
rect 35345 8823 35403 8829
rect 35345 8789 35357 8823
rect 35391 8820 35403 8823
rect 35986 8820 35992 8832
rect 35391 8792 35992 8820
rect 35391 8789 35403 8792
rect 35345 8783 35403 8789
rect 35986 8780 35992 8792
rect 36044 8780 36050 8832
rect 36722 8780 36728 8832
rect 36780 8820 36786 8832
rect 37936 8829 37964 8928
rect 38010 8848 38016 8900
rect 38068 8888 38074 8900
rect 38068 8860 38226 8888
rect 38068 8848 38074 8860
rect 39390 8848 39396 8900
rect 39448 8848 39454 8900
rect 37277 8823 37335 8829
rect 37277 8820 37289 8823
rect 36780 8792 37289 8820
rect 36780 8780 36786 8792
rect 37277 8789 37289 8792
rect 37323 8789 37335 8823
rect 37277 8783 37335 8789
rect 37921 8823 37979 8829
rect 37921 8789 37933 8823
rect 37967 8789 37979 8823
rect 37921 8783 37979 8789
rect 1104 8730 58880 8752
rect 1104 8678 4874 8730
rect 4926 8678 4938 8730
rect 4990 8678 5002 8730
rect 5054 8678 5066 8730
rect 5118 8678 5130 8730
rect 5182 8678 35594 8730
rect 35646 8678 35658 8730
rect 35710 8678 35722 8730
rect 35774 8678 35786 8730
rect 35838 8678 35850 8730
rect 35902 8678 58880 8730
rect 1104 8656 58880 8678
rect 18322 8616 18328 8628
rect 15580 8588 18328 8616
rect 15286 8440 15292 8492
rect 15344 8480 15350 8492
rect 15580 8489 15608 8588
rect 18322 8576 18328 8588
rect 18380 8576 18386 8628
rect 21174 8576 21180 8628
rect 21232 8576 21238 8628
rect 23017 8619 23075 8625
rect 23017 8616 23029 8619
rect 22066 8588 23029 8616
rect 17678 8508 17684 8560
rect 17736 8508 17742 8560
rect 21726 8548 21732 8560
rect 21008 8520 21732 8548
rect 15565 8483 15623 8489
rect 15565 8480 15577 8483
rect 15344 8452 15577 8480
rect 15344 8440 15350 8452
rect 15565 8449 15577 8452
rect 15611 8449 15623 8483
rect 15565 8443 15623 8449
rect 15749 8483 15807 8489
rect 15749 8449 15761 8483
rect 15795 8449 15807 8483
rect 15749 8443 15807 8449
rect 15764 8412 15792 8443
rect 15838 8440 15844 8492
rect 15896 8440 15902 8492
rect 16022 8440 16028 8492
rect 16080 8440 16086 8492
rect 18414 8440 18420 8492
rect 18472 8480 18478 8492
rect 19153 8483 19211 8489
rect 19153 8480 19165 8483
rect 18472 8452 19165 8480
rect 18472 8440 18478 8452
rect 19153 8449 19165 8452
rect 19199 8449 19211 8483
rect 20714 8480 20720 8492
rect 20562 8452 20720 8480
rect 19153 8443 19211 8449
rect 20714 8440 20720 8452
rect 20772 8480 20778 8492
rect 21008 8489 21036 8520
rect 21726 8508 21732 8520
rect 21784 8508 21790 8560
rect 20993 8483 21051 8489
rect 20772 8452 20852 8480
rect 20772 8440 20778 8452
rect 15930 8412 15936 8424
rect 15764 8384 15936 8412
rect 15930 8372 15936 8384
rect 15988 8372 15994 8424
rect 16666 8372 16672 8424
rect 16724 8372 16730 8424
rect 18046 8372 18052 8424
rect 18104 8412 18110 8424
rect 18141 8415 18199 8421
rect 18141 8412 18153 8415
rect 18104 8384 18153 8412
rect 18104 8372 18110 8384
rect 18141 8381 18153 8384
rect 18187 8381 18199 8415
rect 18141 8375 18199 8381
rect 19426 8372 19432 8424
rect 19484 8372 19490 8424
rect 20824 8344 20852 8452
rect 20993 8449 21005 8483
rect 21039 8449 21051 8483
rect 20993 8443 21051 8449
rect 21361 8483 21419 8489
rect 21361 8449 21373 8483
rect 21407 8480 21419 8483
rect 21542 8480 21548 8492
rect 21407 8452 21548 8480
rect 21407 8449 21419 8452
rect 21361 8443 21419 8449
rect 20901 8415 20959 8421
rect 20901 8381 20913 8415
rect 20947 8412 20959 8415
rect 21376 8412 21404 8443
rect 21542 8440 21548 8452
rect 21600 8440 21606 8492
rect 21637 8483 21695 8489
rect 21637 8449 21649 8483
rect 21683 8480 21695 8483
rect 22066 8480 22094 8588
rect 23017 8585 23029 8588
rect 23063 8616 23075 8619
rect 23474 8616 23480 8628
rect 23063 8588 23480 8616
rect 23063 8585 23075 8588
rect 23017 8579 23075 8585
rect 23474 8576 23480 8588
rect 23532 8576 23538 8628
rect 28994 8576 29000 8628
rect 29052 8576 29058 8628
rect 31478 8576 31484 8628
rect 31536 8576 31542 8628
rect 32582 8576 32588 8628
rect 32640 8616 32646 8628
rect 32953 8619 33011 8625
rect 32953 8616 32965 8619
rect 32640 8588 32965 8616
rect 32640 8576 32646 8588
rect 32953 8585 32965 8588
rect 32999 8585 33011 8619
rect 32953 8579 33011 8585
rect 37001 8619 37059 8625
rect 37001 8585 37013 8619
rect 37047 8616 37059 8619
rect 37274 8616 37280 8628
rect 37047 8588 37280 8616
rect 37047 8585 37059 8588
rect 37001 8579 37059 8585
rect 37274 8576 37280 8588
rect 37332 8576 37338 8628
rect 37645 8619 37703 8625
rect 37645 8585 37657 8619
rect 37691 8616 37703 8619
rect 37826 8616 37832 8628
rect 37691 8588 37832 8616
rect 37691 8585 37703 8588
rect 37645 8579 37703 8585
rect 37826 8576 37832 8588
rect 37884 8616 37890 8628
rect 38381 8619 38439 8625
rect 38381 8616 38393 8619
rect 37884 8588 38393 8616
rect 37884 8576 37890 8588
rect 38381 8585 38393 8588
rect 38427 8585 38439 8619
rect 41506 8616 41512 8628
rect 38381 8579 38439 8585
rect 39040 8588 41512 8616
rect 22922 8508 22928 8560
rect 22980 8548 22986 8560
rect 26602 8548 26608 8560
rect 22980 8520 23322 8548
rect 26542 8520 26608 8548
rect 22980 8508 22986 8520
rect 26602 8508 26608 8520
rect 26660 8508 26666 8560
rect 32306 8548 32312 8560
rect 31312 8520 32312 8548
rect 31312 8492 31340 8520
rect 32306 8508 32312 8520
rect 32364 8548 32370 8560
rect 32364 8520 32720 8548
rect 32364 8508 32370 8520
rect 21683 8452 22094 8480
rect 21683 8449 21695 8452
rect 21637 8443 21695 8449
rect 22462 8440 22468 8492
rect 22520 8440 22526 8492
rect 31294 8440 31300 8492
rect 31352 8440 31358 8492
rect 31665 8483 31723 8489
rect 31665 8449 31677 8483
rect 31711 8449 31723 8483
rect 31665 8443 31723 8449
rect 31941 8483 31999 8489
rect 31941 8449 31953 8483
rect 31987 8480 31999 8483
rect 32490 8480 32496 8492
rect 31987 8452 32496 8480
rect 31987 8449 31999 8452
rect 31941 8443 31999 8449
rect 20947 8384 21404 8412
rect 20947 8381 20959 8384
rect 20901 8375 20959 8381
rect 21818 8372 21824 8424
rect 21876 8412 21882 8424
rect 22373 8415 22431 8421
rect 22373 8412 22385 8415
rect 21876 8384 22385 8412
rect 21876 8372 21882 8384
rect 22373 8381 22385 8384
rect 22419 8381 22431 8415
rect 22373 8375 22431 8381
rect 22833 8415 22891 8421
rect 22833 8381 22845 8415
rect 22879 8412 22891 8415
rect 24489 8415 24547 8421
rect 24489 8412 24501 8415
rect 22879 8384 24501 8412
rect 22879 8381 22891 8384
rect 22833 8375 22891 8381
rect 24489 8381 24501 8384
rect 24535 8381 24547 8415
rect 24489 8375 24547 8381
rect 24765 8415 24823 8421
rect 24765 8381 24777 8415
rect 24811 8412 24823 8415
rect 25041 8415 25099 8421
rect 25041 8412 25053 8415
rect 24811 8384 25053 8412
rect 24811 8381 24823 8384
rect 24765 8375 24823 8381
rect 25041 8381 25053 8384
rect 25087 8381 25099 8415
rect 25041 8375 25099 8381
rect 22922 8344 22928 8356
rect 20824 8316 22928 8344
rect 22922 8304 22928 8316
rect 22980 8304 22986 8356
rect 16025 8279 16083 8285
rect 16025 8245 16037 8279
rect 16071 8276 16083 8279
rect 16114 8276 16120 8288
rect 16071 8248 16120 8276
rect 16071 8245 16083 8248
rect 16025 8239 16083 8245
rect 16114 8236 16120 8248
rect 16172 8236 16178 8288
rect 21358 8236 21364 8288
rect 21416 8236 21422 8288
rect 23934 8236 23940 8288
rect 23992 8276 23998 8288
rect 24780 8276 24808 8375
rect 25314 8372 25320 8424
rect 25372 8372 25378 8424
rect 26789 8415 26847 8421
rect 26789 8381 26801 8415
rect 26835 8412 26847 8415
rect 27062 8412 27068 8424
rect 26835 8384 27068 8412
rect 26835 8381 26847 8384
rect 26789 8375 26847 8381
rect 27062 8372 27068 8384
rect 27120 8412 27126 8424
rect 27525 8415 27583 8421
rect 27525 8412 27537 8415
rect 27120 8384 27537 8412
rect 27120 8372 27126 8384
rect 27525 8381 27537 8384
rect 27571 8381 27583 8415
rect 27525 8375 27583 8381
rect 27614 8372 27620 8424
rect 27672 8412 27678 8424
rect 28169 8415 28227 8421
rect 28169 8412 28181 8415
rect 27672 8384 28181 8412
rect 27672 8372 27678 8384
rect 28169 8381 28181 8384
rect 28215 8412 28227 8415
rect 28534 8412 28540 8424
rect 28215 8384 28540 8412
rect 28215 8381 28227 8384
rect 28169 8375 28227 8381
rect 28534 8372 28540 8384
rect 28592 8372 28598 8424
rect 28721 8415 28779 8421
rect 28721 8381 28733 8415
rect 28767 8381 28779 8415
rect 31680 8412 31708 8443
rect 32490 8440 32496 8452
rect 32548 8440 32554 8492
rect 32214 8412 32220 8424
rect 31680 8384 32220 8412
rect 28721 8375 28779 8381
rect 28074 8304 28080 8356
rect 28132 8344 28138 8356
rect 28736 8344 28764 8375
rect 32214 8372 32220 8384
rect 32272 8412 32278 8424
rect 32692 8421 32720 8520
rect 36078 8508 36084 8560
rect 36136 8508 36142 8560
rect 36173 8551 36231 8557
rect 36173 8517 36185 8551
rect 36219 8548 36231 8551
rect 36219 8520 36676 8548
rect 36219 8517 36231 8520
rect 36173 8511 36231 8517
rect 36648 8492 36676 8520
rect 36832 8520 37872 8548
rect 35529 8483 35587 8489
rect 35529 8449 35541 8483
rect 35575 8480 35587 8483
rect 35802 8480 35808 8492
rect 35575 8452 35808 8480
rect 35575 8449 35587 8452
rect 35529 8443 35587 8449
rect 35802 8440 35808 8452
rect 35860 8440 35866 8492
rect 35986 8440 35992 8492
rect 36044 8480 36050 8492
rect 36265 8483 36323 8489
rect 36265 8480 36277 8483
rect 36044 8452 36277 8480
rect 36044 8440 36050 8452
rect 36265 8449 36277 8452
rect 36311 8449 36323 8483
rect 36265 8443 36323 8449
rect 32677 8415 32735 8421
rect 32272 8384 32628 8412
rect 32272 8372 32278 8384
rect 28132 8316 28764 8344
rect 32125 8347 32183 8353
rect 28132 8304 28138 8316
rect 32125 8313 32137 8347
rect 32171 8313 32183 8347
rect 32125 8307 32183 8313
rect 23992 8248 24808 8276
rect 23992 8236 23998 8248
rect 26970 8236 26976 8288
rect 27028 8236 27034 8288
rect 28442 8236 28448 8288
rect 28500 8276 28506 8288
rect 28537 8279 28595 8285
rect 28537 8276 28549 8279
rect 28500 8248 28549 8276
rect 28500 8236 28506 8248
rect 28537 8245 28549 8248
rect 28583 8245 28595 8279
rect 28537 8239 28595 8245
rect 28626 8236 28632 8288
rect 28684 8236 28690 8288
rect 31754 8236 31760 8288
rect 31812 8276 31818 8288
rect 32140 8276 32168 8307
rect 31812 8248 32168 8276
rect 31812 8236 31818 8248
rect 32490 8236 32496 8288
rect 32548 8236 32554 8288
rect 32600 8285 32628 8384
rect 32677 8381 32689 8415
rect 32723 8381 32735 8415
rect 36280 8412 36308 8443
rect 36630 8440 36636 8492
rect 36688 8440 36694 8492
rect 36722 8440 36728 8492
rect 36780 8440 36786 8492
rect 36832 8412 36860 8520
rect 37366 8440 37372 8492
rect 37424 8440 37430 8492
rect 37844 8489 37872 8520
rect 38010 8508 38016 8560
rect 38068 8548 38074 8560
rect 39040 8548 39068 8588
rect 41506 8576 41512 8588
rect 41564 8576 41570 8628
rect 38068 8520 39146 8548
rect 38068 8508 38074 8520
rect 40034 8508 40040 8560
rect 40092 8548 40098 8560
rect 40092 8520 40632 8548
rect 40092 8508 40098 8520
rect 40604 8489 40632 8520
rect 37829 8483 37887 8489
rect 37829 8449 37841 8483
rect 37875 8449 37887 8483
rect 37829 8443 37887 8449
rect 38289 8483 38347 8489
rect 38289 8449 38301 8483
rect 38335 8449 38347 8483
rect 38289 8443 38347 8449
rect 40589 8483 40647 8489
rect 40589 8449 40601 8483
rect 40635 8449 40647 8483
rect 40589 8443 40647 8449
rect 36280 8384 36860 8412
rect 32677 8375 32735 8381
rect 36906 8372 36912 8424
rect 36964 8412 36970 8424
rect 38304 8412 38332 8443
rect 38841 8415 38899 8421
rect 38841 8412 38853 8415
rect 36964 8384 38853 8412
rect 36964 8372 36970 8384
rect 38841 8381 38853 8384
rect 38887 8381 38899 8415
rect 38841 8375 38899 8381
rect 40310 8372 40316 8424
rect 40368 8372 40374 8424
rect 36354 8304 36360 8356
rect 36412 8344 36418 8356
rect 36449 8347 36507 8353
rect 36449 8344 36461 8347
rect 36412 8316 36461 8344
rect 36412 8304 36418 8316
rect 36449 8313 36461 8316
rect 36495 8344 36507 8347
rect 38197 8347 38255 8353
rect 38197 8344 38209 8347
rect 36495 8316 38209 8344
rect 36495 8313 36507 8316
rect 36449 8307 36507 8313
rect 38197 8313 38209 8316
rect 38243 8313 38255 8347
rect 38197 8307 38255 8313
rect 32585 8279 32643 8285
rect 32585 8245 32597 8279
rect 32631 8276 32643 8279
rect 32674 8276 32680 8288
rect 32631 8248 32680 8276
rect 32631 8245 32643 8248
rect 32585 8239 32643 8245
rect 32674 8236 32680 8248
rect 32732 8236 32738 8288
rect 36262 8236 36268 8288
rect 36320 8276 36326 8288
rect 36541 8279 36599 8285
rect 36541 8276 36553 8279
rect 36320 8248 36553 8276
rect 36320 8236 36326 8248
rect 36541 8245 36553 8248
rect 36587 8245 36599 8279
rect 36541 8239 36599 8245
rect 37550 8236 37556 8288
rect 37608 8276 37614 8288
rect 37921 8279 37979 8285
rect 37921 8276 37933 8279
rect 37608 8248 37933 8276
rect 37608 8236 37614 8248
rect 37921 8245 37933 8248
rect 37967 8245 37979 8279
rect 37921 8239 37979 8245
rect 1104 8186 58880 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 58880 8186
rect 1104 8112 58880 8134
rect 16022 8032 16028 8084
rect 16080 8072 16086 8084
rect 16117 8075 16175 8081
rect 16117 8072 16129 8075
rect 16080 8044 16129 8072
rect 16080 8032 16086 8044
rect 16117 8041 16129 8044
rect 16163 8041 16175 8075
rect 16117 8035 16175 8041
rect 12066 7896 12072 7948
rect 12124 7936 12130 7948
rect 12161 7939 12219 7945
rect 12161 7936 12173 7939
rect 12124 7908 12173 7936
rect 12124 7896 12130 7908
rect 12161 7905 12173 7908
rect 12207 7936 12219 7939
rect 12434 7936 12440 7948
rect 12207 7908 12440 7936
rect 12207 7905 12219 7908
rect 12161 7899 12219 7905
rect 12434 7896 12440 7908
rect 12492 7936 12498 7948
rect 14093 7939 14151 7945
rect 14093 7936 14105 7939
rect 12492 7908 14105 7936
rect 12492 7896 12498 7908
rect 14093 7905 14105 7908
rect 14139 7936 14151 7939
rect 15378 7936 15384 7948
rect 14139 7908 15384 7936
rect 14139 7905 14151 7908
rect 14093 7899 14151 7905
rect 15378 7896 15384 7908
rect 15436 7896 15442 7948
rect 15841 7939 15899 7945
rect 15841 7905 15853 7939
rect 15887 7936 15899 7939
rect 16132 7936 16160 8035
rect 19426 8032 19432 8084
rect 19484 8072 19490 8084
rect 19797 8075 19855 8081
rect 19797 8072 19809 8075
rect 19484 8044 19809 8072
rect 19484 8032 19490 8044
rect 19797 8041 19809 8044
rect 19843 8041 19855 8075
rect 19797 8035 19855 8041
rect 21726 8032 21732 8084
rect 21784 8032 21790 8084
rect 21818 8032 21824 8084
rect 21876 8072 21882 8084
rect 21913 8075 21971 8081
rect 21913 8072 21925 8075
rect 21876 8044 21925 8072
rect 21876 8032 21882 8044
rect 21913 8041 21925 8044
rect 21959 8041 21971 8075
rect 21913 8035 21971 8041
rect 25314 8032 25320 8084
rect 25372 8072 25378 8084
rect 26053 8075 26111 8081
rect 26053 8072 26065 8075
rect 25372 8044 26065 8072
rect 25372 8032 25378 8044
rect 26053 8041 26065 8044
rect 26099 8041 26111 8075
rect 26053 8035 26111 8041
rect 28537 8075 28595 8081
rect 28537 8041 28549 8075
rect 28583 8072 28595 8075
rect 28626 8072 28632 8084
rect 28583 8044 28632 8072
rect 28583 8041 28595 8044
rect 28537 8035 28595 8041
rect 28626 8032 28632 8044
rect 28684 8032 28690 8084
rect 28905 8075 28963 8081
rect 28905 8041 28917 8075
rect 28951 8072 28963 8075
rect 29086 8072 29092 8084
rect 28951 8044 29092 8072
rect 28951 8041 28963 8044
rect 28905 8035 28963 8041
rect 29086 8032 29092 8044
rect 29144 8032 29150 8084
rect 32122 8032 32128 8084
rect 32180 8032 32186 8084
rect 37826 8032 37832 8084
rect 37884 8032 37890 8084
rect 38841 8075 38899 8081
rect 38841 8041 38853 8075
rect 38887 8072 38899 8075
rect 40310 8072 40316 8084
rect 38887 8044 40316 8072
rect 38887 8041 38899 8044
rect 38841 8035 38899 8041
rect 40310 8032 40316 8044
rect 40368 8032 40374 8084
rect 40957 8075 41015 8081
rect 40957 8041 40969 8075
rect 41003 8072 41015 8075
rect 41046 8072 41052 8084
rect 41003 8044 41052 8072
rect 41003 8041 41015 8044
rect 40957 8035 41015 8041
rect 16206 7964 16212 8016
rect 16264 8004 16270 8016
rect 16301 8007 16359 8013
rect 16301 8004 16313 8007
rect 16264 7976 16313 8004
rect 16264 7964 16270 7976
rect 16301 7973 16313 7976
rect 16347 8004 16359 8007
rect 27525 8007 27583 8013
rect 27525 8004 27537 8007
rect 16347 7976 18000 8004
rect 16347 7973 16359 7976
rect 16301 7967 16359 7973
rect 16482 7936 16488 7948
rect 15887 7908 16488 7936
rect 15887 7905 15899 7908
rect 15841 7899 15899 7905
rect 16482 7896 16488 7908
rect 16540 7896 16546 7948
rect 17678 7936 17684 7948
rect 16592 7908 17684 7936
rect 15470 7828 15476 7880
rect 15528 7868 15534 7880
rect 16592 7868 16620 7908
rect 17678 7896 17684 7908
rect 17736 7896 17742 7948
rect 15528 7840 16620 7868
rect 15528 7828 15534 7840
rect 16666 7828 16672 7880
rect 16724 7828 16730 7880
rect 16850 7828 16856 7880
rect 16908 7828 16914 7880
rect 17218 7828 17224 7880
rect 17276 7828 17282 7880
rect 17972 7877 18000 7976
rect 26804 7976 27537 8004
rect 26804 7948 26832 7976
rect 27525 7973 27537 7976
rect 27571 7973 27583 8007
rect 27525 7967 27583 7973
rect 27798 7964 27804 8016
rect 27856 8004 27862 8016
rect 28442 8004 28448 8016
rect 27856 7976 28448 8004
rect 27856 7964 27862 7976
rect 28442 7964 28448 7976
rect 28500 7964 28506 8016
rect 31754 7964 31760 8016
rect 31812 8004 31818 8016
rect 32309 8007 32367 8013
rect 32309 8004 32321 8007
rect 31812 7976 32321 8004
rect 31812 7964 31818 7976
rect 32309 7973 32321 7976
rect 32355 7973 32367 8007
rect 32309 7967 32367 7973
rect 32401 8007 32459 8013
rect 32401 7973 32413 8007
rect 32447 8004 32459 8007
rect 32490 8004 32496 8016
rect 32447 7976 32496 8004
rect 32447 7973 32459 7976
rect 32401 7967 32459 7973
rect 32490 7964 32496 7976
rect 32548 8004 32554 8016
rect 33778 8004 33784 8016
rect 32548 7976 33784 8004
rect 32548 7964 32554 7976
rect 33778 7964 33784 7976
rect 33836 7964 33842 8016
rect 36262 7964 36268 8016
rect 36320 8004 36326 8016
rect 36725 8007 36783 8013
rect 36725 8004 36737 8007
rect 36320 7976 36737 8004
rect 36320 7964 36326 7976
rect 36725 7973 36737 7976
rect 36771 7973 36783 8007
rect 37844 8004 37872 8032
rect 36725 7967 36783 7973
rect 36832 7976 37872 8004
rect 20257 7939 20315 7945
rect 20257 7905 20269 7939
rect 20303 7936 20315 7939
rect 21082 7936 21088 7948
rect 20303 7908 21088 7936
rect 20303 7905 20315 7908
rect 20257 7899 20315 7905
rect 21082 7896 21088 7908
rect 21140 7896 21146 7948
rect 21269 7939 21327 7945
rect 21269 7905 21281 7939
rect 21315 7936 21327 7939
rect 21542 7936 21548 7948
rect 21315 7908 21548 7936
rect 21315 7905 21327 7908
rect 21269 7899 21327 7905
rect 21542 7896 21548 7908
rect 21600 7896 21606 7948
rect 26697 7939 26755 7945
rect 26697 7905 26709 7939
rect 26743 7936 26755 7939
rect 26786 7936 26792 7948
rect 26743 7908 26792 7936
rect 26743 7905 26755 7908
rect 26697 7899 26755 7905
rect 26786 7896 26792 7908
rect 26844 7896 26850 7948
rect 27157 7939 27215 7945
rect 27157 7905 27169 7939
rect 27203 7905 27215 7939
rect 27157 7899 27215 7905
rect 17865 7871 17923 7877
rect 17865 7837 17877 7871
rect 17911 7837 17923 7871
rect 17865 7831 17923 7837
rect 17957 7871 18015 7877
rect 17957 7837 17969 7871
rect 18003 7837 18015 7871
rect 17957 7831 18015 7837
rect 12434 7760 12440 7812
rect 12492 7760 12498 7812
rect 13722 7800 13728 7812
rect 13662 7772 13728 7800
rect 13722 7760 13728 7772
rect 13780 7760 13786 7812
rect 14366 7760 14372 7812
rect 14424 7760 14430 7812
rect 15933 7803 15991 7809
rect 15933 7769 15945 7803
rect 15979 7769 15991 7803
rect 17880 7800 17908 7831
rect 18138 7828 18144 7880
rect 18196 7828 18202 7880
rect 20165 7871 20223 7877
rect 20165 7837 20177 7871
rect 20211 7868 20223 7871
rect 20625 7871 20683 7877
rect 20625 7868 20637 7871
rect 20211 7840 20637 7868
rect 20211 7837 20223 7840
rect 20165 7831 20223 7837
rect 20625 7837 20637 7840
rect 20671 7837 20683 7871
rect 20625 7831 20683 7837
rect 21174 7800 21180 7812
rect 17880 7772 21180 7800
rect 15933 7763 15991 7769
rect 13909 7735 13967 7741
rect 13909 7701 13921 7735
rect 13955 7732 13967 7735
rect 13998 7732 14004 7744
rect 13955 7704 14004 7732
rect 13955 7701 13967 7704
rect 13909 7695 13967 7701
rect 13998 7692 14004 7704
rect 14056 7732 14062 7744
rect 15838 7732 15844 7744
rect 14056 7704 15844 7732
rect 14056 7692 14062 7704
rect 15838 7692 15844 7704
rect 15896 7732 15902 7744
rect 15948 7732 15976 7763
rect 21174 7760 21180 7772
rect 21232 7760 21238 7812
rect 21560 7809 21588 7896
rect 26421 7871 26479 7877
rect 26421 7837 26433 7871
rect 26467 7868 26479 7871
rect 26970 7868 26976 7880
rect 26467 7840 26976 7868
rect 26467 7837 26479 7840
rect 26421 7831 26479 7837
rect 26970 7828 26976 7840
rect 27028 7828 27034 7880
rect 27062 7828 27068 7880
rect 27120 7828 27126 7880
rect 27172 7868 27200 7899
rect 27338 7896 27344 7948
rect 27396 7936 27402 7948
rect 27433 7939 27491 7945
rect 27433 7936 27445 7939
rect 27396 7908 27445 7936
rect 27396 7896 27402 7908
rect 27433 7905 27445 7908
rect 27479 7905 27491 7939
rect 27433 7899 27491 7905
rect 28534 7896 28540 7948
rect 28592 7936 28598 7948
rect 28629 7939 28687 7945
rect 28629 7936 28641 7939
rect 28592 7908 28641 7936
rect 28592 7896 28598 7908
rect 28629 7905 28641 7908
rect 28675 7905 28687 7939
rect 28629 7899 28687 7905
rect 30834 7896 30840 7948
rect 30892 7936 30898 7948
rect 31294 7936 31300 7948
rect 30892 7908 31300 7936
rect 30892 7896 30898 7908
rect 31294 7896 31300 7908
rect 31352 7936 31358 7948
rect 32217 7939 32275 7945
rect 32217 7936 32229 7939
rect 31352 7908 32229 7936
rect 31352 7896 31358 7908
rect 32217 7905 32229 7908
rect 32263 7905 32275 7939
rect 32217 7899 32275 7905
rect 32953 7939 33011 7945
rect 32953 7905 32965 7939
rect 32999 7905 33011 7939
rect 32953 7899 33011 7905
rect 33413 7939 33471 7945
rect 33413 7905 33425 7939
rect 33459 7936 33471 7939
rect 34422 7936 34428 7948
rect 33459 7908 34428 7936
rect 33459 7905 33471 7908
rect 33413 7899 33471 7905
rect 28074 7868 28080 7880
rect 27172 7840 28080 7868
rect 21545 7803 21603 7809
rect 21545 7769 21557 7803
rect 21591 7769 21603 7803
rect 27172 7800 27200 7840
rect 28074 7828 28080 7840
rect 28132 7828 28138 7880
rect 28718 7828 28724 7880
rect 28776 7868 28782 7880
rect 29546 7868 29552 7880
rect 28776 7840 29552 7868
rect 28776 7828 28782 7840
rect 29546 7828 29552 7840
rect 29604 7828 29610 7880
rect 32674 7828 32680 7880
rect 32732 7868 32738 7880
rect 32769 7871 32827 7877
rect 32769 7868 32781 7871
rect 32732 7840 32781 7868
rect 32732 7828 32738 7840
rect 32769 7837 32781 7840
rect 32815 7868 32827 7871
rect 32968 7868 32996 7899
rect 34422 7896 34428 7908
rect 34480 7896 34486 7948
rect 34514 7896 34520 7948
rect 34572 7936 34578 7948
rect 35802 7936 35808 7948
rect 34572 7908 35808 7936
rect 34572 7896 34578 7908
rect 35802 7896 35808 7908
rect 35860 7936 35866 7948
rect 35860 7908 36584 7936
rect 35860 7896 35866 7908
rect 32815 7840 32996 7868
rect 33045 7871 33103 7877
rect 32815 7837 32827 7840
rect 32769 7831 32827 7837
rect 33045 7837 33057 7871
rect 33091 7868 33103 7871
rect 33870 7868 33876 7880
rect 33091 7840 33876 7868
rect 33091 7837 33103 7840
rect 33045 7831 33103 7837
rect 33870 7828 33876 7840
rect 33928 7828 33934 7880
rect 36354 7828 36360 7880
rect 36412 7828 36418 7880
rect 36556 7877 36584 7908
rect 36630 7896 36636 7948
rect 36688 7896 36694 7948
rect 36832 7936 36860 7976
rect 36740 7908 36860 7936
rect 36541 7871 36599 7877
rect 36541 7837 36553 7871
rect 36587 7868 36599 7871
rect 36740 7868 36768 7908
rect 36998 7896 37004 7948
rect 37056 7936 37062 7948
rect 37056 7908 38792 7936
rect 37056 7896 37062 7908
rect 36587 7840 36768 7868
rect 36817 7871 36875 7877
rect 36587 7837 36599 7840
rect 36541 7831 36599 7837
rect 36817 7837 36829 7871
rect 36863 7868 36875 7871
rect 37550 7868 37556 7880
rect 36863 7840 37556 7868
rect 36863 7837 36875 7840
rect 36817 7831 36875 7837
rect 37550 7828 37556 7840
rect 37608 7828 37614 7880
rect 37642 7828 37648 7880
rect 37700 7828 37706 7880
rect 38010 7828 38016 7880
rect 38068 7828 38074 7880
rect 38764 7877 38792 7908
rect 38749 7871 38807 7877
rect 38749 7837 38761 7871
rect 38795 7837 38807 7871
rect 38749 7831 38807 7837
rect 39485 7871 39543 7877
rect 39485 7837 39497 7871
rect 39531 7868 39543 7871
rect 40034 7868 40040 7880
rect 39531 7840 40040 7868
rect 39531 7837 39543 7840
rect 39485 7831 39543 7837
rect 40034 7828 40040 7840
rect 40092 7828 40098 7880
rect 40773 7871 40831 7877
rect 40773 7837 40785 7871
rect 40819 7868 40831 7871
rect 40972 7868 41000 8035
rect 41046 8032 41052 8044
rect 41104 8032 41110 8084
rect 40819 7840 41000 7868
rect 40819 7837 40831 7840
rect 40773 7831 40831 7837
rect 21545 7763 21603 7769
rect 26528 7772 27200 7800
rect 15896 7704 15976 7732
rect 15896 7692 15902 7704
rect 16022 7692 16028 7744
rect 16080 7732 16086 7744
rect 16133 7735 16191 7741
rect 16133 7732 16145 7735
rect 16080 7704 16145 7732
rect 16080 7692 16086 7704
rect 16133 7701 16145 7704
rect 16179 7701 16191 7735
rect 16133 7695 16191 7701
rect 16669 7735 16727 7741
rect 16669 7701 16681 7735
rect 16715 7732 16727 7735
rect 16942 7732 16948 7744
rect 16715 7704 16948 7732
rect 16715 7701 16727 7704
rect 16669 7695 16727 7701
rect 16942 7692 16948 7704
rect 17000 7692 17006 7744
rect 17586 7692 17592 7744
rect 17644 7732 17650 7744
rect 18049 7735 18107 7741
rect 18049 7732 18061 7735
rect 17644 7704 18061 7732
rect 17644 7692 17650 7704
rect 18049 7701 18061 7704
rect 18095 7701 18107 7735
rect 18049 7695 18107 7701
rect 21358 7692 21364 7744
rect 21416 7732 21422 7744
rect 21745 7735 21803 7741
rect 21745 7732 21757 7735
rect 21416 7704 21757 7732
rect 21416 7692 21422 7704
rect 21745 7701 21757 7704
rect 21791 7701 21803 7735
rect 21745 7695 21803 7701
rect 26142 7692 26148 7744
rect 26200 7732 26206 7744
rect 26528 7741 26556 7772
rect 29822 7760 29828 7812
rect 29880 7760 29886 7812
rect 30374 7760 30380 7812
rect 30432 7760 30438 7812
rect 26513 7735 26571 7741
rect 26513 7732 26525 7735
rect 26200 7704 26525 7732
rect 26200 7692 26206 7704
rect 26513 7701 26525 7704
rect 26559 7701 26571 7735
rect 26513 7695 26571 7701
rect 31294 7692 31300 7744
rect 31352 7692 31358 7744
rect 37093 7735 37151 7741
rect 37093 7701 37105 7735
rect 37139 7732 37151 7735
rect 37182 7732 37188 7744
rect 37139 7704 37188 7732
rect 37139 7701 37151 7704
rect 37093 7695 37151 7701
rect 37182 7692 37188 7704
rect 37240 7692 37246 7744
rect 38657 7735 38715 7741
rect 38657 7701 38669 7735
rect 38703 7732 38715 7735
rect 38746 7732 38752 7744
rect 38703 7704 38752 7732
rect 38703 7701 38715 7704
rect 38657 7695 38715 7701
rect 38746 7692 38752 7704
rect 38804 7692 38810 7744
rect 1104 7642 58880 7664
rect 1104 7590 4874 7642
rect 4926 7590 4938 7642
rect 4990 7590 5002 7642
rect 5054 7590 5066 7642
rect 5118 7590 5130 7642
rect 5182 7590 35594 7642
rect 35646 7590 35658 7642
rect 35710 7590 35722 7642
rect 35774 7590 35786 7642
rect 35838 7590 35850 7642
rect 35902 7590 58880 7642
rect 1104 7568 58880 7590
rect 14366 7488 14372 7540
rect 14424 7528 14430 7540
rect 16117 7531 16175 7537
rect 16117 7528 16129 7531
rect 14424 7500 16129 7528
rect 14424 7488 14430 7500
rect 16117 7497 16129 7500
rect 16163 7497 16175 7531
rect 16117 7491 16175 7497
rect 16666 7488 16672 7540
rect 16724 7528 16730 7540
rect 16853 7531 16911 7537
rect 16853 7528 16865 7531
rect 16724 7500 16865 7528
rect 16724 7488 16730 7500
rect 16853 7497 16865 7500
rect 16899 7497 16911 7531
rect 16853 7491 16911 7497
rect 17497 7531 17555 7537
rect 17497 7497 17509 7531
rect 17543 7528 17555 7531
rect 18046 7528 18052 7540
rect 17543 7500 18052 7528
rect 17543 7497 17555 7500
rect 17497 7491 17555 7497
rect 18046 7488 18052 7500
rect 18104 7488 18110 7540
rect 20165 7531 20223 7537
rect 20165 7497 20177 7531
rect 20211 7528 20223 7531
rect 21082 7528 21088 7540
rect 20211 7500 21088 7528
rect 20211 7497 20223 7500
rect 20165 7491 20223 7497
rect 21082 7488 21088 7500
rect 21140 7488 21146 7540
rect 23290 7528 23296 7540
rect 22020 7500 23296 7528
rect 15286 7420 15292 7472
rect 15344 7420 15350 7472
rect 16025 7463 16083 7469
rect 16025 7429 16037 7463
rect 16071 7460 16083 7463
rect 16574 7460 16580 7472
rect 16071 7432 16580 7460
rect 16071 7429 16083 7432
rect 16025 7423 16083 7429
rect 16574 7420 16580 7432
rect 16632 7460 16638 7472
rect 22020 7469 22048 7500
rect 23290 7488 23296 7500
rect 23348 7488 23354 7540
rect 27246 7488 27252 7540
rect 27304 7528 27310 7540
rect 28261 7531 28319 7537
rect 28261 7528 28273 7531
rect 27304 7500 28273 7528
rect 27304 7488 27310 7500
rect 28261 7497 28273 7500
rect 28307 7497 28319 7531
rect 30374 7528 30380 7540
rect 28261 7491 28319 7497
rect 29472 7500 30380 7528
rect 22005 7463 22063 7469
rect 22005 7460 22017 7463
rect 16632 7432 22017 7460
rect 16632 7420 16638 7432
rect 22005 7429 22017 7432
rect 22051 7429 22063 7463
rect 28445 7463 28503 7469
rect 28445 7460 28457 7463
rect 22005 7423 22063 7429
rect 27632 7432 28457 7460
rect 27632 7404 27660 7432
rect 28445 7429 28457 7432
rect 28491 7429 28503 7463
rect 28445 7423 28503 7429
rect 12805 7395 12863 7401
rect 12805 7361 12817 7395
rect 12851 7392 12863 7395
rect 13449 7395 13507 7401
rect 13449 7392 13461 7395
rect 12851 7364 13461 7392
rect 12851 7361 12863 7364
rect 12805 7355 12863 7361
rect 13449 7361 13461 7364
rect 13495 7361 13507 7395
rect 13449 7355 13507 7361
rect 13998 7352 14004 7404
rect 14056 7352 14062 7404
rect 16114 7352 16120 7404
rect 16172 7352 16178 7404
rect 16206 7352 16212 7404
rect 16264 7352 16270 7404
rect 16482 7352 16488 7404
rect 16540 7392 16546 7404
rect 16669 7395 16727 7401
rect 16669 7392 16681 7395
rect 16540 7364 16681 7392
rect 16540 7352 16546 7364
rect 16669 7361 16681 7364
rect 16715 7361 16727 7395
rect 16669 7355 16727 7361
rect 17037 7395 17095 7401
rect 17037 7361 17049 7395
rect 17083 7361 17095 7395
rect 17037 7355 17095 7361
rect 17313 7395 17371 7401
rect 17313 7361 17325 7395
rect 17359 7361 17371 7395
rect 17313 7355 17371 7361
rect 12434 7284 12440 7336
rect 12492 7284 12498 7336
rect 12894 7284 12900 7336
rect 12952 7284 12958 7336
rect 16393 7327 16451 7333
rect 16393 7293 16405 7327
rect 16439 7324 16451 7327
rect 16942 7324 16948 7336
rect 16439 7296 16948 7324
rect 16439 7293 16451 7296
rect 16393 7287 16451 7293
rect 16942 7284 16948 7296
rect 17000 7284 17006 7336
rect 15838 7216 15844 7268
rect 15896 7256 15902 7268
rect 17052 7256 17080 7355
rect 17328 7324 17356 7355
rect 17402 7352 17408 7404
rect 17460 7352 17466 7404
rect 17586 7352 17592 7404
rect 17644 7352 17650 7404
rect 20346 7352 20352 7404
rect 20404 7352 20410 7404
rect 20438 7352 20444 7404
rect 20496 7352 20502 7404
rect 20530 7352 20536 7404
rect 20588 7352 20594 7404
rect 21177 7395 21235 7401
rect 21177 7392 21189 7395
rect 20640 7364 21189 7392
rect 20254 7324 20260 7336
rect 17328 7296 20260 7324
rect 20254 7284 20260 7296
rect 20312 7284 20318 7336
rect 15896 7228 17080 7256
rect 15896 7216 15902 7228
rect 17126 7216 17132 7268
rect 17184 7256 17190 7268
rect 20640 7256 20668 7364
rect 21177 7361 21189 7364
rect 21223 7361 21235 7395
rect 21177 7355 21235 7361
rect 17184 7228 20668 7256
rect 17184 7216 17190 7228
rect 20714 7216 20720 7268
rect 20772 7216 20778 7268
rect 21192 7256 21220 7355
rect 21358 7352 21364 7404
rect 21416 7352 21422 7404
rect 23014 7352 23020 7404
rect 23072 7352 23078 7404
rect 23106 7352 23112 7404
rect 23164 7392 23170 7404
rect 23201 7395 23259 7401
rect 23201 7392 23213 7395
rect 23164 7364 23213 7392
rect 23164 7352 23170 7364
rect 23201 7361 23213 7364
rect 23247 7361 23259 7395
rect 23201 7355 23259 7361
rect 26329 7395 26387 7401
rect 26329 7361 26341 7395
rect 26375 7392 26387 7395
rect 26973 7395 27031 7401
rect 26973 7392 26985 7395
rect 26375 7364 26985 7392
rect 26375 7361 26387 7364
rect 26329 7355 26387 7361
rect 26973 7361 26985 7364
rect 27019 7361 27031 7395
rect 26973 7355 27031 7361
rect 27614 7352 27620 7404
rect 27672 7352 27678 7404
rect 28077 7395 28135 7401
rect 28077 7361 28089 7395
rect 28123 7361 28135 7395
rect 28077 7355 28135 7361
rect 22002 7284 22008 7336
rect 22060 7324 22066 7336
rect 22741 7327 22799 7333
rect 22741 7324 22753 7327
rect 22060 7296 22753 7324
rect 22060 7284 22066 7296
rect 22741 7293 22753 7296
rect 22787 7324 22799 7327
rect 23934 7324 23940 7336
rect 22787 7296 23940 7324
rect 22787 7293 22799 7296
rect 22741 7287 22799 7293
rect 23934 7284 23940 7296
rect 23992 7284 23998 7336
rect 26234 7284 26240 7336
rect 26292 7324 26298 7336
rect 26421 7327 26479 7333
rect 26421 7324 26433 7327
rect 26292 7296 26433 7324
rect 26292 7284 26298 7296
rect 26421 7293 26433 7296
rect 26467 7293 26479 7327
rect 26421 7287 26479 7293
rect 26513 7327 26571 7333
rect 26513 7293 26525 7327
rect 26559 7293 26571 7327
rect 26513 7287 26571 7293
rect 23106 7256 23112 7268
rect 21192 7228 23112 7256
rect 23106 7216 23112 7228
rect 23164 7216 23170 7268
rect 25869 7259 25927 7265
rect 25869 7225 25881 7259
rect 25915 7256 25927 7259
rect 26528 7256 26556 7287
rect 26602 7284 26608 7336
rect 26660 7324 26666 7336
rect 28092 7324 28120 7355
rect 28534 7352 28540 7404
rect 28592 7392 28598 7404
rect 28629 7395 28687 7401
rect 28629 7392 28641 7395
rect 28592 7364 28641 7392
rect 28592 7352 28598 7364
rect 28629 7361 28641 7364
rect 28675 7361 28687 7395
rect 28629 7355 28687 7361
rect 29472 7324 29500 7500
rect 30374 7488 30380 7500
rect 30432 7488 30438 7540
rect 31846 7488 31852 7540
rect 31904 7488 31910 7540
rect 33870 7488 33876 7540
rect 33928 7528 33934 7540
rect 35805 7531 35863 7537
rect 35805 7528 35817 7531
rect 33928 7500 34560 7528
rect 33928 7488 33934 7500
rect 29546 7420 29552 7472
rect 29604 7460 29610 7472
rect 31864 7460 31892 7488
rect 32858 7460 32864 7472
rect 29604 7432 31754 7460
rect 31864 7432 32864 7460
rect 29604 7420 29610 7432
rect 29917 7395 29975 7401
rect 29917 7361 29929 7395
rect 29963 7392 29975 7395
rect 30653 7395 30711 7401
rect 30653 7392 30665 7395
rect 29963 7364 30665 7392
rect 29963 7361 29975 7364
rect 29917 7355 29975 7361
rect 30653 7361 30665 7364
rect 30699 7361 30711 7395
rect 30653 7355 30711 7361
rect 31294 7352 31300 7404
rect 31352 7352 31358 7404
rect 31726 7392 31754 7432
rect 32858 7420 32864 7432
rect 32916 7420 32922 7472
rect 34532 7401 34560 7500
rect 35176 7500 35817 7528
rect 34790 7420 34796 7472
rect 34848 7460 34854 7472
rect 35176 7469 35204 7500
rect 35805 7497 35817 7500
rect 35851 7497 35863 7531
rect 35805 7491 35863 7497
rect 36265 7531 36323 7537
rect 36265 7497 36277 7531
rect 36311 7528 36323 7531
rect 36630 7528 36636 7540
rect 36311 7500 36636 7528
rect 36311 7497 36323 7500
rect 36265 7491 36323 7497
rect 36630 7488 36636 7500
rect 36688 7488 36694 7540
rect 37093 7531 37151 7537
rect 37093 7497 37105 7531
rect 37139 7528 37151 7531
rect 38010 7528 38016 7540
rect 37139 7500 38016 7528
rect 37139 7497 37151 7500
rect 37093 7491 37151 7497
rect 38010 7488 38016 7500
rect 38068 7488 38074 7540
rect 35161 7463 35219 7469
rect 35161 7460 35173 7463
rect 34848 7432 35173 7460
rect 34848 7420 34854 7432
rect 35161 7429 35173 7432
rect 35207 7429 35219 7463
rect 35161 7423 35219 7429
rect 35366 7463 35424 7469
rect 35366 7429 35378 7463
rect 35412 7460 35424 7463
rect 36817 7463 36875 7469
rect 35412 7432 35480 7460
rect 35412 7429 35424 7432
rect 35366 7423 35424 7429
rect 32125 7395 32183 7401
rect 32125 7392 32137 7395
rect 31726 7364 32137 7392
rect 32125 7361 32137 7364
rect 32171 7361 32183 7395
rect 32125 7355 32183 7361
rect 34517 7395 34575 7401
rect 34517 7361 34529 7395
rect 34563 7361 34575 7395
rect 34517 7355 34575 7361
rect 35452 7336 35480 7432
rect 36817 7429 36829 7463
rect 36863 7460 36875 7463
rect 37182 7460 37188 7472
rect 36863 7432 37188 7460
rect 36863 7429 36875 7432
rect 36817 7423 36875 7429
rect 37182 7420 37188 7432
rect 37240 7420 37246 7472
rect 37918 7420 37924 7472
rect 37976 7420 37982 7472
rect 35989 7395 36047 7401
rect 35989 7361 36001 7395
rect 36035 7392 36047 7395
rect 36035 7364 36492 7392
rect 36035 7361 36047 7364
rect 35989 7355 36047 7361
rect 26660 7296 29500 7324
rect 30009 7327 30067 7333
rect 26660 7284 26666 7296
rect 30009 7293 30021 7327
rect 30055 7293 30067 7327
rect 30009 7287 30067 7293
rect 30193 7327 30251 7333
rect 30193 7293 30205 7327
rect 30239 7324 30251 7327
rect 30239 7296 30788 7324
rect 30239 7293 30251 7296
rect 30193 7287 30251 7293
rect 26786 7256 26792 7268
rect 25915 7228 26792 7256
rect 25915 7225 25927 7228
rect 25869 7219 25927 7225
rect 26786 7216 26792 7228
rect 26844 7256 26850 7268
rect 29549 7259 29607 7265
rect 26844 7228 28994 7256
rect 26844 7216 26850 7228
rect 16758 7148 16764 7200
rect 16816 7188 16822 7200
rect 17037 7191 17095 7197
rect 17037 7188 17049 7191
rect 16816 7160 17049 7188
rect 16816 7148 16822 7160
rect 17037 7157 17049 7160
rect 17083 7157 17095 7191
rect 17037 7151 17095 7157
rect 21266 7148 21272 7200
rect 21324 7188 21330 7200
rect 21361 7191 21419 7197
rect 21361 7188 21373 7191
rect 21324 7160 21373 7188
rect 21324 7148 21330 7160
rect 21361 7157 21373 7160
rect 21407 7157 21419 7191
rect 21361 7151 21419 7157
rect 23017 7191 23075 7197
rect 23017 7157 23029 7191
rect 23063 7188 23075 7191
rect 23842 7188 23848 7200
rect 23063 7160 23848 7188
rect 23063 7157 23075 7160
rect 23017 7151 23075 7157
rect 23842 7148 23848 7160
rect 23900 7148 23906 7200
rect 25958 7148 25964 7200
rect 26016 7148 26022 7200
rect 27985 7191 28043 7197
rect 27985 7157 27997 7191
rect 28031 7188 28043 7191
rect 28166 7188 28172 7200
rect 28031 7160 28172 7188
rect 28031 7157 28043 7160
rect 27985 7151 28043 7157
rect 28166 7148 28172 7160
rect 28224 7148 28230 7200
rect 28966 7188 28994 7228
rect 29549 7225 29561 7259
rect 29595 7256 29607 7259
rect 29822 7256 29828 7268
rect 29595 7228 29828 7256
rect 29595 7225 29607 7228
rect 29549 7219 29607 7225
rect 29822 7216 29828 7228
rect 29880 7216 29886 7268
rect 30024 7256 30052 7287
rect 30650 7256 30656 7268
rect 30024 7228 30656 7256
rect 30650 7216 30656 7228
rect 30708 7216 30714 7268
rect 29270 7188 29276 7200
rect 28966 7160 29276 7188
rect 29270 7148 29276 7160
rect 29328 7188 29334 7200
rect 30469 7191 30527 7197
rect 30469 7188 30481 7191
rect 29328 7160 30481 7188
rect 29328 7148 29334 7160
rect 30469 7157 30481 7160
rect 30515 7188 30527 7191
rect 30760 7188 30788 7296
rect 32398 7284 32404 7336
rect 32456 7284 32462 7336
rect 35434 7284 35440 7336
rect 35492 7324 35498 7336
rect 35621 7327 35679 7333
rect 35621 7324 35633 7327
rect 35492 7296 35633 7324
rect 35492 7284 35498 7296
rect 35621 7293 35633 7296
rect 35667 7293 35679 7327
rect 35621 7287 35679 7293
rect 35713 7327 35771 7333
rect 35713 7293 35725 7327
rect 35759 7293 35771 7327
rect 35713 7287 35771 7293
rect 36081 7327 36139 7333
rect 36081 7293 36093 7327
rect 36127 7324 36139 7327
rect 36354 7324 36360 7336
rect 36127 7296 36360 7324
rect 36127 7293 36139 7296
rect 36081 7287 36139 7293
rect 35728 7256 35756 7287
rect 36354 7284 36360 7296
rect 36412 7284 36418 7336
rect 36464 7324 36492 7364
rect 36538 7352 36544 7404
rect 36596 7352 36602 7404
rect 36722 7352 36728 7404
rect 36780 7352 36786 7404
rect 36909 7395 36967 7401
rect 36909 7361 36921 7395
rect 36955 7392 36967 7395
rect 36998 7392 37004 7404
rect 36955 7364 37004 7392
rect 36955 7361 36967 7364
rect 36909 7355 36967 7361
rect 36998 7352 37004 7364
rect 37056 7352 37062 7404
rect 38746 7352 38752 7404
rect 38804 7352 38810 7404
rect 39117 7395 39175 7401
rect 39117 7361 39129 7395
rect 39163 7392 39175 7395
rect 40034 7392 40040 7404
rect 39163 7364 40040 7392
rect 39163 7361 39175 7364
rect 39117 7355 39175 7361
rect 40034 7352 40040 7364
rect 40092 7352 40098 7404
rect 37323 7327 37381 7333
rect 37323 7324 37335 7327
rect 36464 7296 37335 7324
rect 37323 7293 37335 7296
rect 37369 7324 37381 7327
rect 37642 7324 37648 7336
rect 37369 7296 37648 7324
rect 37369 7293 37381 7296
rect 37323 7287 37381 7293
rect 37642 7284 37648 7296
rect 37700 7284 37706 7336
rect 35360 7228 35756 7256
rect 36372 7256 36400 7284
rect 36998 7256 37004 7268
rect 36372 7228 37004 7256
rect 35360 7200 35388 7228
rect 36998 7216 37004 7228
rect 37056 7216 37062 7268
rect 31662 7188 31668 7200
rect 30515 7160 31668 7188
rect 30515 7157 30527 7160
rect 30469 7151 30527 7157
rect 31662 7148 31668 7160
rect 31720 7188 31726 7200
rect 32950 7188 32956 7200
rect 31720 7160 32956 7188
rect 31720 7148 31726 7160
rect 32950 7148 32956 7160
rect 33008 7148 33014 7200
rect 33134 7148 33140 7200
rect 33192 7188 33198 7200
rect 33965 7191 34023 7197
rect 33965 7188 33977 7191
rect 33192 7160 33977 7188
rect 33192 7148 33198 7160
rect 33965 7157 33977 7160
rect 34011 7157 34023 7191
rect 33965 7151 34023 7157
rect 35342 7148 35348 7200
rect 35400 7148 35406 7200
rect 35529 7191 35587 7197
rect 35529 7157 35541 7191
rect 35575 7188 35587 7191
rect 36170 7188 36176 7200
rect 35575 7160 36176 7188
rect 35575 7157 35587 7160
rect 35529 7151 35587 7157
rect 36170 7148 36176 7160
rect 36228 7148 36234 7200
rect 1104 7098 58880 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 58880 7098
rect 1104 7024 58880 7046
rect 23842 6944 23848 6996
rect 23900 6984 23906 6996
rect 23949 6987 24007 6993
rect 23949 6984 23961 6987
rect 23900 6956 23961 6984
rect 23900 6944 23906 6956
rect 23949 6953 23961 6956
rect 23995 6953 24007 6987
rect 23949 6947 24007 6953
rect 25488 6987 25546 6993
rect 25488 6953 25500 6987
rect 25534 6984 25546 6987
rect 25958 6984 25964 6996
rect 25534 6956 25964 6984
rect 25534 6953 25546 6956
rect 25488 6947 25546 6953
rect 25958 6944 25964 6956
rect 26016 6944 26022 6996
rect 26234 6944 26240 6996
rect 26292 6984 26298 6996
rect 28534 6984 28540 6996
rect 26292 6956 28540 6984
rect 26292 6944 26298 6956
rect 15838 6876 15844 6928
rect 15896 6916 15902 6928
rect 15933 6919 15991 6925
rect 15933 6916 15945 6919
rect 15896 6888 15945 6916
rect 15896 6876 15902 6888
rect 15933 6885 15945 6888
rect 15979 6885 15991 6919
rect 15933 6879 15991 6885
rect 27341 6919 27399 6925
rect 27341 6885 27353 6919
rect 27387 6916 27399 6919
rect 27387 6888 27568 6916
rect 27387 6885 27399 6888
rect 27341 6879 27399 6885
rect 16482 6848 16488 6860
rect 16132 6820 16488 6848
rect 14734 6740 14740 6792
rect 14792 6740 14798 6792
rect 16132 6789 16160 6820
rect 16482 6808 16488 6820
rect 16540 6808 16546 6860
rect 16574 6808 16580 6860
rect 16632 6808 16638 6860
rect 20349 6851 20407 6857
rect 20349 6848 20361 6851
rect 18340 6820 20361 6848
rect 16117 6783 16175 6789
rect 16117 6749 16129 6783
rect 16163 6749 16175 6783
rect 16117 6743 16175 6749
rect 16209 6783 16267 6789
rect 16209 6749 16221 6783
rect 16255 6780 16267 6783
rect 16758 6780 16764 6792
rect 16255 6752 16764 6780
rect 16255 6749 16267 6752
rect 16209 6743 16267 6749
rect 16758 6740 16764 6752
rect 16816 6740 16822 6792
rect 17678 6740 17684 6792
rect 17736 6780 17742 6792
rect 18340 6789 18368 6820
rect 20349 6817 20361 6820
rect 20395 6848 20407 6851
rect 20714 6848 20720 6860
rect 20395 6820 20720 6848
rect 20395 6817 20407 6820
rect 20349 6811 20407 6817
rect 20714 6808 20720 6820
rect 20772 6808 20778 6860
rect 20901 6851 20959 6857
rect 20901 6817 20913 6851
rect 20947 6848 20959 6851
rect 21269 6851 21327 6857
rect 21269 6848 21281 6851
rect 20947 6820 21281 6848
rect 20947 6817 20959 6820
rect 20901 6811 20959 6817
rect 21269 6817 21281 6820
rect 21315 6848 21327 6851
rect 21358 6848 21364 6860
rect 21315 6820 21364 6848
rect 21315 6817 21327 6820
rect 21269 6811 21327 6817
rect 21358 6808 21364 6820
rect 21416 6808 21422 6860
rect 22465 6851 22523 6857
rect 22465 6848 22477 6851
rect 21928 6820 22477 6848
rect 18325 6783 18383 6789
rect 18325 6780 18337 6783
rect 17736 6752 18337 6780
rect 17736 6740 17742 6752
rect 18325 6749 18337 6752
rect 18371 6749 18383 6783
rect 18325 6743 18383 6749
rect 20254 6740 20260 6792
rect 20312 6780 20318 6792
rect 20530 6780 20536 6792
rect 20312 6752 20536 6780
rect 20312 6740 20318 6752
rect 20530 6740 20536 6752
rect 20588 6740 20594 6792
rect 20806 6740 20812 6792
rect 20864 6780 20870 6792
rect 21177 6783 21235 6789
rect 21177 6780 21189 6783
rect 20864 6752 21189 6780
rect 20864 6740 20870 6752
rect 21177 6749 21189 6752
rect 21223 6780 21235 6783
rect 21726 6780 21732 6792
rect 21223 6752 21732 6780
rect 21223 6749 21235 6752
rect 21177 6743 21235 6749
rect 21726 6740 21732 6752
rect 21784 6780 21790 6792
rect 21928 6780 21956 6820
rect 22465 6817 22477 6820
rect 22511 6817 22523 6851
rect 22922 6848 22928 6860
rect 22465 6811 22523 6817
rect 22572 6820 22928 6848
rect 21784 6752 21956 6780
rect 21784 6740 21790 6752
rect 22002 6740 22008 6792
rect 22060 6740 22066 6792
rect 16485 6715 16543 6721
rect 16485 6681 16497 6715
rect 16531 6712 16543 6715
rect 17402 6712 17408 6724
rect 16531 6684 17408 6712
rect 16531 6681 16543 6684
rect 16485 6675 16543 6681
rect 17402 6672 17408 6684
rect 17460 6712 17466 6724
rect 18509 6715 18567 6721
rect 18509 6712 18521 6715
rect 17460 6684 18521 6712
rect 17460 6672 17466 6684
rect 18509 6681 18521 6684
rect 18555 6712 18567 6715
rect 20346 6712 20352 6724
rect 18555 6684 20352 6712
rect 18555 6681 18567 6684
rect 18509 6675 18567 6681
rect 20346 6672 20352 6684
rect 20404 6712 20410 6724
rect 20404 6684 20760 6712
rect 20404 6672 20410 6684
rect 14090 6604 14096 6656
rect 14148 6604 14154 6656
rect 14918 6604 14924 6656
rect 14976 6644 14982 6656
rect 16022 6644 16028 6656
rect 14976 6616 16028 6644
rect 14976 6604 14982 6616
rect 16022 6604 16028 6616
rect 16080 6644 16086 6656
rect 16301 6647 16359 6653
rect 16301 6644 16313 6647
rect 16080 6616 16313 6644
rect 16080 6604 16086 6616
rect 16301 6613 16313 6616
rect 16347 6613 16359 6647
rect 16301 6607 16359 6613
rect 18138 6604 18144 6656
rect 18196 6604 18202 6656
rect 20622 6604 20628 6656
rect 20680 6604 20686 6656
rect 20732 6653 20760 6684
rect 21910 6672 21916 6724
rect 21968 6712 21974 6724
rect 22572 6712 22600 6820
rect 22922 6808 22928 6820
rect 22980 6808 22986 6860
rect 23566 6808 23572 6860
rect 23624 6848 23630 6860
rect 24213 6851 24271 6857
rect 24213 6848 24225 6851
rect 23624 6820 24225 6848
rect 23624 6808 23630 6820
rect 24213 6817 24225 6820
rect 24259 6848 24271 6851
rect 25225 6851 25283 6857
rect 25225 6848 25237 6851
rect 24259 6820 25237 6848
rect 24259 6817 24271 6820
rect 24213 6811 24271 6817
rect 25225 6817 25237 6820
rect 25271 6817 25283 6851
rect 25225 6811 25283 6817
rect 27065 6783 27123 6789
rect 27065 6749 27077 6783
rect 27111 6780 27123 6783
rect 27246 6780 27252 6792
rect 27111 6752 27252 6780
rect 27111 6749 27123 6752
rect 27065 6743 27123 6749
rect 27246 6740 27252 6752
rect 27304 6740 27310 6792
rect 27338 6740 27344 6792
rect 27396 6740 27402 6792
rect 27430 6740 27436 6792
rect 27488 6740 27494 6792
rect 21968 6684 22600 6712
rect 21968 6672 21974 6684
rect 22922 6672 22928 6724
rect 22980 6672 22986 6724
rect 26050 6672 26056 6724
rect 26108 6672 26114 6724
rect 27448 6712 27476 6740
rect 26988 6684 27476 6712
rect 27540 6712 27568 6888
rect 27632 6789 27660 6956
rect 28534 6944 28540 6956
rect 28592 6944 28598 6996
rect 32309 6987 32367 6993
rect 32309 6953 32321 6987
rect 32355 6984 32367 6987
rect 32398 6984 32404 6996
rect 32355 6956 32404 6984
rect 32355 6953 32367 6956
rect 32309 6947 32367 6953
rect 32398 6944 32404 6956
rect 32456 6944 32462 6996
rect 32858 6944 32864 6996
rect 32916 6984 32922 6996
rect 34606 6984 34612 6996
rect 32916 6956 34612 6984
rect 32916 6944 32922 6956
rect 34606 6944 34612 6956
rect 34664 6944 34670 6996
rect 36538 6944 36544 6996
rect 36596 6944 36602 6996
rect 36722 6944 36728 6996
rect 36780 6984 36786 6996
rect 36817 6987 36875 6993
rect 36817 6984 36829 6987
rect 36780 6956 36829 6984
rect 36780 6944 36786 6956
rect 36817 6953 36829 6956
rect 36863 6953 36875 6987
rect 36817 6947 36875 6953
rect 33042 6876 33048 6928
rect 33100 6916 33106 6928
rect 33229 6919 33287 6925
rect 33229 6916 33241 6919
rect 33100 6888 33241 6916
rect 33100 6876 33106 6888
rect 33229 6885 33241 6888
rect 33275 6916 33287 6919
rect 34514 6916 34520 6928
rect 33275 6888 34520 6916
rect 33275 6885 33287 6888
rect 33229 6879 33287 6885
rect 34514 6876 34520 6888
rect 34572 6876 34578 6928
rect 30650 6808 30656 6860
rect 30708 6808 30714 6860
rect 32858 6808 32864 6860
rect 32916 6808 32922 6860
rect 34333 6851 34391 6857
rect 34333 6817 34345 6851
rect 34379 6848 34391 6851
rect 35342 6848 35348 6860
rect 34379 6820 35348 6848
rect 34379 6817 34391 6820
rect 34333 6811 34391 6817
rect 35342 6808 35348 6820
rect 35400 6808 35406 6860
rect 27617 6783 27675 6789
rect 27617 6749 27629 6783
rect 27663 6749 27675 6783
rect 27617 6743 27675 6749
rect 30745 6783 30803 6789
rect 30745 6749 30757 6783
rect 30791 6780 30803 6783
rect 31294 6780 31300 6792
rect 30791 6752 31300 6780
rect 30791 6749 30803 6752
rect 30745 6743 30803 6749
rect 31294 6740 31300 6752
rect 31352 6740 31358 6792
rect 32677 6783 32735 6789
rect 32677 6749 32689 6783
rect 32723 6780 32735 6783
rect 33134 6780 33140 6792
rect 32723 6752 33140 6780
rect 32723 6749 32735 6752
rect 32677 6743 32735 6749
rect 33134 6740 33140 6752
rect 33192 6740 33198 6792
rect 33962 6740 33968 6792
rect 34020 6780 34026 6792
rect 34241 6783 34299 6789
rect 34241 6780 34253 6783
rect 34020 6752 34253 6780
rect 34020 6740 34026 6752
rect 34241 6749 34253 6752
rect 34287 6749 34299 6783
rect 34241 6743 34299 6749
rect 34422 6740 34428 6792
rect 34480 6740 34486 6792
rect 35360 6780 35388 6808
rect 35621 6783 35679 6789
rect 35621 6780 35633 6783
rect 35360 6752 35633 6780
rect 35621 6749 35633 6752
rect 35667 6749 35679 6783
rect 35621 6743 35679 6749
rect 35713 6783 35771 6789
rect 35713 6749 35725 6783
rect 35759 6749 35771 6783
rect 35713 6743 35771 6749
rect 35434 6712 35440 6724
rect 27540 6684 35440 6712
rect 20717 6647 20775 6653
rect 20717 6613 20729 6647
rect 20763 6644 20775 6647
rect 20898 6644 20904 6656
rect 20763 6616 20904 6644
rect 20763 6613 20775 6616
rect 20717 6607 20775 6613
rect 20898 6604 20904 6616
rect 20956 6604 20962 6656
rect 21545 6647 21603 6653
rect 21545 6613 21557 6647
rect 21591 6644 21603 6647
rect 23014 6644 23020 6656
rect 21591 6616 23020 6644
rect 21591 6613 21603 6616
rect 21545 6607 21603 6613
rect 23014 6604 23020 6616
rect 23072 6604 23078 6656
rect 26988 6653 27016 6684
rect 35434 6672 35440 6684
rect 35492 6672 35498 6724
rect 35728 6712 35756 6743
rect 36170 6740 36176 6792
rect 36228 6780 36234 6792
rect 36265 6783 36323 6789
rect 36265 6780 36277 6783
rect 36228 6752 36277 6780
rect 36228 6740 36234 6752
rect 36265 6749 36277 6752
rect 36311 6780 36323 6783
rect 36725 6783 36783 6789
rect 36725 6780 36737 6783
rect 36311 6752 36737 6780
rect 36311 6749 36323 6752
rect 36265 6743 36323 6749
rect 36725 6749 36737 6752
rect 36771 6749 36783 6783
rect 36725 6743 36783 6749
rect 36906 6740 36912 6792
rect 36964 6740 36970 6792
rect 35636 6684 35756 6712
rect 26973 6647 27031 6653
rect 26973 6613 26985 6647
rect 27019 6613 27031 6647
rect 26973 6607 27031 6613
rect 27157 6647 27215 6653
rect 27157 6613 27169 6647
rect 27203 6644 27215 6647
rect 27433 6647 27491 6653
rect 27433 6644 27445 6647
rect 27203 6616 27445 6644
rect 27203 6613 27215 6616
rect 27157 6607 27215 6613
rect 27433 6613 27445 6616
rect 27479 6613 27491 6647
rect 27433 6607 27491 6613
rect 30374 6604 30380 6656
rect 30432 6604 30438 6656
rect 32674 6604 32680 6656
rect 32732 6644 32738 6656
rect 32769 6647 32827 6653
rect 32769 6644 32781 6647
rect 32732 6616 32781 6644
rect 32732 6604 32738 6616
rect 32769 6613 32781 6616
rect 32815 6613 32827 6647
rect 32769 6607 32827 6613
rect 35342 6604 35348 6656
rect 35400 6644 35406 6656
rect 35636 6644 35664 6684
rect 35986 6672 35992 6724
rect 36044 6712 36050 6724
rect 36357 6715 36415 6721
rect 36357 6712 36369 6715
rect 36044 6684 36369 6712
rect 36044 6672 36050 6684
rect 36357 6681 36369 6684
rect 36403 6681 36415 6715
rect 36357 6675 36415 6681
rect 36541 6715 36599 6721
rect 36541 6681 36553 6715
rect 36587 6712 36599 6715
rect 36630 6712 36636 6724
rect 36587 6684 36636 6712
rect 36587 6681 36599 6684
rect 36541 6675 36599 6681
rect 36630 6672 36636 6684
rect 36688 6672 36694 6724
rect 35400 6616 35664 6644
rect 35713 6647 35771 6653
rect 35400 6604 35406 6616
rect 35713 6613 35725 6647
rect 35759 6644 35771 6647
rect 36262 6644 36268 6656
rect 35759 6616 36268 6644
rect 35759 6613 35771 6616
rect 35713 6607 35771 6613
rect 36262 6604 36268 6616
rect 36320 6604 36326 6656
rect 1104 6554 58880 6576
rect 1104 6502 4874 6554
rect 4926 6502 4938 6554
rect 4990 6502 5002 6554
rect 5054 6502 5066 6554
rect 5118 6502 5130 6554
rect 5182 6502 35594 6554
rect 35646 6502 35658 6554
rect 35710 6502 35722 6554
rect 35774 6502 35786 6554
rect 35838 6502 35850 6554
rect 35902 6502 58880 6554
rect 1104 6480 58880 6502
rect 12986 6400 12992 6452
rect 13044 6440 13050 6452
rect 13817 6443 13875 6449
rect 13044 6412 13768 6440
rect 13044 6400 13050 6412
rect 13630 6372 13636 6384
rect 13570 6344 13636 6372
rect 13630 6332 13636 6344
rect 13688 6332 13694 6384
rect 13740 6372 13768 6412
rect 13817 6409 13829 6443
rect 13863 6440 13875 6443
rect 14734 6440 14740 6452
rect 13863 6412 14740 6440
rect 13863 6409 13875 6412
rect 13817 6403 13875 6409
rect 14734 6400 14740 6412
rect 14792 6440 14798 6452
rect 15197 6443 15255 6449
rect 15197 6440 15209 6443
rect 14792 6412 15209 6440
rect 14792 6400 14798 6412
rect 15197 6409 15209 6412
rect 15243 6409 15255 6443
rect 15197 6403 15255 6409
rect 15565 6443 15623 6449
rect 15565 6409 15577 6443
rect 15611 6440 15623 6443
rect 19705 6443 19763 6449
rect 19705 6440 19717 6443
rect 15611 6412 15976 6440
rect 15611 6409 15623 6412
rect 15565 6403 15623 6409
rect 14918 6372 14924 6384
rect 13740 6344 14924 6372
rect 14918 6332 14924 6344
rect 14976 6332 14982 6384
rect 15212 6372 15240 6403
rect 15212 6344 15792 6372
rect 13909 6307 13967 6313
rect 13909 6273 13921 6307
rect 13955 6304 13967 6307
rect 13998 6304 14004 6316
rect 13955 6276 14004 6304
rect 13955 6273 13967 6276
rect 13909 6267 13967 6273
rect 13998 6264 14004 6276
rect 14056 6264 14062 6316
rect 14090 6264 14096 6316
rect 14148 6264 14154 6316
rect 14550 6264 14556 6316
rect 14608 6264 14614 6316
rect 14645 6307 14703 6313
rect 14645 6273 14657 6307
rect 14691 6304 14703 6307
rect 14691 6276 14780 6304
rect 14691 6273 14703 6276
rect 14645 6267 14703 6273
rect 12066 6196 12072 6248
rect 12124 6196 12130 6248
rect 12345 6239 12403 6245
rect 12345 6205 12357 6239
rect 12391 6236 12403 6239
rect 12986 6236 12992 6248
rect 12391 6208 12992 6236
rect 12391 6205 12403 6208
rect 12345 6199 12403 6205
rect 12986 6196 12992 6208
rect 13044 6196 13050 6248
rect 12084 6100 12112 6196
rect 14752 6180 14780 6276
rect 14826 6264 14832 6316
rect 14884 6264 14890 6316
rect 15105 6307 15163 6313
rect 15105 6273 15117 6307
rect 15151 6273 15163 6307
rect 15105 6267 15163 6273
rect 15289 6307 15347 6313
rect 15289 6273 15301 6307
rect 15335 6304 15347 6307
rect 15378 6304 15384 6316
rect 15335 6276 15384 6304
rect 15335 6273 15347 6276
rect 15289 6267 15347 6273
rect 15120 6236 15148 6267
rect 15378 6264 15384 6276
rect 15436 6264 15442 6316
rect 15764 6313 15792 6344
rect 15749 6307 15807 6313
rect 15749 6273 15761 6307
rect 15795 6273 15807 6307
rect 15948 6304 15976 6412
rect 16040 6412 19717 6440
rect 16040 6381 16068 6412
rect 19705 6409 19717 6412
rect 19751 6409 19763 6443
rect 19705 6403 19763 6409
rect 20438 6400 20444 6452
rect 20496 6440 20502 6452
rect 20533 6443 20591 6449
rect 20533 6440 20545 6443
rect 20496 6412 20545 6440
rect 20496 6400 20502 6412
rect 20533 6409 20545 6412
rect 20579 6409 20591 6443
rect 20533 6403 20591 6409
rect 20714 6400 20720 6452
rect 20772 6440 20778 6452
rect 21358 6440 21364 6452
rect 20772 6412 21364 6440
rect 20772 6400 20778 6412
rect 21358 6400 21364 6412
rect 21416 6400 21422 6452
rect 29089 6443 29147 6449
rect 29089 6409 29101 6443
rect 29135 6409 29147 6443
rect 29089 6403 29147 6409
rect 16025 6375 16083 6381
rect 16025 6341 16037 6375
rect 16071 6341 16083 6375
rect 19978 6372 19984 6384
rect 18722 6344 19984 6372
rect 16025 6335 16083 6341
rect 19978 6332 19984 6344
rect 20036 6332 20042 6384
rect 20622 6332 20628 6384
rect 20680 6372 20686 6384
rect 20680 6344 20944 6372
rect 20680 6332 20686 6344
rect 16850 6304 16856 6316
rect 15948 6276 16856 6304
rect 15749 6267 15807 6273
rect 16850 6264 16856 6276
rect 16908 6264 16914 6316
rect 17402 6264 17408 6316
rect 17460 6264 17466 6316
rect 17589 6307 17647 6313
rect 17589 6273 17601 6307
rect 17635 6304 17647 6307
rect 19705 6307 19763 6313
rect 17635 6276 17724 6304
rect 17635 6273 17647 6276
rect 17589 6267 17647 6273
rect 17696 6248 17724 6276
rect 19705 6273 19717 6307
rect 19751 6273 19763 6307
rect 19705 6267 19763 6273
rect 19889 6307 19947 6313
rect 19889 6273 19901 6307
rect 19935 6304 19947 6307
rect 20640 6304 20668 6332
rect 19935 6276 20668 6304
rect 20717 6307 20775 6313
rect 19935 6273 19947 6276
rect 19889 6267 19947 6273
rect 20717 6273 20729 6307
rect 20763 6304 20775 6307
rect 20806 6304 20812 6316
rect 20763 6276 20812 6304
rect 20763 6273 20775 6276
rect 20717 6267 20775 6273
rect 15120 6208 15792 6236
rect 14734 6128 14740 6180
rect 14792 6168 14798 6180
rect 15473 6171 15531 6177
rect 15473 6168 15485 6171
rect 14792 6140 15485 6168
rect 14792 6128 14798 6140
rect 15473 6137 15485 6140
rect 15519 6137 15531 6171
rect 15473 6131 15531 6137
rect 15764 6112 15792 6208
rect 15838 6196 15844 6248
rect 15896 6196 15902 6248
rect 17678 6196 17684 6248
rect 17736 6196 17742 6248
rect 19150 6196 19156 6248
rect 19208 6196 19214 6248
rect 19429 6239 19487 6245
rect 19429 6205 19441 6239
rect 19475 6205 19487 6239
rect 19720 6236 19748 6267
rect 20806 6264 20812 6276
rect 20864 6264 20870 6316
rect 20916 6313 20944 6344
rect 20990 6332 20996 6384
rect 21048 6372 21054 6384
rect 21910 6372 21916 6384
rect 21048 6344 21916 6372
rect 21048 6332 21054 6344
rect 21910 6332 21916 6344
rect 21968 6372 21974 6384
rect 29104 6372 29132 6403
rect 30374 6400 30380 6452
rect 30432 6400 30438 6452
rect 30561 6443 30619 6449
rect 30561 6409 30573 6443
rect 30607 6440 30619 6443
rect 30837 6443 30895 6449
rect 30837 6440 30849 6443
rect 30607 6412 30849 6440
rect 30607 6409 30619 6412
rect 30561 6403 30619 6409
rect 30837 6409 30849 6412
rect 30883 6409 30895 6443
rect 30837 6403 30895 6409
rect 35897 6443 35955 6449
rect 35897 6409 35909 6443
rect 35943 6440 35955 6443
rect 36354 6440 36360 6452
rect 35943 6412 36360 6440
rect 35943 6409 35955 6412
rect 35897 6403 35955 6409
rect 36354 6400 36360 6412
rect 36412 6400 36418 6452
rect 30469 6375 30527 6381
rect 30469 6372 30481 6375
rect 21968 6344 22126 6372
rect 29104 6344 30481 6372
rect 21968 6332 21974 6344
rect 30469 6341 30481 6344
rect 30515 6341 30527 6375
rect 30469 6335 30527 6341
rect 30745 6375 30803 6381
rect 30745 6341 30757 6375
rect 30791 6372 30803 6375
rect 34790 6372 34796 6384
rect 30791 6344 34796 6372
rect 30791 6341 30803 6344
rect 30745 6335 30803 6341
rect 34790 6332 34796 6344
rect 34848 6372 34854 6384
rect 35342 6372 35348 6384
rect 34848 6344 35348 6372
rect 34848 6332 34854 6344
rect 35342 6332 35348 6344
rect 35400 6332 35406 6384
rect 20901 6307 20959 6313
rect 20901 6273 20913 6307
rect 20947 6304 20959 6307
rect 27249 6307 27307 6313
rect 20947 6276 21496 6304
rect 20947 6273 20959 6276
rect 20901 6267 20959 6273
rect 20622 6236 20628 6248
rect 19720 6208 20628 6236
rect 19429 6199 19487 6205
rect 19444 6168 19472 6199
rect 20622 6196 20628 6208
rect 20680 6196 20686 6248
rect 21177 6239 21235 6245
rect 21177 6205 21189 6239
rect 21223 6205 21235 6239
rect 21177 6199 21235 6205
rect 21269 6239 21327 6245
rect 21269 6205 21281 6239
rect 21315 6205 21327 6239
rect 21269 6199 21327 6205
rect 19702 6168 19708 6180
rect 19444 6140 19708 6168
rect 19702 6128 19708 6140
rect 19760 6128 19766 6180
rect 20898 6128 20904 6180
rect 20956 6168 20962 6180
rect 21192 6168 21220 6199
rect 20956 6140 21220 6168
rect 21284 6168 21312 6199
rect 21358 6196 21364 6248
rect 21416 6196 21422 6248
rect 21468 6245 21496 6276
rect 27249 6273 27261 6307
rect 27295 6304 27307 6307
rect 27430 6304 27436 6316
rect 27295 6276 27436 6304
rect 27295 6273 27307 6276
rect 27249 6267 27307 6273
rect 27430 6264 27436 6276
rect 27488 6304 27494 6316
rect 27709 6307 27767 6313
rect 27709 6304 27721 6307
rect 27488 6276 27721 6304
rect 27488 6264 27494 6276
rect 27709 6273 27721 6276
rect 27755 6273 27767 6307
rect 27709 6267 27767 6273
rect 28721 6307 28779 6313
rect 28721 6273 28733 6307
rect 28767 6304 28779 6307
rect 29454 6304 29460 6316
rect 28767 6276 29460 6304
rect 28767 6273 28779 6276
rect 28721 6267 28779 6273
rect 29454 6264 29460 6276
rect 29512 6304 29518 6316
rect 29733 6307 29791 6313
rect 29733 6304 29745 6307
rect 29512 6276 29745 6304
rect 29512 6264 29518 6276
rect 29733 6273 29745 6276
rect 29779 6273 29791 6307
rect 29733 6267 29791 6273
rect 31205 6307 31263 6313
rect 31205 6273 31217 6307
rect 31251 6304 31263 6307
rect 31846 6304 31852 6316
rect 31251 6276 31852 6304
rect 31251 6273 31263 6276
rect 31205 6267 31263 6273
rect 31846 6264 31852 6276
rect 31904 6264 31910 6316
rect 33597 6307 33655 6313
rect 33597 6273 33609 6307
rect 33643 6304 33655 6307
rect 34514 6304 34520 6316
rect 33643 6276 34520 6304
rect 33643 6273 33655 6276
rect 33597 6267 33655 6273
rect 34514 6264 34520 6276
rect 34572 6264 34578 6316
rect 36170 6304 36176 6316
rect 36131 6276 36176 6304
rect 36170 6264 36176 6276
rect 36228 6264 36234 6316
rect 36262 6264 36268 6316
rect 36320 6264 36326 6316
rect 21453 6239 21511 6245
rect 21453 6205 21465 6239
rect 21499 6236 21511 6239
rect 21821 6239 21879 6245
rect 21821 6236 21833 6239
rect 21499 6208 21833 6236
rect 21499 6205 21511 6208
rect 21453 6199 21511 6205
rect 21821 6205 21833 6208
rect 21867 6205 21879 6239
rect 21821 6199 21879 6205
rect 23290 6196 23296 6248
rect 23348 6196 23354 6248
rect 23566 6196 23572 6248
rect 23624 6196 23630 6248
rect 27341 6239 27399 6245
rect 27341 6205 27353 6239
rect 27387 6236 27399 6239
rect 27798 6236 27804 6248
rect 27387 6208 27804 6236
rect 27387 6205 27399 6208
rect 27341 6199 27399 6205
rect 27798 6196 27804 6208
rect 27856 6196 27862 6248
rect 28626 6196 28632 6248
rect 28684 6196 28690 6248
rect 31297 6239 31355 6245
rect 31297 6205 31309 6239
rect 31343 6236 31355 6239
rect 31386 6236 31392 6248
rect 31343 6208 31392 6236
rect 31343 6205 31355 6208
rect 31297 6199 31355 6205
rect 31386 6196 31392 6208
rect 31444 6236 31450 6248
rect 31754 6236 31760 6248
rect 31444 6208 31760 6236
rect 31444 6196 31450 6208
rect 31754 6196 31760 6208
rect 31812 6196 31818 6248
rect 33689 6239 33747 6245
rect 33689 6205 33701 6239
rect 33735 6236 33747 6239
rect 33778 6236 33784 6248
rect 33735 6208 33784 6236
rect 33735 6205 33747 6208
rect 33689 6199 33747 6205
rect 33778 6196 33784 6208
rect 33836 6196 33842 6248
rect 33962 6196 33968 6248
rect 34020 6196 34026 6248
rect 36449 6239 36507 6245
rect 36449 6205 36461 6239
rect 36495 6236 36507 6239
rect 36630 6236 36636 6248
rect 36495 6208 36636 6236
rect 36495 6205 36507 6208
rect 36449 6199 36507 6205
rect 36630 6196 36636 6208
rect 36688 6196 36694 6248
rect 27617 6171 27675 6177
rect 21284 6140 21404 6168
rect 20956 6128 20962 6140
rect 21376 6112 21404 6140
rect 27617 6137 27629 6171
rect 27663 6168 27675 6171
rect 30193 6171 30251 6177
rect 30193 6168 30205 6171
rect 27663 6140 30205 6168
rect 27663 6137 27675 6140
rect 27617 6131 27675 6137
rect 30193 6137 30205 6140
rect 30239 6137 30251 6171
rect 30193 6131 30251 6137
rect 12342 6100 12348 6112
rect 12084 6072 12348 6100
rect 12342 6060 12348 6072
rect 12400 6060 12406 6112
rect 13906 6060 13912 6112
rect 13964 6060 13970 6112
rect 14274 6060 14280 6112
rect 14332 6100 14338 6112
rect 14829 6103 14887 6109
rect 14829 6100 14841 6103
rect 14332 6072 14841 6100
rect 14332 6060 14338 6072
rect 14829 6069 14841 6072
rect 14875 6069 14887 6103
rect 14829 6063 14887 6069
rect 15746 6060 15752 6112
rect 15804 6060 15810 6112
rect 17494 6060 17500 6112
rect 17552 6060 17558 6112
rect 20993 6103 21051 6109
rect 20993 6069 21005 6103
rect 21039 6100 21051 6103
rect 21082 6100 21088 6112
rect 21039 6072 21088 6100
rect 21039 6069 21051 6072
rect 20993 6063 21051 6069
rect 21082 6060 21088 6072
rect 21140 6060 21146 6112
rect 21358 6060 21364 6112
rect 21416 6060 21422 6112
rect 27890 6060 27896 6112
rect 27948 6100 27954 6112
rect 28353 6103 28411 6109
rect 28353 6100 28365 6103
rect 27948 6072 28365 6100
rect 27948 6060 27954 6072
rect 28353 6069 28365 6072
rect 28399 6069 28411 6103
rect 28353 6063 28411 6069
rect 29178 6060 29184 6112
rect 29236 6060 29242 6112
rect 36998 6060 37004 6112
rect 37056 6060 37062 6112
rect 1104 6010 58880 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 58880 6010
rect 1104 5936 58880 5958
rect 12986 5856 12992 5908
rect 13044 5856 13050 5908
rect 14550 5856 14556 5908
rect 14608 5856 14614 5908
rect 14826 5856 14832 5908
rect 14884 5856 14890 5908
rect 18138 5856 18144 5908
rect 18196 5856 18202 5908
rect 18325 5899 18383 5905
rect 18325 5865 18337 5899
rect 18371 5896 18383 5899
rect 19150 5896 19156 5908
rect 18371 5868 19156 5896
rect 18371 5865 18383 5868
rect 18325 5859 18383 5865
rect 19150 5856 19156 5868
rect 19208 5856 19214 5908
rect 20530 5856 20536 5908
rect 20588 5896 20594 5908
rect 20993 5899 21051 5905
rect 20993 5896 21005 5899
rect 20588 5868 21005 5896
rect 20588 5856 20594 5868
rect 20993 5865 21005 5868
rect 21039 5896 21051 5899
rect 21358 5896 21364 5908
rect 21039 5868 21364 5896
rect 21039 5865 21051 5868
rect 20993 5859 21051 5865
rect 21358 5856 21364 5868
rect 21416 5856 21422 5908
rect 21453 5899 21511 5905
rect 21453 5865 21465 5899
rect 21499 5896 21511 5899
rect 23290 5896 23296 5908
rect 21499 5868 23296 5896
rect 21499 5865 21511 5868
rect 21453 5859 21511 5865
rect 23290 5856 23296 5868
rect 23348 5856 23354 5908
rect 27430 5856 27436 5908
rect 27488 5856 27494 5908
rect 29270 5856 29276 5908
rect 29328 5896 29334 5908
rect 29549 5899 29607 5905
rect 29549 5896 29561 5899
rect 29328 5868 29561 5896
rect 29328 5856 29334 5868
rect 29549 5865 29561 5868
rect 29595 5865 29607 5899
rect 29549 5859 29607 5865
rect 31846 5856 31852 5908
rect 31904 5856 31910 5908
rect 34514 5856 34520 5908
rect 34572 5856 34578 5908
rect 36170 5856 36176 5908
rect 36228 5896 36234 5908
rect 36228 5868 36308 5896
rect 36228 5856 36234 5868
rect 14369 5831 14427 5837
rect 14369 5828 14381 5831
rect 14108 5800 14381 5828
rect 12805 5695 12863 5701
rect 12805 5661 12817 5695
rect 12851 5692 12863 5695
rect 12894 5692 12900 5704
rect 12851 5664 12900 5692
rect 12851 5661 12863 5664
rect 12805 5655 12863 5661
rect 12894 5652 12900 5664
rect 12952 5652 12958 5704
rect 12989 5695 13047 5701
rect 12989 5661 13001 5695
rect 13035 5692 13047 5695
rect 13906 5692 13912 5704
rect 13035 5664 13912 5692
rect 13035 5661 13047 5664
rect 12989 5655 13047 5661
rect 13906 5652 13912 5664
rect 13964 5652 13970 5704
rect 13998 5652 14004 5704
rect 14056 5692 14062 5704
rect 14108 5701 14136 5800
rect 14369 5797 14381 5800
rect 14415 5797 14427 5831
rect 14568 5828 14596 5856
rect 15378 5828 15384 5840
rect 14568 5800 15384 5828
rect 14369 5791 14427 5797
rect 15378 5788 15384 5800
rect 15436 5828 15442 5840
rect 27525 5831 27583 5837
rect 15436 5800 16712 5828
rect 15436 5788 15442 5800
rect 15473 5763 15531 5769
rect 15473 5729 15485 5763
rect 15519 5760 15531 5763
rect 15746 5760 15752 5772
rect 15519 5732 15752 5760
rect 15519 5729 15531 5732
rect 15473 5723 15531 5729
rect 14093 5695 14151 5701
rect 14093 5692 14105 5695
rect 14056 5664 14105 5692
rect 14056 5652 14062 5664
rect 14093 5661 14105 5664
rect 14139 5661 14151 5695
rect 14093 5655 14151 5661
rect 14274 5652 14280 5704
rect 14332 5652 14338 5704
rect 15488 5692 15516 5723
rect 15746 5720 15752 5732
rect 15804 5720 15810 5772
rect 15838 5720 15844 5772
rect 15896 5760 15902 5772
rect 16301 5763 16359 5769
rect 16301 5760 16313 5763
rect 15896 5732 16313 5760
rect 15896 5720 15902 5732
rect 16301 5729 16313 5732
rect 16347 5729 16359 5763
rect 16301 5723 16359 5729
rect 14660 5664 15516 5692
rect 16025 5695 16083 5701
rect 14550 5633 14556 5636
rect 14537 5627 14556 5633
rect 14537 5593 14549 5627
rect 14608 5624 14614 5636
rect 14660 5624 14688 5664
rect 16025 5661 16037 5695
rect 16071 5692 16083 5695
rect 16574 5692 16580 5704
rect 16071 5664 16580 5692
rect 16071 5661 16083 5664
rect 16025 5655 16083 5661
rect 16574 5652 16580 5664
rect 16632 5652 16638 5704
rect 14608 5596 14688 5624
rect 14537 5587 14556 5593
rect 14550 5584 14556 5587
rect 14608 5584 14614 5596
rect 14734 5584 14740 5636
rect 14792 5624 14798 5636
rect 16482 5624 16488 5636
rect 14792 5596 16488 5624
rect 14792 5584 14798 5596
rect 16482 5584 16488 5596
rect 16540 5584 16546 5636
rect 16684 5633 16712 5800
rect 27525 5797 27537 5831
rect 27571 5797 27583 5831
rect 27525 5791 27583 5797
rect 18509 5763 18567 5769
rect 18509 5760 18521 5763
rect 18156 5732 18521 5760
rect 16942 5652 16948 5704
rect 17000 5692 17006 5704
rect 17770 5692 17776 5704
rect 17000 5664 17776 5692
rect 17000 5652 17006 5664
rect 17770 5652 17776 5664
rect 17828 5652 17834 5704
rect 16669 5627 16727 5633
rect 16669 5593 16681 5627
rect 16715 5624 16727 5627
rect 16850 5624 16856 5636
rect 16715 5596 16856 5624
rect 16715 5593 16727 5596
rect 16669 5587 16727 5593
rect 16850 5584 16856 5596
rect 16908 5584 16914 5636
rect 17494 5584 17500 5636
rect 17552 5624 17558 5636
rect 18156 5633 18184 5732
rect 18509 5729 18521 5732
rect 18555 5729 18567 5763
rect 18509 5723 18567 5729
rect 19245 5763 19303 5769
rect 19245 5729 19257 5763
rect 19291 5760 19303 5763
rect 19610 5760 19616 5772
rect 19291 5732 19616 5760
rect 19291 5729 19303 5732
rect 19245 5723 19303 5729
rect 19610 5720 19616 5732
rect 19668 5720 19674 5772
rect 19978 5720 19984 5772
rect 20036 5760 20042 5772
rect 20714 5760 20720 5772
rect 20036 5732 20720 5760
rect 20036 5720 20042 5732
rect 20714 5720 20720 5732
rect 20772 5760 20778 5772
rect 20990 5760 20996 5772
rect 20772 5732 20996 5760
rect 20772 5720 20778 5732
rect 20990 5720 20996 5732
rect 21048 5720 21054 5772
rect 21082 5720 21088 5772
rect 21140 5720 21146 5772
rect 25961 5763 26019 5769
rect 25961 5729 25973 5763
rect 26007 5760 26019 5763
rect 27540 5760 27568 5791
rect 26007 5732 27568 5760
rect 28169 5763 28227 5769
rect 26007 5729 26019 5732
rect 25961 5723 26019 5729
rect 28169 5729 28181 5763
rect 28215 5760 28227 5763
rect 28997 5763 29055 5769
rect 28997 5760 29009 5763
rect 28215 5732 29009 5760
rect 28215 5729 28227 5732
rect 28169 5723 28227 5729
rect 28997 5729 29009 5732
rect 29043 5760 29055 5763
rect 29288 5760 29316 5856
rect 29043 5732 29316 5760
rect 30101 5763 30159 5769
rect 29043 5729 29055 5732
rect 28997 5723 29055 5729
rect 30101 5729 30113 5763
rect 30147 5760 30159 5763
rect 34532 5760 34560 5856
rect 36280 5828 36308 5868
rect 36630 5856 36636 5908
rect 36688 5856 36694 5908
rect 37366 5856 37372 5908
rect 37424 5896 37430 5908
rect 37461 5899 37519 5905
rect 37461 5896 37473 5899
rect 37424 5868 37473 5896
rect 37424 5856 37430 5868
rect 37461 5865 37473 5868
rect 37507 5865 37519 5899
rect 37461 5859 37519 5865
rect 37553 5831 37611 5837
rect 37553 5828 37565 5831
rect 36280 5800 37565 5828
rect 37553 5797 37565 5800
rect 37599 5797 37611 5831
rect 37553 5791 37611 5797
rect 35253 5763 35311 5769
rect 35253 5760 35265 5763
rect 30147 5732 32812 5760
rect 34532 5732 35265 5760
rect 30147 5729 30159 5732
rect 30101 5723 30159 5729
rect 32784 5704 32812 5732
rect 35253 5729 35265 5732
rect 35299 5729 35311 5763
rect 35253 5723 35311 5729
rect 36081 5763 36139 5769
rect 36081 5729 36093 5763
rect 36127 5729 36139 5763
rect 36081 5723 36139 5729
rect 18601 5695 18659 5701
rect 18601 5661 18613 5695
rect 18647 5661 18659 5695
rect 18601 5655 18659 5661
rect 18141 5627 18199 5633
rect 18141 5624 18153 5627
rect 17552 5596 18153 5624
rect 17552 5584 17558 5596
rect 18141 5593 18153 5596
rect 18187 5593 18199 5627
rect 18616 5624 18644 5655
rect 21266 5652 21272 5704
rect 21324 5652 21330 5704
rect 24762 5652 24768 5704
rect 24820 5692 24826 5704
rect 25685 5695 25743 5701
rect 25685 5692 25697 5695
rect 24820 5664 25697 5692
rect 24820 5652 24826 5664
rect 25685 5661 25697 5664
rect 25731 5661 25743 5695
rect 25685 5655 25743 5661
rect 27890 5652 27896 5704
rect 27948 5652 27954 5704
rect 28721 5695 28779 5701
rect 28721 5661 28733 5695
rect 28767 5692 28779 5695
rect 29178 5692 29184 5704
rect 28767 5664 29184 5692
rect 28767 5661 28779 5664
rect 28721 5655 28779 5661
rect 29178 5652 29184 5664
rect 29236 5652 29242 5704
rect 31846 5652 31852 5704
rect 31904 5692 31910 5704
rect 32493 5695 32551 5701
rect 32493 5692 32505 5695
rect 31904 5664 32505 5692
rect 31904 5652 31910 5664
rect 32493 5661 32505 5664
rect 32539 5661 32551 5695
rect 32493 5655 32551 5661
rect 32766 5652 32772 5704
rect 32824 5652 32830 5704
rect 36096 5692 36124 5723
rect 36096 5664 36216 5692
rect 19426 5624 19432 5636
rect 18616 5596 19432 5624
rect 18141 5587 18199 5593
rect 19426 5584 19432 5596
rect 19484 5584 19490 5636
rect 19521 5627 19579 5633
rect 19521 5593 19533 5627
rect 19567 5593 19579 5627
rect 19521 5587 19579 5593
rect 13814 5516 13820 5568
rect 13872 5556 13878 5568
rect 14185 5559 14243 5565
rect 14185 5556 14197 5559
rect 13872 5528 14197 5556
rect 13872 5516 13878 5528
rect 14185 5525 14197 5528
rect 14231 5525 14243 5559
rect 14185 5519 14243 5525
rect 16206 5516 16212 5568
rect 16264 5516 16270 5568
rect 18969 5559 19027 5565
rect 18969 5525 18981 5559
rect 19015 5556 19027 5559
rect 19536 5556 19564 5587
rect 19978 5584 19984 5636
rect 20036 5584 20042 5636
rect 27614 5624 27620 5636
rect 27186 5596 27620 5624
rect 27614 5584 27620 5596
rect 27672 5584 27678 5636
rect 30374 5584 30380 5636
rect 30432 5584 30438 5636
rect 30466 5584 30472 5636
rect 30524 5624 30530 5636
rect 33045 5627 33103 5633
rect 30524 5596 30866 5624
rect 31726 5596 32904 5624
rect 30524 5584 30530 5596
rect 19015 5528 19564 5556
rect 19015 5525 19027 5528
rect 18969 5519 19027 5525
rect 27890 5516 27896 5568
rect 27948 5556 27954 5568
rect 27985 5559 28043 5565
rect 27985 5556 27997 5559
rect 27948 5528 27997 5556
rect 27948 5516 27954 5528
rect 27985 5525 27997 5528
rect 28031 5525 28043 5559
rect 27985 5519 28043 5525
rect 28074 5516 28080 5568
rect 28132 5556 28138 5568
rect 28353 5559 28411 5565
rect 28353 5556 28365 5559
rect 28132 5528 28365 5556
rect 28132 5516 28138 5528
rect 28353 5525 28365 5528
rect 28399 5525 28411 5559
rect 28353 5519 28411 5525
rect 28718 5516 28724 5568
rect 28776 5556 28782 5568
rect 28813 5559 28871 5565
rect 28813 5556 28825 5559
rect 28776 5528 28825 5556
rect 28776 5516 28782 5528
rect 28813 5525 28825 5528
rect 28859 5525 28871 5559
rect 30760 5556 30788 5596
rect 31726 5556 31754 5596
rect 32876 5568 32904 5596
rect 33045 5593 33057 5627
rect 33091 5624 33103 5627
rect 33318 5624 33324 5636
rect 33091 5596 33324 5624
rect 33091 5593 33103 5596
rect 33045 5587 33103 5593
rect 33318 5584 33324 5596
rect 33376 5584 33382 5636
rect 36188 5624 36216 5664
rect 36262 5652 36268 5704
rect 36320 5692 36326 5704
rect 37277 5695 37335 5701
rect 37277 5692 37289 5695
rect 36320 5664 37289 5692
rect 36320 5652 36326 5664
rect 37277 5661 37289 5664
rect 37323 5692 37335 5695
rect 37921 5695 37979 5701
rect 37921 5692 37933 5695
rect 37323 5664 37933 5692
rect 37323 5661 37335 5664
rect 37277 5655 37335 5661
rect 37921 5661 37933 5664
rect 37967 5661 37979 5695
rect 37921 5655 37979 5661
rect 37826 5624 37832 5636
rect 33428 5596 33534 5624
rect 36188 5596 37832 5624
rect 30760 5528 31754 5556
rect 28813 5519 28871 5525
rect 31938 5516 31944 5568
rect 31996 5516 32002 5568
rect 32858 5516 32864 5568
rect 32916 5556 32922 5568
rect 33428 5556 33456 5596
rect 37826 5584 37832 5596
rect 37884 5584 37890 5636
rect 32916 5528 33456 5556
rect 32916 5516 32922 5528
rect 34698 5516 34704 5568
rect 34756 5516 34762 5568
rect 36170 5516 36176 5568
rect 36228 5516 36234 5568
rect 36265 5559 36323 5565
rect 36265 5525 36277 5559
rect 36311 5556 36323 5559
rect 36725 5559 36783 5565
rect 36725 5556 36737 5559
rect 36311 5528 36737 5556
rect 36311 5525 36323 5528
rect 36265 5519 36323 5525
rect 36725 5525 36737 5528
rect 36771 5525 36783 5559
rect 36725 5519 36783 5525
rect 1104 5466 58880 5488
rect 1104 5414 4874 5466
rect 4926 5414 4938 5466
rect 4990 5414 5002 5466
rect 5054 5414 5066 5466
rect 5118 5414 5130 5466
rect 5182 5414 35594 5466
rect 35646 5414 35658 5466
rect 35710 5414 35722 5466
rect 35774 5414 35786 5466
rect 35838 5414 35850 5466
rect 35902 5414 58880 5466
rect 1104 5392 58880 5414
rect 13464 5324 14504 5352
rect 13464 5284 13492 5324
rect 13538 5284 13544 5296
rect 13464 5256 13544 5284
rect 13538 5244 13544 5256
rect 13596 5244 13602 5296
rect 14476 5284 14504 5324
rect 14550 5312 14556 5364
rect 14608 5312 14614 5364
rect 14734 5312 14740 5364
rect 14792 5312 14798 5364
rect 15286 5312 15292 5364
rect 15344 5352 15350 5364
rect 15562 5352 15568 5364
rect 15344 5324 15568 5352
rect 15344 5312 15350 5324
rect 15562 5312 15568 5324
rect 15620 5352 15626 5364
rect 15620 5324 16528 5352
rect 15620 5312 15626 5324
rect 14476 5270 15042 5284
rect 14476 5256 15056 5270
rect 12342 5176 12348 5228
rect 12400 5216 12406 5228
rect 12805 5219 12863 5225
rect 12805 5216 12817 5219
rect 12400 5188 12817 5216
rect 12400 5176 12406 5188
rect 12805 5185 12817 5188
rect 12851 5185 12863 5219
rect 12805 5179 12863 5185
rect 13081 5151 13139 5157
rect 13081 5117 13093 5151
rect 13127 5148 13139 5151
rect 13814 5148 13820 5160
rect 13127 5120 13820 5148
rect 13127 5117 13139 5120
rect 13081 5111 13139 5117
rect 13814 5108 13820 5120
rect 13872 5108 13878 5160
rect 15028 5148 15056 5256
rect 16206 5244 16212 5296
rect 16264 5244 16270 5296
rect 16500 5225 16528 5324
rect 16574 5312 16580 5364
rect 16632 5352 16638 5364
rect 16669 5355 16727 5361
rect 16669 5352 16681 5355
rect 16632 5324 16681 5352
rect 16632 5312 16638 5324
rect 16669 5321 16681 5324
rect 16715 5321 16727 5355
rect 16669 5315 16727 5321
rect 19426 5312 19432 5364
rect 19484 5352 19490 5364
rect 19889 5355 19947 5361
rect 19889 5352 19901 5355
rect 19484 5324 19901 5352
rect 19484 5312 19490 5324
rect 19889 5321 19901 5324
rect 19935 5321 19947 5355
rect 24762 5352 24768 5364
rect 19889 5315 19947 5321
rect 23768 5324 24768 5352
rect 23566 5244 23572 5296
rect 23624 5284 23630 5296
rect 23768 5284 23796 5324
rect 24762 5312 24768 5324
rect 24820 5312 24826 5364
rect 25409 5355 25467 5361
rect 25409 5321 25421 5355
rect 25455 5352 25467 5355
rect 26234 5352 26240 5364
rect 25455 5324 26240 5352
rect 25455 5321 25467 5324
rect 25409 5315 25467 5321
rect 26234 5312 26240 5324
rect 26292 5312 26298 5364
rect 27614 5312 27620 5364
rect 27672 5352 27678 5364
rect 27798 5352 27804 5364
rect 27672 5324 27804 5352
rect 27672 5312 27678 5324
rect 27798 5312 27804 5324
rect 27856 5352 27862 5364
rect 28166 5352 28172 5364
rect 27856 5324 28172 5352
rect 27856 5312 27862 5324
rect 28166 5312 28172 5324
rect 28224 5312 28230 5364
rect 29454 5312 29460 5364
rect 29512 5312 29518 5364
rect 30374 5312 30380 5364
rect 30432 5352 30438 5364
rect 30929 5355 30987 5361
rect 30929 5352 30941 5355
rect 30432 5324 30941 5352
rect 30432 5312 30438 5324
rect 30929 5321 30941 5324
rect 30975 5321 30987 5355
rect 30929 5315 30987 5321
rect 31297 5355 31355 5361
rect 31297 5321 31309 5355
rect 31343 5352 31355 5355
rect 31938 5352 31944 5364
rect 31343 5324 31944 5352
rect 31343 5321 31355 5324
rect 31297 5315 31355 5321
rect 31938 5312 31944 5324
rect 31996 5312 32002 5364
rect 33318 5312 33324 5364
rect 33376 5312 33382 5364
rect 33689 5355 33747 5361
rect 33689 5321 33701 5355
rect 33735 5352 33747 5355
rect 34698 5352 34704 5364
rect 33735 5324 34704 5352
rect 33735 5321 33747 5324
rect 33689 5315 33747 5321
rect 34698 5312 34704 5324
rect 34756 5312 34762 5364
rect 35529 5355 35587 5361
rect 35529 5321 35541 5355
rect 35575 5352 35587 5355
rect 36262 5352 36268 5364
rect 35575 5324 36268 5352
rect 35575 5321 35587 5324
rect 35529 5315 35587 5321
rect 36262 5312 36268 5324
rect 36320 5312 36326 5364
rect 37366 5352 37372 5364
rect 36372 5324 37372 5352
rect 26050 5284 26056 5296
rect 23624 5256 23796 5284
rect 25162 5256 26056 5284
rect 23624 5244 23630 5256
rect 16485 5219 16543 5225
rect 16485 5185 16497 5219
rect 16531 5185 16543 5219
rect 16485 5179 16543 5185
rect 16574 5176 16580 5228
rect 16632 5216 16638 5228
rect 16669 5219 16727 5225
rect 16669 5216 16681 5219
rect 16632 5188 16681 5216
rect 16632 5176 16638 5188
rect 16669 5185 16681 5188
rect 16715 5185 16727 5219
rect 16669 5179 16727 5185
rect 16850 5176 16856 5228
rect 16908 5216 16914 5228
rect 17310 5216 17316 5228
rect 16908 5188 17316 5216
rect 16908 5176 16914 5188
rect 17310 5176 17316 5188
rect 17368 5176 17374 5228
rect 20530 5176 20536 5228
rect 20588 5176 20594 5228
rect 23676 5225 23704 5256
rect 26050 5244 26056 5256
rect 26108 5244 26114 5296
rect 27985 5287 28043 5293
rect 27985 5253 27997 5287
rect 28031 5284 28043 5287
rect 28074 5284 28080 5296
rect 28031 5256 28080 5284
rect 28031 5253 28043 5256
rect 27985 5247 28043 5253
rect 28074 5244 28080 5256
rect 28132 5244 28138 5296
rect 28184 5284 28212 5312
rect 28184 5256 28474 5284
rect 31662 5244 31668 5296
rect 31720 5284 31726 5296
rect 31757 5287 31815 5293
rect 31757 5284 31769 5287
rect 31720 5256 31769 5284
rect 31720 5244 31726 5256
rect 31757 5253 31769 5256
rect 31803 5253 31815 5287
rect 31757 5247 31815 5253
rect 23661 5219 23719 5225
rect 23661 5185 23673 5219
rect 23707 5185 23719 5219
rect 23661 5179 23719 5185
rect 16114 5148 16120 5160
rect 15028 5120 16120 5148
rect 16114 5108 16120 5120
rect 16172 5108 16178 5160
rect 23934 5108 23940 5160
rect 23992 5108 23998 5160
rect 27709 5151 27767 5157
rect 27709 5117 27721 5151
rect 27755 5117 27767 5151
rect 27709 5111 27767 5117
rect 27724 5012 27752 5111
rect 31386 5108 31392 5160
rect 31444 5108 31450 5160
rect 31573 5151 31631 5157
rect 31573 5117 31585 5151
rect 31619 5148 31631 5151
rect 31680 5148 31708 5244
rect 36372 5216 36400 5324
rect 37366 5312 37372 5324
rect 37424 5312 37430 5364
rect 36664 5287 36722 5293
rect 36664 5253 36676 5287
rect 36710 5284 36722 5287
rect 36998 5284 37004 5296
rect 36710 5256 37004 5284
rect 36710 5253 36722 5256
rect 36664 5247 36722 5253
rect 36998 5244 37004 5256
rect 37056 5244 37062 5296
rect 33980 5188 36400 5216
rect 36909 5219 36967 5225
rect 31619 5120 31708 5148
rect 31619 5117 31631 5120
rect 31573 5111 31631 5117
rect 33778 5108 33784 5160
rect 33836 5108 33842 5160
rect 33980 5157 34008 5188
rect 36909 5185 36921 5219
rect 36955 5216 36967 5219
rect 37090 5216 37096 5228
rect 36955 5188 37096 5216
rect 36955 5185 36967 5188
rect 36909 5179 36967 5185
rect 37090 5176 37096 5188
rect 37148 5176 37154 5228
rect 33965 5151 34023 5157
rect 33965 5117 33977 5151
rect 34011 5117 34023 5151
rect 33965 5111 34023 5117
rect 34146 5108 34152 5160
rect 34204 5108 34210 5160
rect 28074 5012 28080 5024
rect 27724 4984 28080 5012
rect 28074 4972 28080 4984
rect 28132 4972 28138 5024
rect 34790 4972 34796 5024
rect 34848 4972 34854 5024
rect 1104 4922 58880 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 58880 4922
rect 1104 4848 58880 4870
rect 17770 4808 17776 4820
rect 15488 4780 17776 4808
rect 15488 4613 15516 4780
rect 17770 4768 17776 4780
rect 17828 4768 17834 4820
rect 23753 4811 23811 4817
rect 23753 4777 23765 4811
rect 23799 4808 23811 4811
rect 23934 4808 23940 4820
rect 23799 4780 23940 4808
rect 23799 4777 23811 4780
rect 23753 4771 23811 4777
rect 23934 4768 23940 4780
rect 23992 4768 23998 4820
rect 26142 4768 26148 4820
rect 26200 4768 26206 4820
rect 27706 4768 27712 4820
rect 27764 4768 27770 4820
rect 33229 4811 33287 4817
rect 33229 4777 33241 4811
rect 33275 4808 33287 4811
rect 34146 4808 34152 4820
rect 33275 4780 34152 4808
rect 33275 4777 33287 4780
rect 33229 4771 33287 4777
rect 34146 4768 34152 4780
rect 34204 4768 34210 4820
rect 34517 4811 34575 4817
rect 34517 4777 34529 4811
rect 34563 4808 34575 4811
rect 34606 4808 34612 4820
rect 34563 4780 34612 4808
rect 34563 4777 34575 4780
rect 34517 4771 34575 4777
rect 34606 4768 34612 4780
rect 34664 4768 34670 4820
rect 34790 4768 34796 4820
rect 34848 4768 34854 4820
rect 36170 4768 36176 4820
rect 36228 4808 36234 4820
rect 36449 4811 36507 4817
rect 36449 4808 36461 4811
rect 36228 4780 36461 4808
rect 36228 4768 36234 4780
rect 36449 4777 36461 4780
rect 36495 4777 36507 4811
rect 36449 4771 36507 4777
rect 15562 4632 15568 4684
rect 15620 4632 15626 4684
rect 21177 4675 21235 4681
rect 21177 4641 21189 4675
rect 21223 4672 21235 4675
rect 21910 4672 21916 4684
rect 21223 4644 21916 4672
rect 21223 4641 21235 4644
rect 21177 4635 21235 4641
rect 21910 4632 21916 4644
rect 21968 4672 21974 4684
rect 22557 4675 22615 4681
rect 22557 4672 22569 4675
rect 21968 4644 22569 4672
rect 21968 4632 21974 4644
rect 22557 4641 22569 4644
rect 22603 4641 22615 4675
rect 22557 4635 22615 4641
rect 24397 4675 24455 4681
rect 24397 4641 24409 4675
rect 24443 4672 24455 4675
rect 24762 4672 24768 4684
rect 24443 4644 24768 4672
rect 24443 4641 24455 4644
rect 24397 4635 24455 4641
rect 24762 4632 24768 4644
rect 24820 4632 24826 4684
rect 31478 4672 31484 4684
rect 31439 4644 31484 4672
rect 31478 4632 31484 4644
rect 31536 4672 31542 4684
rect 32766 4672 32772 4684
rect 31536 4644 32772 4672
rect 31536 4632 31542 4644
rect 32766 4632 32772 4644
rect 32824 4672 32830 4684
rect 34701 4675 34759 4681
rect 34701 4672 34713 4675
rect 32824 4644 34713 4672
rect 32824 4632 32830 4644
rect 34701 4641 34713 4644
rect 34747 4641 34759 4675
rect 34808 4672 34836 4768
rect 34977 4675 35035 4681
rect 34977 4672 34989 4675
rect 34808 4644 34989 4672
rect 34701 4635 34759 4641
rect 34977 4641 34989 4644
rect 35023 4641 35035 4675
rect 34977 4635 35035 4641
rect 15289 4607 15347 4613
rect 15289 4573 15301 4607
rect 15335 4573 15347 4607
rect 15289 4567 15347 4573
rect 15473 4607 15531 4613
rect 15473 4573 15485 4607
rect 15519 4573 15531 4607
rect 23569 4607 23627 4613
rect 23569 4604 23581 4607
rect 15473 4567 15531 4573
rect 23216 4576 23581 4604
rect 15304 4468 15332 4567
rect 15381 4539 15439 4545
rect 15381 4505 15393 4539
rect 15427 4536 15439 4539
rect 15841 4539 15899 4545
rect 15841 4536 15853 4539
rect 15427 4508 15853 4536
rect 15427 4505 15439 4508
rect 15381 4499 15439 4505
rect 15841 4505 15853 4508
rect 15887 4505 15899 4539
rect 15841 4499 15899 4505
rect 16114 4496 16120 4548
rect 16172 4536 16178 4548
rect 20901 4539 20959 4545
rect 16172 4508 16330 4536
rect 16172 4496 16178 4508
rect 20901 4505 20913 4539
rect 20947 4536 20959 4539
rect 22922 4536 22928 4548
rect 20947 4508 22928 4536
rect 20947 4505 20959 4508
rect 20901 4499 20959 4505
rect 22922 4496 22928 4508
rect 22980 4496 22986 4548
rect 23216 4480 23244 4576
rect 23569 4573 23581 4576
rect 23615 4573 23627 4607
rect 23569 4567 23627 4573
rect 23753 4607 23811 4613
rect 23753 4573 23765 4607
rect 23799 4573 23811 4607
rect 23753 4567 23811 4573
rect 23382 4496 23388 4548
rect 23440 4536 23446 4548
rect 23768 4536 23796 4567
rect 27706 4564 27712 4616
rect 27764 4604 27770 4616
rect 28813 4607 28871 4613
rect 28813 4604 28825 4607
rect 27764 4576 28825 4604
rect 27764 4564 27770 4576
rect 28813 4573 28825 4576
rect 28859 4573 28871 4607
rect 28813 4567 28871 4573
rect 30742 4564 30748 4616
rect 30800 4604 30806 4616
rect 30837 4607 30895 4613
rect 30837 4604 30849 4607
rect 30800 4576 30849 4604
rect 30800 4564 30806 4576
rect 30837 4573 30849 4576
rect 30883 4573 30895 4607
rect 30837 4567 30895 4573
rect 32858 4564 32864 4616
rect 32916 4564 32922 4616
rect 23440 4508 23796 4536
rect 23440 4496 23446 4508
rect 24670 4496 24676 4548
rect 24728 4496 24734 4548
rect 26050 4536 26056 4548
rect 25898 4508 26056 4536
rect 26050 4496 26056 4508
rect 26108 4536 26114 4548
rect 27798 4536 27804 4548
rect 26108 4508 27804 4536
rect 26108 4496 26114 4508
rect 27798 4496 27804 4508
rect 27856 4496 27862 4548
rect 28074 4496 28080 4548
rect 28132 4496 28138 4548
rect 30929 4539 30987 4545
rect 30929 4505 30941 4539
rect 30975 4536 30987 4539
rect 31757 4539 31815 4545
rect 31757 4536 31769 4539
rect 30975 4508 31769 4536
rect 30975 4505 30987 4508
rect 30929 4499 30987 4505
rect 31757 4505 31769 4508
rect 31803 4505 31815 4539
rect 31757 4499 31815 4505
rect 34606 4496 34612 4548
rect 34664 4536 34670 4548
rect 34664 4508 35466 4536
rect 34664 4496 34670 4508
rect 16666 4468 16672 4480
rect 15304 4440 16672 4468
rect 16666 4428 16672 4440
rect 16724 4428 16730 4480
rect 17310 4428 17316 4480
rect 17368 4428 17374 4480
rect 19978 4428 19984 4480
rect 20036 4468 20042 4480
rect 20533 4471 20591 4477
rect 20533 4468 20545 4471
rect 20036 4440 20545 4468
rect 20036 4428 20042 4440
rect 20533 4437 20545 4440
rect 20579 4437 20591 4471
rect 20533 4431 20591 4437
rect 20993 4471 21051 4477
rect 20993 4437 21005 4471
rect 21039 4468 21051 4471
rect 21174 4468 21180 4480
rect 21039 4440 21180 4468
rect 21039 4437 21051 4440
rect 20993 4431 21051 4437
rect 21174 4428 21180 4440
rect 21232 4428 21238 4480
rect 23198 4428 23204 4480
rect 23256 4428 23262 4480
rect 1104 4378 58880 4400
rect 1104 4326 4874 4378
rect 4926 4326 4938 4378
rect 4990 4326 5002 4378
rect 5054 4326 5066 4378
rect 5118 4326 5130 4378
rect 5182 4326 35594 4378
rect 35646 4326 35658 4378
rect 35710 4326 35722 4378
rect 35774 4326 35786 4378
rect 35838 4326 35850 4378
rect 35902 4326 58880 4378
rect 1104 4304 58880 4326
rect 22649 4267 22707 4273
rect 22649 4233 22661 4267
rect 22695 4264 22707 4267
rect 23198 4264 23204 4276
rect 22695 4236 23204 4264
rect 22695 4233 22707 4236
rect 22649 4227 22707 4233
rect 23198 4224 23204 4236
rect 23256 4224 23262 4276
rect 19978 4156 19984 4208
rect 20036 4156 20042 4208
rect 20714 4156 20720 4208
rect 20772 4156 20778 4208
rect 22833 4199 22891 4205
rect 22833 4165 22845 4199
rect 22879 4196 22891 4199
rect 23474 4196 23480 4208
rect 22879 4168 23480 4196
rect 22879 4165 22891 4168
rect 22833 4159 22891 4165
rect 23474 4156 23480 4168
rect 23532 4156 23538 4208
rect 26050 4196 26056 4208
rect 24978 4168 26056 4196
rect 26050 4156 26056 4168
rect 26108 4156 26114 4208
rect 27249 4199 27307 4205
rect 27249 4196 27261 4199
rect 26988 4168 27261 4196
rect 16666 4088 16672 4140
rect 16724 4088 16730 4140
rect 17310 4088 17316 4140
rect 17368 4088 17374 4140
rect 22554 4088 22560 4140
rect 22612 4088 22618 4140
rect 22922 4088 22928 4140
rect 22980 4088 22986 4140
rect 23106 4088 23112 4140
rect 23164 4088 23170 4140
rect 25314 4088 25320 4140
rect 25372 4128 25378 4140
rect 26329 4131 26387 4137
rect 26329 4128 26341 4131
rect 25372 4100 26341 4128
rect 25372 4088 25378 4100
rect 26329 4097 26341 4100
rect 26375 4097 26387 4131
rect 26329 4091 26387 4097
rect 26510 4088 26516 4140
rect 26568 4088 26574 4140
rect 26988 4128 27016 4168
rect 27249 4165 27261 4168
rect 27295 4165 27307 4199
rect 27249 4159 27307 4165
rect 27798 4156 27804 4208
rect 27856 4156 27862 4208
rect 26896 4100 27016 4128
rect 19702 4020 19708 4072
rect 19760 4060 19766 4072
rect 19760 4032 21036 4060
rect 19760 4020 19766 4032
rect 21008 3992 21036 4032
rect 21358 4020 21364 4072
rect 21416 4060 21422 4072
rect 21910 4060 21916 4072
rect 21416 4032 21916 4060
rect 21416 4020 21422 4032
rect 21910 4020 21916 4032
rect 21968 4060 21974 4072
rect 22373 4063 22431 4069
rect 22373 4060 22385 4063
rect 21968 4032 22385 4060
rect 21968 4020 21974 4032
rect 22373 4029 22385 4032
rect 22419 4029 22431 4063
rect 22373 4023 22431 4029
rect 23293 4063 23351 4069
rect 23293 4029 23305 4063
rect 23339 4060 23351 4063
rect 23382 4060 23388 4072
rect 23339 4032 23388 4060
rect 23339 4029 23351 4032
rect 23293 4023 23351 4029
rect 23382 4020 23388 4032
rect 23440 4020 23446 4072
rect 23477 4063 23535 4069
rect 23477 4029 23489 4063
rect 23523 4029 23535 4063
rect 23477 4023 23535 4029
rect 22002 3992 22008 4004
rect 21008 3964 22008 3992
rect 22002 3952 22008 3964
rect 22060 3992 22066 4004
rect 23492 3992 23520 4023
rect 23750 4020 23756 4072
rect 23808 4020 23814 4072
rect 25225 4063 25283 4069
rect 25225 4029 25237 4063
rect 25271 4060 25283 4063
rect 25593 4063 25651 4069
rect 25593 4060 25605 4063
rect 25271 4032 25605 4060
rect 25271 4029 25283 4032
rect 25225 4023 25283 4029
rect 25593 4029 25605 4032
rect 25639 4029 25651 4063
rect 25593 4023 25651 4029
rect 26421 4063 26479 4069
rect 26421 4029 26433 4063
rect 26467 4060 26479 4063
rect 26896 4060 26924 4100
rect 26467 4032 26924 4060
rect 26973 4063 27031 4069
rect 26467 4029 26479 4032
rect 26421 4023 26479 4029
rect 26973 4029 26985 4063
rect 27019 4060 27031 4063
rect 27019 4032 27108 4060
rect 27019 4029 27031 4032
rect 26973 4023 27031 4029
rect 22060 3964 23520 3992
rect 22060 3952 22066 3964
rect 21358 3884 21364 3936
rect 21416 3924 21422 3936
rect 21453 3927 21511 3933
rect 21453 3924 21465 3927
rect 21416 3896 21465 3924
rect 21416 3884 21422 3896
rect 21453 3893 21465 3896
rect 21499 3893 21511 3927
rect 21453 3887 21511 3893
rect 21542 3884 21548 3936
rect 21600 3924 21606 3936
rect 21821 3927 21879 3933
rect 21821 3924 21833 3927
rect 21600 3896 21833 3924
rect 21600 3884 21606 3896
rect 21821 3893 21833 3896
rect 21867 3893 21879 3927
rect 21821 3887 21879 3893
rect 22830 3884 22836 3936
rect 22888 3884 22894 3936
rect 23290 3884 23296 3936
rect 23348 3924 23354 3936
rect 25240 3924 25268 4023
rect 23348 3896 25268 3924
rect 23348 3884 23354 3896
rect 25958 3884 25964 3936
rect 26016 3924 26022 3936
rect 26237 3927 26295 3933
rect 26237 3924 26249 3927
rect 26016 3896 26249 3924
rect 26016 3884 26022 3896
rect 26237 3893 26249 3896
rect 26283 3893 26295 3927
rect 27080 3924 27108 4032
rect 28718 4020 28724 4072
rect 28776 4020 28782 4072
rect 27982 3924 27988 3936
rect 27080 3896 27988 3924
rect 26237 3887 26295 3893
rect 27982 3884 27988 3896
rect 28040 3884 28046 3936
rect 1104 3834 58880 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 58880 3834
rect 1104 3760 58880 3782
rect 23385 3723 23443 3729
rect 23385 3689 23397 3723
rect 23431 3720 23443 3723
rect 24670 3720 24676 3732
rect 23431 3692 24676 3720
rect 23431 3689 23443 3692
rect 23385 3683 23443 3689
rect 24670 3680 24676 3692
rect 24728 3680 24734 3732
rect 25314 3680 25320 3732
rect 25372 3680 25378 3732
rect 25774 3680 25780 3732
rect 25832 3720 25838 3732
rect 26510 3720 26516 3732
rect 25832 3692 26516 3720
rect 25832 3680 25838 3692
rect 26510 3680 26516 3692
rect 26568 3720 26574 3732
rect 26568 3692 27568 3720
rect 26568 3680 26574 3692
rect 23474 3612 23480 3664
rect 23532 3612 23538 3664
rect 25792 3652 25820 3680
rect 23584 3624 25820 3652
rect 27540 3652 27568 3692
rect 27890 3680 27896 3732
rect 27948 3720 27954 3732
rect 27985 3723 28043 3729
rect 27985 3720 27997 3723
rect 27948 3692 27997 3720
rect 27948 3680 27954 3692
rect 27985 3689 27997 3692
rect 28031 3689 28043 3723
rect 27985 3683 28043 3689
rect 30742 3680 30748 3732
rect 30800 3680 30806 3732
rect 31386 3680 31392 3732
rect 31444 3720 31450 3732
rect 32401 3723 32459 3729
rect 32401 3720 32413 3723
rect 31444 3692 32413 3720
rect 31444 3680 31450 3692
rect 32401 3689 32413 3692
rect 32447 3689 32459 3723
rect 32401 3683 32459 3689
rect 30760 3652 30788 3680
rect 27540 3624 30788 3652
rect 19702 3544 19708 3596
rect 19760 3544 19766 3596
rect 23584 3584 23612 3624
rect 23308 3556 23612 3584
rect 22373 3519 22431 3525
rect 22373 3516 22385 3519
rect 22112 3488 22385 3516
rect 19978 3408 19984 3460
rect 20036 3408 20042 3460
rect 20714 3408 20720 3460
rect 20772 3408 20778 3460
rect 21818 3448 21824 3460
rect 21468 3420 21824 3448
rect 21468 3389 21496 3420
rect 21818 3408 21824 3420
rect 21876 3448 21882 3460
rect 22112 3457 22140 3488
rect 22373 3485 22385 3488
rect 22419 3485 22431 3519
rect 22373 3479 22431 3485
rect 23017 3519 23075 3525
rect 23017 3485 23029 3519
rect 23063 3516 23075 3519
rect 23201 3519 23259 3525
rect 23201 3516 23213 3519
rect 23063 3488 23213 3516
rect 23063 3485 23075 3488
rect 23017 3479 23075 3485
rect 23201 3485 23213 3488
rect 23247 3485 23259 3519
rect 23308 3516 23336 3556
rect 23934 3544 23940 3596
rect 23992 3584 23998 3596
rect 24762 3584 24768 3596
rect 23992 3556 24768 3584
rect 23992 3544 23998 3556
rect 24762 3544 24768 3556
rect 24820 3584 24826 3596
rect 26237 3587 26295 3593
rect 26237 3584 26249 3587
rect 24820 3556 26249 3584
rect 24820 3544 24826 3556
rect 26237 3553 26249 3556
rect 26283 3584 26295 3587
rect 28074 3584 28080 3596
rect 26283 3556 28080 3584
rect 26283 3553 26295 3556
rect 26237 3547 26295 3553
rect 28074 3544 28080 3556
rect 28132 3544 28138 3596
rect 30374 3544 30380 3596
rect 30432 3584 30438 3596
rect 30653 3587 30711 3593
rect 30653 3584 30665 3587
rect 30432 3556 30665 3584
rect 30432 3544 30438 3556
rect 30653 3553 30665 3556
rect 30699 3584 30711 3587
rect 31478 3584 31484 3596
rect 30699 3556 31484 3584
rect 30699 3553 30711 3556
rect 30653 3547 30711 3553
rect 31478 3544 31484 3556
rect 31536 3544 31542 3596
rect 23382 3516 23388 3528
rect 23308 3488 23388 3516
rect 23201 3479 23259 3485
rect 23382 3476 23388 3488
rect 23440 3476 23446 3528
rect 23477 3519 23535 3525
rect 23477 3485 23489 3519
rect 23523 3485 23535 3519
rect 23477 3479 23535 3485
rect 23661 3519 23719 3525
rect 23661 3485 23673 3519
rect 23707 3516 23719 3519
rect 24673 3519 24731 3525
rect 24673 3516 24685 3519
rect 23707 3488 24685 3516
rect 23707 3485 23719 3488
rect 23661 3479 23719 3485
rect 24673 3485 24685 3488
rect 24719 3516 24731 3519
rect 25682 3516 25688 3528
rect 24719 3488 25688 3516
rect 24719 3485 24731 3488
rect 24673 3479 24731 3485
rect 22097 3451 22155 3457
rect 22097 3448 22109 3451
rect 21876 3420 22109 3448
rect 21876 3408 21882 3420
rect 22097 3417 22109 3420
rect 22143 3448 22155 3451
rect 22281 3451 22339 3457
rect 22143 3420 22197 3448
rect 22143 3417 22155 3420
rect 22097 3411 22155 3417
rect 22281 3417 22293 3451
rect 22327 3448 22339 3451
rect 22922 3448 22928 3460
rect 22327 3420 22928 3448
rect 22327 3417 22339 3420
rect 22281 3411 22339 3417
rect 22922 3408 22928 3420
rect 22980 3448 22986 3460
rect 23492 3448 23520 3479
rect 22980 3420 23520 3448
rect 22980 3408 22986 3420
rect 21453 3383 21511 3389
rect 21453 3349 21465 3383
rect 21499 3349 21511 3383
rect 21453 3343 21511 3349
rect 21910 3340 21916 3392
rect 21968 3340 21974 3392
rect 22646 3340 22652 3392
rect 22704 3380 22710 3392
rect 23290 3380 23296 3392
rect 22704 3352 23296 3380
rect 22704 3340 22710 3352
rect 23290 3340 23296 3352
rect 23348 3340 23354 3392
rect 23382 3340 23388 3392
rect 23440 3380 23446 3392
rect 23676 3380 23704 3479
rect 25682 3476 25688 3488
rect 25740 3476 25746 3528
rect 25774 3476 25780 3528
rect 25832 3476 25838 3528
rect 25958 3476 25964 3528
rect 26016 3476 26022 3528
rect 28629 3519 28687 3525
rect 28629 3485 28641 3519
rect 28675 3516 28687 3519
rect 29362 3516 29368 3528
rect 28675 3488 29368 3516
rect 28675 3485 28687 3488
rect 28629 3479 28687 3485
rect 29362 3476 29368 3488
rect 29420 3476 29426 3528
rect 30282 3476 30288 3528
rect 30340 3476 30346 3528
rect 25869 3451 25927 3457
rect 25869 3417 25881 3451
rect 25915 3448 25927 3451
rect 26513 3451 26571 3457
rect 26513 3448 26525 3451
rect 25915 3420 26525 3448
rect 25915 3417 25927 3420
rect 25869 3411 25927 3417
rect 26513 3417 26525 3420
rect 26559 3417 26571 3451
rect 27798 3448 27804 3460
rect 27738 3420 27804 3448
rect 26513 3411 26571 3417
rect 27798 3408 27804 3420
rect 27856 3448 27862 3460
rect 28810 3448 28816 3460
rect 27856 3420 28816 3448
rect 27856 3408 27862 3420
rect 28810 3408 28816 3420
rect 28868 3408 28874 3460
rect 30558 3408 30564 3460
rect 30616 3448 30622 3460
rect 30929 3451 30987 3457
rect 30929 3448 30941 3451
rect 30616 3420 30941 3448
rect 30616 3408 30622 3420
rect 30929 3417 30941 3420
rect 30975 3417 30987 3451
rect 32306 3448 32312 3460
rect 32154 3420 32312 3448
rect 30929 3411 30987 3417
rect 32306 3408 32312 3420
rect 32364 3448 32370 3460
rect 32858 3448 32864 3460
rect 32364 3420 32864 3448
rect 32364 3408 32370 3420
rect 32858 3408 32864 3420
rect 32916 3408 32922 3460
rect 23440 3352 23704 3380
rect 23440 3340 23446 3352
rect 28350 3340 28356 3392
rect 28408 3380 28414 3392
rect 28445 3383 28503 3389
rect 28445 3380 28457 3383
rect 28408 3352 28457 3380
rect 28408 3340 28414 3352
rect 28445 3349 28457 3352
rect 28491 3349 28503 3383
rect 28445 3343 28503 3349
rect 30469 3383 30527 3389
rect 30469 3349 30481 3383
rect 30515 3380 30527 3383
rect 32398 3380 32404 3392
rect 30515 3352 32404 3380
rect 30515 3349 30527 3352
rect 30469 3343 30527 3349
rect 32398 3340 32404 3352
rect 32456 3340 32462 3392
rect 1104 3290 58880 3312
rect 1104 3238 4874 3290
rect 4926 3238 4938 3290
rect 4990 3238 5002 3290
rect 5054 3238 5066 3290
rect 5118 3238 5130 3290
rect 5182 3238 35594 3290
rect 35646 3238 35658 3290
rect 35710 3238 35722 3290
rect 35774 3238 35786 3290
rect 35838 3238 35850 3290
rect 35902 3238 58880 3290
rect 1104 3216 58880 3238
rect 19978 3136 19984 3188
rect 20036 3176 20042 3188
rect 20809 3179 20867 3185
rect 20809 3176 20821 3179
rect 20036 3148 20821 3176
rect 20036 3136 20042 3148
rect 20809 3145 20821 3148
rect 20855 3145 20867 3179
rect 20809 3139 20867 3145
rect 22005 3179 22063 3185
rect 22005 3145 22017 3179
rect 22051 3176 22063 3179
rect 22186 3176 22192 3188
rect 22051 3148 22192 3176
rect 22051 3145 22063 3148
rect 22005 3139 22063 3145
rect 22186 3136 22192 3148
rect 22244 3136 22250 3188
rect 22554 3136 22560 3188
rect 22612 3176 22618 3188
rect 22925 3179 22983 3185
rect 22925 3176 22937 3179
rect 22612 3148 22937 3176
rect 22612 3136 22618 3148
rect 22925 3145 22937 3148
rect 22971 3145 22983 3179
rect 22925 3139 22983 3145
rect 23290 3136 23296 3188
rect 23348 3176 23354 3188
rect 23385 3179 23443 3185
rect 23385 3176 23397 3179
rect 23348 3148 23397 3176
rect 23348 3136 23354 3148
rect 23385 3145 23397 3148
rect 23431 3145 23443 3179
rect 23385 3139 23443 3145
rect 23750 3136 23756 3188
rect 23808 3136 23814 3188
rect 25682 3136 25688 3188
rect 25740 3136 25746 3188
rect 28074 3136 28080 3188
rect 28132 3176 28138 3188
rect 31757 3179 31815 3185
rect 28132 3148 30052 3176
rect 28132 3136 28138 3148
rect 22097 3111 22155 3117
rect 22097 3077 22109 3111
rect 22143 3108 22155 3111
rect 22646 3108 22652 3120
rect 22143 3080 22652 3108
rect 22143 3077 22155 3080
rect 22097 3071 22155 3077
rect 22646 3068 22652 3080
rect 22704 3068 22710 3120
rect 22830 3068 22836 3120
rect 22888 3108 22894 3120
rect 24213 3111 24271 3117
rect 24213 3108 24225 3111
rect 22888 3080 24225 3108
rect 22888 3068 22894 3080
rect 24213 3077 24225 3080
rect 24259 3077 24271 3111
rect 26050 3108 26056 3120
rect 25438 3080 26056 3108
rect 24213 3071 24271 3077
rect 26050 3068 26056 3080
rect 26108 3068 26114 3120
rect 20993 3043 21051 3049
rect 20993 3009 21005 3043
rect 21039 3040 21051 3043
rect 21910 3040 21916 3052
rect 21039 3012 21916 3040
rect 21039 3009 21051 3012
rect 20993 3003 21051 3009
rect 21910 3000 21916 3012
rect 21968 3000 21974 3052
rect 22189 3043 22247 3049
rect 22189 3009 22201 3043
rect 22235 3040 22247 3043
rect 22235 3012 22968 3040
rect 22235 3009 22247 3012
rect 22189 3003 22247 3009
rect 22940 2984 22968 3012
rect 23934 3000 23940 3052
rect 23992 3000 23998 3052
rect 28092 3049 28120 3136
rect 28350 3068 28356 3120
rect 28408 3068 28414 3120
rect 28810 3068 28816 3120
rect 28868 3068 28874 3120
rect 30024 3108 30052 3148
rect 31757 3145 31769 3179
rect 31803 3176 31815 3179
rect 32674 3176 32680 3188
rect 31803 3148 32680 3176
rect 31803 3145 31815 3148
rect 31757 3139 31815 3145
rect 32674 3136 32680 3148
rect 32732 3136 32738 3188
rect 33778 3136 33784 3188
rect 33836 3176 33842 3188
rect 33873 3179 33931 3185
rect 33873 3176 33885 3179
rect 33836 3148 33885 3176
rect 33836 3136 33842 3148
rect 33873 3145 33885 3148
rect 33919 3145 33931 3179
rect 33873 3139 33931 3145
rect 30374 3108 30380 3120
rect 30024 3080 30380 3108
rect 30024 3049 30052 3080
rect 30374 3068 30380 3080
rect 30432 3068 30438 3120
rect 32306 3108 32312 3120
rect 31510 3080 32312 3108
rect 32306 3068 32312 3080
rect 32364 3068 32370 3120
rect 32398 3068 32404 3120
rect 32456 3068 32462 3120
rect 32858 3068 32864 3120
rect 32916 3068 32922 3120
rect 28077 3043 28135 3049
rect 28077 3009 28089 3043
rect 28123 3009 28135 3043
rect 28077 3003 28135 3009
rect 30009 3043 30067 3049
rect 30009 3009 30021 3043
rect 30055 3009 30067 3043
rect 30009 3003 30067 3009
rect 34333 3043 34391 3049
rect 34333 3009 34345 3043
rect 34379 3040 34391 3043
rect 34425 3043 34483 3049
rect 34425 3040 34437 3043
rect 34379 3012 34437 3040
rect 34379 3009 34391 3012
rect 34333 3003 34391 3009
rect 34425 3009 34437 3012
rect 34471 3009 34483 3043
rect 34425 3003 34483 3009
rect 35069 3043 35127 3049
rect 35069 3009 35081 3043
rect 35115 3009 35127 3043
rect 35069 3003 35127 3009
rect 35253 3043 35311 3049
rect 35253 3009 35265 3043
rect 35299 3040 35311 3043
rect 35342 3040 35348 3052
rect 35299 3012 35348 3040
rect 35299 3009 35311 3012
rect 35253 3003 35311 3009
rect 21174 2932 21180 2984
rect 21232 2932 21238 2984
rect 21269 2975 21327 2981
rect 21269 2941 21281 2975
rect 21315 2972 21327 2975
rect 21542 2972 21548 2984
rect 21315 2944 21548 2972
rect 21315 2941 21327 2944
rect 21269 2935 21327 2941
rect 21542 2932 21548 2944
rect 21600 2932 21606 2984
rect 21818 2932 21824 2984
rect 21876 2972 21882 2984
rect 22281 2975 22339 2981
rect 22281 2972 22293 2975
rect 21876 2944 22293 2972
rect 21876 2932 21882 2944
rect 22281 2941 22293 2944
rect 22327 2941 22339 2975
rect 22281 2935 22339 2941
rect 22557 2975 22615 2981
rect 22557 2941 22569 2975
rect 22603 2941 22615 2975
rect 22557 2935 22615 2941
rect 22766 2975 22824 2981
rect 22766 2941 22778 2975
rect 22812 2972 22824 2975
rect 22922 2972 22928 2984
rect 22812 2944 22928 2972
rect 22812 2941 22824 2944
rect 22766 2935 22824 2941
rect 21192 2904 21220 2932
rect 21913 2907 21971 2913
rect 21913 2904 21925 2907
rect 21192 2876 21925 2904
rect 21913 2873 21925 2876
rect 21959 2873 21971 2907
rect 21913 2867 21971 2873
rect 22186 2864 22192 2916
rect 22244 2904 22250 2916
rect 22572 2904 22600 2935
rect 22922 2932 22928 2944
rect 22980 2972 22986 2984
rect 23109 2975 23167 2981
rect 23109 2972 23121 2975
rect 22980 2944 23121 2972
rect 22980 2932 22986 2944
rect 23109 2941 23121 2944
rect 23155 2941 23167 2975
rect 23109 2935 23167 2941
rect 23290 2932 23296 2984
rect 23348 2932 23354 2984
rect 28994 2932 29000 2984
rect 29052 2972 29058 2984
rect 30285 2975 30343 2981
rect 30285 2972 30297 2975
rect 29052 2944 30297 2972
rect 29052 2932 29058 2944
rect 30285 2941 30297 2944
rect 30331 2941 30343 2975
rect 30285 2935 30343 2941
rect 31478 2932 31484 2984
rect 31536 2972 31542 2984
rect 32125 2975 32183 2981
rect 32125 2972 32137 2975
rect 31536 2944 32137 2972
rect 31536 2932 31542 2944
rect 32125 2941 32137 2944
rect 32171 2941 32183 2975
rect 35084 2972 35112 3003
rect 35342 3000 35348 3012
rect 35400 3000 35406 3052
rect 36173 3043 36231 3049
rect 36173 3009 36185 3043
rect 36219 3040 36231 3043
rect 36265 3043 36323 3049
rect 36265 3040 36277 3043
rect 36219 3012 36277 3040
rect 36219 3009 36231 3012
rect 36173 3003 36231 3009
rect 36265 3009 36277 3012
rect 36311 3009 36323 3043
rect 36265 3003 36323 3009
rect 36817 3043 36875 3049
rect 36817 3009 36829 3043
rect 36863 3040 36875 3043
rect 36909 3043 36967 3049
rect 36909 3040 36921 3043
rect 36863 3012 36921 3040
rect 36863 3009 36875 3012
rect 36817 3003 36875 3009
rect 36909 3009 36921 3012
rect 36955 3009 36967 3043
rect 36909 3003 36967 3009
rect 37274 3000 37280 3052
rect 37332 3000 37338 3052
rect 38105 3043 38163 3049
rect 38105 3009 38117 3043
rect 38151 3040 38163 3043
rect 38197 3043 38255 3049
rect 38197 3040 38209 3043
rect 38151 3012 38209 3040
rect 38151 3009 38163 3012
rect 38105 3003 38163 3009
rect 38197 3009 38209 3012
rect 38243 3009 38255 3043
rect 38197 3003 38255 3009
rect 38749 3043 38807 3049
rect 38749 3009 38761 3043
rect 38795 3040 38807 3043
rect 38841 3043 38899 3049
rect 38841 3040 38853 3043
rect 38795 3012 38853 3040
rect 38795 3009 38807 3012
rect 38749 3003 38807 3009
rect 38841 3009 38853 3012
rect 38887 3009 38899 3043
rect 38841 3003 38899 3009
rect 39393 3043 39451 3049
rect 39393 3009 39405 3043
rect 39439 3040 39451 3043
rect 39485 3043 39543 3049
rect 39485 3040 39497 3043
rect 39439 3012 39497 3040
rect 39439 3009 39451 3012
rect 39393 3003 39451 3009
rect 39485 3009 39497 3012
rect 39531 3009 39543 3043
rect 39485 3003 39543 3009
rect 40037 3043 40095 3049
rect 40037 3009 40049 3043
rect 40083 3040 40095 3043
rect 40129 3043 40187 3049
rect 40129 3040 40141 3043
rect 40083 3012 40141 3040
rect 40083 3009 40095 3012
rect 40037 3003 40095 3009
rect 40129 3009 40141 3012
rect 40175 3009 40187 3043
rect 40129 3003 40187 3009
rect 40681 3043 40739 3049
rect 40681 3009 40693 3043
rect 40727 3040 40739 3043
rect 40773 3043 40831 3049
rect 40773 3040 40785 3043
rect 40727 3012 40785 3040
rect 40727 3009 40739 3012
rect 40681 3003 40739 3009
rect 40773 3009 40785 3012
rect 40819 3009 40831 3043
rect 40773 3003 40831 3009
rect 41325 3043 41383 3049
rect 41325 3009 41337 3043
rect 41371 3040 41383 3043
rect 41417 3043 41475 3049
rect 41417 3040 41429 3043
rect 41371 3012 41429 3040
rect 41371 3009 41383 3012
rect 41325 3003 41383 3009
rect 41417 3009 41429 3012
rect 41463 3009 41475 3043
rect 41417 3003 41475 3009
rect 41969 3043 42027 3049
rect 41969 3009 41981 3043
rect 42015 3040 42027 3043
rect 42061 3043 42119 3049
rect 42061 3040 42073 3043
rect 42015 3012 42073 3040
rect 42015 3009 42027 3012
rect 41969 3003 42027 3009
rect 42061 3009 42073 3012
rect 42107 3009 42119 3043
rect 42061 3003 42119 3009
rect 42426 3000 42432 3052
rect 42484 3000 42490 3052
rect 43257 3043 43315 3049
rect 43257 3009 43269 3043
rect 43303 3040 43315 3043
rect 43349 3043 43407 3049
rect 43349 3040 43361 3043
rect 43303 3012 43361 3040
rect 43303 3009 43315 3012
rect 43257 3003 43315 3009
rect 43349 3009 43361 3012
rect 43395 3009 43407 3043
rect 43349 3003 43407 3009
rect 43622 3000 43628 3052
rect 43680 3000 43686 3052
rect 44361 3043 44419 3049
rect 44361 3009 44373 3043
rect 44407 3009 44419 3043
rect 44361 3003 44419 3009
rect 44729 3043 44787 3049
rect 44729 3009 44741 3043
rect 44775 3040 44787 3043
rect 45097 3043 45155 3049
rect 45097 3040 45109 3043
rect 44775 3012 45109 3040
rect 44775 3009 44787 3012
rect 44729 3003 44787 3009
rect 45097 3009 45109 3012
rect 45143 3009 45155 3043
rect 45097 3003 45155 3009
rect 35621 2975 35679 2981
rect 35621 2972 35633 2975
rect 35084 2944 35633 2972
rect 32125 2935 32183 2941
rect 35621 2941 35633 2944
rect 35667 2941 35679 2975
rect 44376 2972 44404 3003
rect 44821 2975 44879 2981
rect 44821 2972 44833 2975
rect 44376 2944 44833 2972
rect 35621 2935 35679 2941
rect 44821 2941 44833 2944
rect 44867 2941 44879 2975
rect 44821 2935 44879 2941
rect 23382 2904 23388 2916
rect 22244 2876 23388 2904
rect 22244 2864 22250 2876
rect 23382 2864 23388 2876
rect 23440 2864 23446 2916
rect 29825 2839 29883 2845
rect 29825 2805 29837 2839
rect 29871 2836 29883 2839
rect 30650 2836 30656 2848
rect 29871 2808 30656 2836
rect 29871 2805 29883 2808
rect 29825 2799 29883 2805
rect 30650 2796 30656 2808
rect 30708 2796 30714 2848
rect 34146 2796 34152 2848
rect 34204 2836 34210 2848
rect 34609 2839 34667 2845
rect 34609 2836 34621 2839
rect 34204 2808 34621 2836
rect 34204 2796 34210 2808
rect 34609 2805 34621 2808
rect 34655 2805 34667 2839
rect 34609 2799 34667 2805
rect 34790 2796 34796 2848
rect 34848 2836 34854 2848
rect 34885 2839 34943 2845
rect 34885 2836 34897 2839
rect 34848 2808 34897 2836
rect 34848 2796 34854 2808
rect 34885 2805 34897 2808
rect 34931 2805 34943 2839
rect 34885 2799 34943 2805
rect 35434 2796 35440 2848
rect 35492 2796 35498 2848
rect 35989 2839 36047 2845
rect 35989 2805 36001 2839
rect 36035 2836 36047 2839
rect 36078 2836 36084 2848
rect 36035 2808 36084 2836
rect 36035 2805 36047 2808
rect 35989 2799 36047 2805
rect 36078 2796 36084 2808
rect 36136 2796 36142 2848
rect 36633 2839 36691 2845
rect 36633 2805 36645 2839
rect 36679 2836 36691 2839
rect 36722 2836 36728 2848
rect 36679 2808 36728 2836
rect 36679 2805 36691 2808
rect 36633 2799 36691 2805
rect 36722 2796 36728 2808
rect 36780 2796 36786 2848
rect 37366 2796 37372 2848
rect 37424 2836 37430 2848
rect 37461 2839 37519 2845
rect 37461 2836 37473 2839
rect 37424 2808 37473 2836
rect 37424 2796 37430 2808
rect 37461 2805 37473 2808
rect 37507 2805 37519 2839
rect 37461 2799 37519 2805
rect 37921 2839 37979 2845
rect 37921 2805 37933 2839
rect 37967 2836 37979 2839
rect 38010 2836 38016 2848
rect 37967 2808 38016 2836
rect 37967 2805 37979 2808
rect 37921 2799 37979 2805
rect 38010 2796 38016 2808
rect 38068 2796 38074 2848
rect 38565 2839 38623 2845
rect 38565 2805 38577 2839
rect 38611 2836 38623 2839
rect 38654 2836 38660 2848
rect 38611 2808 38660 2836
rect 38611 2805 38623 2808
rect 38565 2799 38623 2805
rect 38654 2796 38660 2808
rect 38712 2796 38718 2848
rect 39209 2839 39267 2845
rect 39209 2805 39221 2839
rect 39255 2836 39267 2839
rect 39298 2836 39304 2848
rect 39255 2808 39304 2836
rect 39255 2805 39267 2808
rect 39209 2799 39267 2805
rect 39298 2796 39304 2808
rect 39356 2796 39362 2848
rect 39853 2839 39911 2845
rect 39853 2805 39865 2839
rect 39899 2836 39911 2839
rect 39942 2836 39948 2848
rect 39899 2808 39948 2836
rect 39899 2805 39911 2808
rect 39853 2799 39911 2805
rect 39942 2796 39948 2808
rect 40000 2796 40006 2848
rect 40497 2839 40555 2845
rect 40497 2805 40509 2839
rect 40543 2836 40555 2839
rect 40586 2836 40592 2848
rect 40543 2808 40592 2836
rect 40543 2805 40555 2808
rect 40497 2799 40555 2805
rect 40586 2796 40592 2808
rect 40644 2796 40650 2848
rect 41141 2839 41199 2845
rect 41141 2805 41153 2839
rect 41187 2836 41199 2839
rect 41230 2836 41236 2848
rect 41187 2808 41236 2836
rect 41187 2805 41199 2808
rect 41141 2799 41199 2805
rect 41230 2796 41236 2808
rect 41288 2796 41294 2848
rect 41785 2839 41843 2845
rect 41785 2805 41797 2839
rect 41831 2836 41843 2839
rect 41874 2836 41880 2848
rect 41831 2808 41880 2836
rect 41831 2805 41843 2808
rect 41785 2799 41843 2805
rect 41874 2796 41880 2808
rect 41932 2796 41938 2848
rect 42518 2796 42524 2848
rect 42576 2836 42582 2848
rect 42613 2839 42671 2845
rect 42613 2836 42625 2839
rect 42576 2808 42625 2836
rect 42576 2796 42582 2808
rect 42613 2805 42625 2808
rect 42659 2805 42671 2839
rect 42613 2799 42671 2805
rect 43073 2839 43131 2845
rect 43073 2805 43085 2839
rect 43119 2836 43131 2839
rect 43162 2836 43168 2848
rect 43119 2808 43168 2836
rect 43119 2805 43131 2808
rect 43073 2799 43131 2805
rect 43162 2796 43168 2808
rect 43220 2796 43226 2848
rect 43806 2796 43812 2848
rect 43864 2796 43870 2848
rect 44177 2839 44235 2845
rect 44177 2805 44189 2839
rect 44223 2836 44235 2839
rect 44450 2836 44456 2848
rect 44223 2808 44456 2836
rect 44223 2805 44235 2808
rect 44177 2799 44235 2805
rect 44450 2796 44456 2808
rect 44508 2796 44514 2848
rect 44545 2839 44603 2845
rect 44545 2805 44557 2839
rect 44591 2836 44603 2839
rect 45094 2836 45100 2848
rect 44591 2808 45100 2836
rect 44591 2805 44603 2808
rect 44545 2799 44603 2805
rect 45094 2796 45100 2808
rect 45152 2796 45158 2848
rect 1104 2746 58880 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 58880 2746
rect 1104 2672 58880 2694
rect 19334 2592 19340 2644
rect 19392 2632 19398 2644
rect 19429 2635 19487 2641
rect 19429 2632 19441 2635
rect 19392 2604 19441 2632
rect 19392 2592 19398 2604
rect 19429 2601 19441 2604
rect 19475 2601 19487 2635
rect 19429 2595 19487 2601
rect 28905 2635 28963 2641
rect 28905 2601 28917 2635
rect 28951 2632 28963 2635
rect 28994 2632 29000 2644
rect 28951 2604 29000 2632
rect 28951 2601 28963 2604
rect 28905 2595 28963 2601
rect 28994 2592 29000 2604
rect 29052 2592 29058 2644
rect 29362 2592 29368 2644
rect 29420 2632 29426 2644
rect 30098 2632 30104 2644
rect 29420 2604 30104 2632
rect 29420 2592 29426 2604
rect 30098 2592 30104 2604
rect 30156 2592 30162 2644
rect 30282 2592 30288 2644
rect 30340 2632 30346 2644
rect 31021 2635 31079 2641
rect 31021 2632 31033 2635
rect 30340 2604 31033 2632
rect 30340 2592 30346 2604
rect 31021 2601 31033 2604
rect 31067 2601 31079 2635
rect 31021 2595 31079 2601
rect 22554 2524 22560 2576
rect 22612 2564 22618 2576
rect 22833 2567 22891 2573
rect 22833 2564 22845 2567
rect 22612 2536 22845 2564
rect 22612 2524 22618 2536
rect 22833 2533 22845 2536
rect 22879 2533 22891 2567
rect 22833 2527 22891 2533
rect 29733 2567 29791 2573
rect 29733 2533 29745 2567
rect 29779 2564 29791 2567
rect 30374 2564 30380 2576
rect 29779 2536 30380 2564
rect 29779 2533 29791 2536
rect 29733 2527 29791 2533
rect 30374 2524 30380 2536
rect 30432 2524 30438 2576
rect 30745 2567 30803 2573
rect 30745 2533 30757 2567
rect 30791 2533 30803 2567
rect 30745 2527 30803 2533
rect 21818 2456 21824 2508
rect 21876 2496 21882 2508
rect 22649 2499 22707 2505
rect 21876 2468 22324 2496
rect 21876 2456 21882 2468
rect 19613 2431 19671 2437
rect 19613 2428 19625 2431
rect 19352 2400 19625 2428
rect 19352 2304 19380 2400
rect 19613 2397 19625 2400
rect 19659 2397 19671 2431
rect 19613 2391 19671 2397
rect 20993 2431 21051 2437
rect 20993 2397 21005 2431
rect 21039 2397 21051 2431
rect 20993 2391 21051 2397
rect 21637 2431 21695 2437
rect 21637 2397 21649 2431
rect 21683 2428 21695 2431
rect 21836 2428 21864 2456
rect 21683 2400 21864 2428
rect 21683 2397 21695 2400
rect 21637 2391 21695 2397
rect 21008 2360 21036 2391
rect 22186 2388 22192 2440
rect 22244 2388 22250 2440
rect 22296 2437 22324 2468
rect 22649 2465 22661 2499
rect 22695 2496 22707 2499
rect 23290 2496 23296 2508
rect 22695 2468 23296 2496
rect 22695 2465 22707 2468
rect 22649 2459 22707 2465
rect 23290 2456 23296 2468
rect 23348 2456 23354 2508
rect 28353 2499 28411 2505
rect 28353 2465 28365 2499
rect 28399 2496 28411 2499
rect 28994 2496 29000 2508
rect 28399 2468 29000 2496
rect 28399 2465 28411 2468
rect 28353 2459 28411 2465
rect 22281 2431 22339 2437
rect 22281 2397 22293 2431
rect 22327 2397 22339 2431
rect 22281 2391 22339 2397
rect 23017 2431 23075 2437
rect 23017 2397 23029 2431
rect 23063 2397 23075 2431
rect 23017 2391 23075 2397
rect 21358 2360 21364 2372
rect 21008 2332 21364 2360
rect 21358 2320 21364 2332
rect 21416 2360 21422 2372
rect 22373 2363 22431 2369
rect 22373 2360 22385 2363
rect 21416 2332 22385 2360
rect 21416 2320 21422 2332
rect 22373 2329 22385 2332
rect 22419 2329 22431 2363
rect 22373 2323 22431 2329
rect 22465 2363 22523 2369
rect 22465 2329 22477 2363
rect 22511 2360 22523 2363
rect 22646 2360 22652 2372
rect 22511 2332 22652 2360
rect 22511 2329 22523 2332
rect 22465 2323 22523 2329
rect 22646 2320 22652 2332
rect 22704 2360 22710 2372
rect 23032 2360 23060 2391
rect 23382 2388 23388 2440
rect 23440 2428 23446 2440
rect 28460 2437 28488 2468
rect 28994 2456 29000 2468
rect 29052 2456 29058 2508
rect 30760 2496 30788 2527
rect 31481 2499 31539 2505
rect 31481 2496 31493 2499
rect 29564 2468 30788 2496
rect 30944 2468 31493 2496
rect 29564 2437 29592 2468
rect 23569 2431 23627 2437
rect 23569 2428 23581 2431
rect 23440 2400 23581 2428
rect 23440 2388 23446 2400
rect 23569 2397 23581 2400
rect 23615 2397 23627 2431
rect 23569 2391 23627 2397
rect 28445 2431 28503 2437
rect 28445 2397 28457 2431
rect 28491 2428 28503 2431
rect 28721 2431 28779 2437
rect 28491 2400 28525 2428
rect 28491 2397 28503 2400
rect 28445 2391 28503 2397
rect 28721 2397 28733 2431
rect 28767 2397 28779 2431
rect 28721 2391 28779 2397
rect 29181 2431 29239 2437
rect 29181 2397 29193 2431
rect 29227 2428 29239 2431
rect 29549 2431 29607 2437
rect 29227 2400 29261 2428
rect 29227 2397 29239 2400
rect 29181 2391 29239 2397
rect 29549 2397 29561 2431
rect 29595 2397 29607 2431
rect 29549 2391 29607 2397
rect 29825 2431 29883 2437
rect 29825 2397 29837 2431
rect 29871 2397 29883 2431
rect 29825 2391 29883 2397
rect 22704 2332 23060 2360
rect 22704 2320 22710 2332
rect 19334 2252 19340 2304
rect 19392 2252 19398 2304
rect 20622 2252 20628 2304
rect 20680 2292 20686 2304
rect 20809 2295 20867 2301
rect 20809 2292 20821 2295
rect 20680 2264 20821 2292
rect 20680 2252 20686 2264
rect 20809 2261 20821 2264
rect 20855 2261 20867 2295
rect 20809 2255 20867 2261
rect 21266 2252 21272 2304
rect 21324 2292 21330 2304
rect 21453 2295 21511 2301
rect 21453 2292 21465 2295
rect 21324 2264 21465 2292
rect 21324 2252 21330 2264
rect 21453 2261 21465 2264
rect 21499 2261 21511 2295
rect 21453 2255 21511 2261
rect 23198 2252 23204 2304
rect 23256 2292 23262 2304
rect 23385 2295 23443 2301
rect 23385 2292 23397 2295
rect 23256 2264 23397 2292
rect 23256 2252 23262 2264
rect 23385 2261 23397 2264
rect 23431 2261 23443 2295
rect 23385 2255 23443 2261
rect 28629 2295 28687 2301
rect 28629 2261 28641 2295
rect 28675 2292 28687 2295
rect 28736 2292 28764 2391
rect 29089 2363 29147 2369
rect 29089 2329 29101 2363
rect 29135 2360 29147 2363
rect 29196 2360 29224 2391
rect 29638 2360 29644 2372
rect 29135 2332 29644 2360
rect 29135 2329 29147 2332
rect 29089 2323 29147 2329
rect 29638 2320 29644 2332
rect 29696 2320 29702 2372
rect 29840 2292 29868 2391
rect 30098 2388 30104 2440
rect 30156 2388 30162 2440
rect 30282 2388 30288 2440
rect 30340 2388 30346 2440
rect 30484 2437 30512 2468
rect 30469 2431 30527 2437
rect 30469 2397 30481 2431
rect 30515 2397 30527 2431
rect 30469 2391 30527 2397
rect 30653 2431 30711 2437
rect 30653 2397 30665 2431
rect 30699 2428 30711 2431
rect 30742 2428 30748 2440
rect 30699 2400 30748 2428
rect 30699 2397 30711 2400
rect 30653 2391 30711 2397
rect 30742 2388 30748 2400
rect 30800 2388 30806 2440
rect 30944 2437 30972 2468
rect 31481 2465 31493 2468
rect 31527 2465 31539 2499
rect 31481 2459 31539 2465
rect 35342 2456 35348 2508
rect 35400 2456 35406 2508
rect 37274 2456 37280 2508
rect 37332 2456 37338 2508
rect 42426 2456 42432 2508
rect 42484 2456 42490 2508
rect 43622 2456 43628 2508
rect 43680 2456 43686 2508
rect 30929 2431 30987 2437
rect 30929 2428 30941 2431
rect 30852 2400 30941 2428
rect 30852 2360 30880 2400
rect 30929 2397 30941 2400
rect 30975 2397 30987 2431
rect 30929 2391 30987 2397
rect 31205 2431 31263 2437
rect 31205 2397 31217 2431
rect 31251 2428 31263 2431
rect 31251 2400 31285 2428
rect 31251 2397 31263 2400
rect 31205 2391 31263 2397
rect 31220 2360 31248 2391
rect 31297 2363 31355 2369
rect 31297 2360 31309 2363
rect 30300 2332 30880 2360
rect 30944 2332 31309 2360
rect 30300 2304 30328 2332
rect 30944 2304 30972 2332
rect 31297 2329 31309 2332
rect 31343 2329 31355 2363
rect 31297 2323 31355 2329
rect 28675 2264 29868 2292
rect 28675 2261 28687 2264
rect 28629 2255 28687 2261
rect 30282 2252 30288 2304
rect 30340 2252 30346 2304
rect 30926 2252 30932 2304
rect 30984 2252 30990 2304
rect 1104 2202 58880 2224
rect 1104 2150 4874 2202
rect 4926 2150 4938 2202
rect 4990 2150 5002 2202
rect 5054 2150 5066 2202
rect 5118 2150 5130 2202
rect 5182 2150 35594 2202
rect 35646 2150 35658 2202
rect 35710 2150 35722 2202
rect 35774 2150 35786 2202
rect 35838 2150 35850 2202
rect 35902 2150 58880 2202
rect 1104 2128 58880 2150
<< via1 >>
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 22560 37408 22612 37460
rect 23204 37408 23256 37460
rect 26424 37408 26476 37460
rect 28356 37408 28408 37460
rect 31668 37204 31720 37256
rect 23020 37179 23072 37188
rect 23020 37145 23029 37179
rect 23029 37145 23063 37179
rect 23063 37145 23072 37179
rect 23020 37136 23072 37145
rect 24216 37136 24268 37188
rect 29736 37136 29788 37188
rect 4874 36966 4926 37018
rect 4938 36966 4990 37018
rect 5002 36966 5054 37018
rect 5066 36966 5118 37018
rect 5130 36966 5182 37018
rect 35594 36966 35646 37018
rect 35658 36966 35710 37018
rect 35722 36966 35774 37018
rect 35786 36966 35838 37018
rect 35850 36966 35902 37018
rect 24492 36864 24544 36916
rect 25136 36864 25188 36916
rect 25780 36864 25832 36916
rect 27068 36864 27120 36916
rect 27712 36864 27764 36916
rect 29000 36864 29052 36916
rect 29644 36864 29696 36916
rect 30288 36864 30340 36916
rect 30932 36864 30984 36916
rect 31576 36864 31628 36916
rect 32220 36864 32272 36916
rect 32864 36864 32916 36916
rect 33508 36864 33560 36916
rect 34152 36864 34204 36916
rect 34796 36864 34848 36916
rect 35440 36907 35492 36916
rect 35440 36873 35449 36907
rect 35449 36873 35483 36907
rect 35483 36873 35492 36907
rect 35440 36864 35492 36873
rect 36084 36864 36136 36916
rect 36728 36864 36780 36916
rect 37372 36864 37424 36916
rect 38016 36864 38068 36916
rect 38660 36864 38712 36916
rect 39304 36864 39356 36916
rect 39948 36864 40000 36916
rect 40592 36864 40644 36916
rect 41236 36864 41288 36916
rect 41880 36864 41932 36916
rect 42524 36864 42576 36916
rect 43168 36864 43220 36916
rect 43812 36864 43864 36916
rect 44456 36864 44508 36916
rect 45100 36864 45152 36916
rect 45744 36864 45796 36916
rect 46388 36907 46440 36916
rect 46388 36873 46397 36907
rect 46397 36873 46431 36907
rect 46431 36873 46440 36907
rect 46388 36864 46440 36873
rect 47032 36864 47084 36916
rect 47676 36864 47728 36916
rect 25320 36728 25372 36780
rect 32220 36728 32272 36780
rect 35348 36728 35400 36780
rect 37372 36728 37424 36780
rect 42524 36728 42576 36780
rect 46204 36771 46256 36780
rect 46204 36737 46213 36771
rect 46213 36737 46247 36771
rect 46247 36737 46256 36771
rect 46204 36728 46256 36737
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 24216 36363 24268 36372
rect 24216 36329 24225 36363
rect 24225 36329 24259 36363
rect 24259 36329 24268 36363
rect 24216 36320 24268 36329
rect 25320 36363 25372 36372
rect 25320 36329 25329 36363
rect 25329 36329 25363 36363
rect 25363 36329 25372 36363
rect 25320 36320 25372 36329
rect 32220 36363 32272 36372
rect 32220 36329 32229 36363
rect 32229 36329 32263 36363
rect 32263 36329 32272 36363
rect 32220 36320 32272 36329
rect 35348 36320 35400 36372
rect 37372 36363 37424 36372
rect 37372 36329 37381 36363
rect 37381 36329 37415 36363
rect 37415 36329 37424 36363
rect 37372 36320 37424 36329
rect 42524 36363 42576 36372
rect 42524 36329 42533 36363
rect 42533 36329 42567 36363
rect 42567 36329 42576 36363
rect 42524 36320 42576 36329
rect 46204 36363 46256 36372
rect 46204 36329 46213 36363
rect 46213 36329 46247 36363
rect 46247 36329 46256 36363
rect 46204 36320 46256 36329
rect 22100 36116 22152 36168
rect 23296 36048 23348 36100
rect 23572 36048 23624 36100
rect 28816 36091 28868 36100
rect 28816 36057 28825 36091
rect 28825 36057 28859 36091
rect 28859 36057 28868 36091
rect 28816 36048 28868 36057
rect 29552 36023 29604 36032
rect 29552 35989 29561 36023
rect 29561 35989 29595 36023
rect 29595 35989 29604 36023
rect 29552 35980 29604 35989
rect 29736 36091 29788 36100
rect 29736 36057 29745 36091
rect 29745 36057 29779 36091
rect 29779 36057 29788 36091
rect 29736 36048 29788 36057
rect 33324 35980 33376 36032
rect 4874 35878 4926 35930
rect 4938 35878 4990 35930
rect 5002 35878 5054 35930
rect 5066 35878 5118 35930
rect 5130 35878 5182 35930
rect 35594 35878 35646 35930
rect 35658 35878 35710 35930
rect 35722 35878 35774 35930
rect 35786 35878 35838 35930
rect 35850 35878 35902 35930
rect 23020 35776 23072 35828
rect 23296 35819 23348 35828
rect 23296 35785 23305 35819
rect 23305 35785 23339 35819
rect 23339 35785 23348 35819
rect 23296 35776 23348 35785
rect 25228 35776 25280 35828
rect 28816 35776 28868 35828
rect 29736 35776 29788 35828
rect 26700 35708 26752 35760
rect 29276 35708 29328 35760
rect 21916 35640 21968 35692
rect 23572 35683 23624 35692
rect 23572 35649 23581 35683
rect 23581 35649 23615 35683
rect 23615 35649 23624 35683
rect 23572 35640 23624 35649
rect 23664 35683 23716 35692
rect 23664 35649 23673 35683
rect 23673 35649 23707 35683
rect 23707 35649 23716 35683
rect 23664 35640 23716 35649
rect 23756 35683 23808 35692
rect 23756 35649 23765 35683
rect 23765 35649 23799 35683
rect 23799 35649 23808 35683
rect 23756 35640 23808 35649
rect 28816 35683 28868 35692
rect 28816 35649 28850 35683
rect 28850 35649 28868 35683
rect 28816 35640 28868 35649
rect 25044 35615 25096 35624
rect 25044 35581 25053 35615
rect 25053 35581 25087 35615
rect 25087 35581 25096 35615
rect 25044 35572 25096 35581
rect 25320 35615 25372 35624
rect 25320 35581 25329 35615
rect 25329 35581 25363 35615
rect 25363 35581 25372 35615
rect 25320 35572 25372 35581
rect 27804 35572 27856 35624
rect 22100 35436 22152 35488
rect 25136 35436 25188 35488
rect 26792 35479 26844 35488
rect 26792 35445 26801 35479
rect 26801 35445 26835 35479
rect 26835 35445 26844 35479
rect 26792 35436 26844 35445
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 21916 35275 21968 35284
rect 21916 35241 21925 35275
rect 21925 35241 21959 35275
rect 21959 35241 21968 35275
rect 21916 35232 21968 35241
rect 22284 35232 22336 35284
rect 23664 35232 23716 35284
rect 25320 35232 25372 35284
rect 28816 35232 28868 35284
rect 29552 35232 29604 35284
rect 31668 35275 31720 35284
rect 31668 35241 31677 35275
rect 31677 35241 31711 35275
rect 31711 35241 31720 35275
rect 31668 35232 31720 35241
rect 18604 35071 18656 35080
rect 18604 35037 18613 35071
rect 18613 35037 18647 35071
rect 18647 35037 18656 35071
rect 18604 35028 18656 35037
rect 23020 35096 23072 35148
rect 22284 35071 22336 35080
rect 22284 35037 22293 35071
rect 22293 35037 22327 35071
rect 22327 35037 22336 35071
rect 22284 35028 22336 35037
rect 22468 35028 22520 35080
rect 22652 35028 22704 35080
rect 24860 35028 24912 35080
rect 25688 35071 25740 35080
rect 25688 35037 25697 35071
rect 25697 35037 25731 35071
rect 25731 35037 25740 35071
rect 25688 35028 25740 35037
rect 27804 35096 27856 35148
rect 28816 35139 28868 35148
rect 28816 35105 28825 35139
rect 28825 35105 28859 35139
rect 28859 35105 28868 35139
rect 28816 35096 28868 35105
rect 25872 35028 25924 35080
rect 26056 35071 26108 35080
rect 26056 35037 26065 35071
rect 26065 35037 26099 35071
rect 26099 35037 26108 35071
rect 26056 35028 26108 35037
rect 26332 35028 26384 35080
rect 26424 34960 26476 35012
rect 26792 34960 26844 35012
rect 30380 35028 30432 35080
rect 30656 35028 30708 35080
rect 31852 35071 31904 35080
rect 31852 35037 31861 35071
rect 31861 35037 31895 35071
rect 31895 35037 31904 35071
rect 31852 35028 31904 35037
rect 29276 35003 29328 35012
rect 29276 34969 29285 35003
rect 29285 34969 29319 35003
rect 29319 34969 29328 35003
rect 29276 34960 29328 34969
rect 16856 34892 16908 34944
rect 26608 34892 26660 34944
rect 27068 34935 27120 34944
rect 27068 34901 27077 34935
rect 27077 34901 27111 34935
rect 27111 34901 27120 34935
rect 27068 34892 27120 34901
rect 29184 34892 29236 34944
rect 31208 34935 31260 34944
rect 31208 34901 31217 34935
rect 31217 34901 31251 34935
rect 31251 34901 31260 34935
rect 31208 34892 31260 34901
rect 4874 34790 4926 34842
rect 4938 34790 4990 34842
rect 5002 34790 5054 34842
rect 5066 34790 5118 34842
rect 5130 34790 5182 34842
rect 35594 34790 35646 34842
rect 35658 34790 35710 34842
rect 35722 34790 35774 34842
rect 35786 34790 35838 34842
rect 35850 34790 35902 34842
rect 24860 34731 24912 34740
rect 24860 34697 24869 34731
rect 24869 34697 24903 34731
rect 24903 34697 24912 34731
rect 24860 34688 24912 34697
rect 25044 34688 25096 34740
rect 27804 34688 27856 34740
rect 18052 34620 18104 34672
rect 16856 34595 16908 34604
rect 16856 34561 16865 34595
rect 16865 34561 16899 34595
rect 16899 34561 16908 34595
rect 16856 34552 16908 34561
rect 21272 34595 21324 34604
rect 21272 34561 21281 34595
rect 21281 34561 21315 34595
rect 21315 34561 21324 34595
rect 21272 34552 21324 34561
rect 22652 34595 22704 34604
rect 22652 34561 22661 34595
rect 22661 34561 22695 34595
rect 22695 34561 22704 34595
rect 22652 34552 22704 34561
rect 25688 34620 25740 34672
rect 27068 34620 27120 34672
rect 30380 34620 30432 34672
rect 16948 34527 17000 34536
rect 16948 34493 16957 34527
rect 16957 34493 16991 34527
rect 16991 34493 17000 34527
rect 16948 34484 17000 34493
rect 17224 34484 17276 34536
rect 18144 34484 18196 34536
rect 18604 34484 18656 34536
rect 22100 34484 22152 34536
rect 23112 34527 23164 34536
rect 23112 34493 23121 34527
rect 23121 34493 23155 34527
rect 23155 34493 23164 34527
rect 23112 34484 23164 34493
rect 23388 34527 23440 34536
rect 23388 34493 23397 34527
rect 23397 34493 23431 34527
rect 23431 34493 23440 34527
rect 23388 34484 23440 34493
rect 26424 34595 26476 34604
rect 26424 34561 26433 34595
rect 26433 34561 26467 34595
rect 26467 34561 26476 34595
rect 26424 34552 26476 34561
rect 26056 34484 26108 34536
rect 26792 34595 26844 34604
rect 26792 34561 26801 34595
rect 26801 34561 26835 34595
rect 26835 34561 26844 34595
rect 26792 34552 26844 34561
rect 28816 34552 28868 34604
rect 26608 34484 26660 34536
rect 30472 34527 30524 34536
rect 30472 34493 30481 34527
rect 30481 34493 30515 34527
rect 30515 34493 30524 34527
rect 30472 34484 30524 34493
rect 32312 34484 32364 34536
rect 33232 34527 33284 34536
rect 33232 34493 33241 34527
rect 33241 34493 33275 34527
rect 33275 34493 33284 34527
rect 33232 34484 33284 34493
rect 34428 34484 34480 34536
rect 21180 34391 21232 34400
rect 21180 34357 21189 34391
rect 21189 34357 21223 34391
rect 21223 34357 21232 34391
rect 21180 34348 21232 34357
rect 24952 34391 25004 34400
rect 24952 34357 24961 34391
rect 24961 34357 24995 34391
rect 24995 34357 25004 34391
rect 24952 34348 25004 34357
rect 26700 34348 26752 34400
rect 26792 34348 26844 34400
rect 27252 34348 27304 34400
rect 32128 34348 32180 34400
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 17132 33940 17184 33992
rect 18144 34144 18196 34196
rect 21272 34187 21324 34196
rect 21272 34153 21281 34187
rect 21281 34153 21315 34187
rect 21315 34153 21324 34187
rect 21272 34144 21324 34153
rect 20260 34119 20312 34128
rect 20260 34085 20269 34119
rect 20269 34085 20303 34119
rect 20303 34085 20312 34119
rect 20260 34076 20312 34085
rect 18052 34008 18104 34060
rect 19800 34008 19852 34060
rect 21640 34076 21692 34128
rect 25780 34144 25832 34196
rect 26240 34076 26292 34128
rect 30472 34144 30524 34196
rect 30656 34076 30708 34128
rect 17868 33983 17920 33992
rect 17868 33949 17877 33983
rect 17877 33949 17911 33983
rect 17911 33949 17920 33983
rect 17868 33940 17920 33949
rect 16948 33804 17000 33856
rect 17776 33804 17828 33856
rect 22008 33940 22060 33992
rect 23112 33940 23164 33992
rect 30288 34008 30340 34060
rect 31852 34144 31904 34196
rect 32680 34144 32732 34196
rect 31116 34076 31168 34128
rect 33232 34144 33284 34196
rect 33784 34076 33836 34128
rect 31208 34008 31260 34060
rect 32036 34008 32088 34060
rect 18328 33804 18380 33856
rect 21180 33872 21232 33924
rect 22560 33872 22612 33924
rect 25780 33983 25832 33992
rect 25780 33949 25789 33983
rect 25789 33949 25823 33983
rect 25823 33949 25832 33983
rect 25780 33940 25832 33949
rect 26332 33983 26384 33992
rect 26332 33949 26341 33983
rect 26341 33949 26375 33983
rect 26375 33949 26384 33983
rect 26332 33940 26384 33949
rect 26516 33940 26568 33992
rect 27160 33940 27212 33992
rect 30656 33940 30708 33992
rect 31116 33983 31168 33992
rect 31116 33949 31125 33983
rect 31125 33949 31159 33983
rect 31159 33949 31168 33983
rect 31116 33940 31168 33949
rect 32128 33983 32180 33992
rect 32128 33949 32137 33983
rect 32137 33949 32171 33983
rect 32171 33949 32180 33983
rect 32128 33940 32180 33949
rect 33048 34008 33100 34060
rect 25044 33872 25096 33924
rect 31668 33872 31720 33924
rect 22192 33804 22244 33856
rect 25872 33847 25924 33856
rect 25872 33813 25881 33847
rect 25881 33813 25915 33847
rect 25915 33813 25924 33847
rect 25872 33804 25924 33813
rect 26332 33804 26384 33856
rect 27344 33804 27396 33856
rect 32680 33983 32732 33992
rect 32680 33949 32689 33983
rect 32689 33949 32723 33983
rect 32723 33949 32732 33983
rect 32680 33940 32732 33949
rect 32772 33983 32824 33992
rect 32772 33949 32781 33983
rect 32781 33949 32815 33983
rect 32815 33949 32824 33983
rect 32772 33940 32824 33949
rect 33140 33872 33192 33924
rect 33416 33983 33468 33992
rect 33416 33949 33425 33983
rect 33425 33949 33459 33983
rect 33459 33949 33468 33983
rect 33416 33940 33468 33949
rect 32772 33804 32824 33856
rect 34428 34051 34480 34060
rect 33784 33915 33836 33924
rect 33784 33881 33793 33915
rect 33793 33881 33827 33915
rect 33827 33881 33836 33915
rect 34428 34017 34437 34051
rect 34437 34017 34471 34051
rect 34471 34017 34480 34051
rect 34428 34008 34480 34017
rect 33784 33872 33836 33881
rect 37096 33847 37148 33856
rect 37096 33813 37105 33847
rect 37105 33813 37139 33847
rect 37139 33813 37148 33847
rect 37096 33804 37148 33813
rect 4874 33702 4926 33754
rect 4938 33702 4990 33754
rect 5002 33702 5054 33754
rect 5066 33702 5118 33754
rect 5130 33702 5182 33754
rect 35594 33702 35646 33754
rect 35658 33702 35710 33754
rect 35722 33702 35774 33754
rect 35786 33702 35838 33754
rect 35850 33702 35902 33754
rect 15936 33532 15988 33584
rect 17960 33532 18012 33584
rect 20260 33532 20312 33584
rect 21640 33643 21692 33652
rect 21640 33609 21649 33643
rect 21649 33609 21683 33643
rect 21683 33609 21692 33643
rect 21640 33600 21692 33609
rect 23388 33600 23440 33652
rect 26608 33600 26660 33652
rect 27252 33600 27304 33652
rect 32036 33600 32088 33652
rect 33416 33600 33468 33652
rect 22284 33532 22336 33584
rect 16948 33507 17000 33516
rect 16948 33473 16957 33507
rect 16957 33473 16991 33507
rect 16991 33473 17000 33507
rect 16948 33464 17000 33473
rect 17132 33507 17184 33516
rect 17132 33473 17141 33507
rect 17141 33473 17175 33507
rect 17175 33473 17184 33507
rect 17132 33464 17184 33473
rect 22008 33507 22060 33516
rect 22008 33473 22017 33507
rect 22017 33473 22051 33507
rect 22051 33473 22060 33507
rect 22008 33464 22060 33473
rect 22192 33507 22244 33516
rect 22192 33473 22201 33507
rect 22201 33473 22235 33507
rect 22235 33473 22244 33507
rect 24952 33532 25004 33584
rect 26700 33532 26752 33584
rect 27344 33575 27396 33584
rect 27344 33541 27353 33575
rect 27353 33541 27387 33575
rect 27387 33541 27396 33575
rect 27344 33532 27396 33541
rect 30380 33532 30432 33584
rect 22192 33464 22244 33473
rect 17224 33439 17276 33448
rect 17224 33405 17233 33439
rect 17233 33405 17267 33439
rect 17267 33405 17276 33439
rect 17224 33396 17276 33405
rect 18236 33396 18288 33448
rect 20628 33396 20680 33448
rect 22560 33396 22612 33448
rect 17040 33303 17092 33312
rect 17040 33269 17049 33303
rect 17049 33269 17083 33303
rect 17083 33269 17092 33303
rect 17040 33260 17092 33269
rect 18052 33260 18104 33312
rect 18972 33303 19024 33312
rect 18972 33269 18981 33303
rect 18981 33269 19015 33303
rect 19015 33269 19024 33303
rect 18972 33260 19024 33269
rect 21824 33303 21876 33312
rect 21824 33269 21833 33303
rect 21833 33269 21867 33303
rect 21867 33269 21876 33303
rect 21824 33260 21876 33269
rect 23572 33303 23624 33312
rect 23572 33269 23581 33303
rect 23581 33269 23615 33303
rect 23615 33269 23624 33303
rect 23572 33260 23624 33269
rect 24860 33464 24912 33516
rect 25044 33507 25096 33516
rect 25044 33473 25053 33507
rect 25053 33473 25087 33507
rect 25087 33473 25096 33507
rect 25044 33464 25096 33473
rect 27804 33464 27856 33516
rect 31116 33507 31168 33516
rect 31116 33473 31125 33507
rect 31125 33473 31159 33507
rect 31159 33473 31168 33507
rect 31116 33464 31168 33473
rect 25320 33439 25372 33448
rect 25320 33405 25329 33439
rect 25329 33405 25363 33439
rect 25363 33405 25372 33439
rect 25320 33396 25372 33405
rect 30656 33328 30708 33380
rect 25964 33260 26016 33312
rect 27160 33303 27212 33312
rect 27160 33269 27169 33303
rect 27169 33269 27203 33303
rect 27203 33269 27212 33303
rect 27160 33260 27212 33269
rect 30564 33260 30616 33312
rect 31668 33396 31720 33448
rect 32956 33464 33008 33516
rect 33692 33396 33744 33448
rect 33048 33303 33100 33312
rect 33048 33269 33057 33303
rect 33057 33269 33091 33303
rect 33091 33269 33100 33303
rect 33048 33260 33100 33269
rect 33416 33303 33468 33312
rect 33416 33269 33425 33303
rect 33425 33269 33459 33303
rect 33459 33269 33468 33303
rect 33416 33260 33468 33269
rect 33784 33303 33836 33312
rect 33784 33269 33793 33303
rect 33793 33269 33827 33303
rect 33827 33269 33836 33303
rect 33784 33260 33836 33269
rect 34060 33303 34112 33312
rect 34060 33269 34069 33303
rect 34069 33269 34103 33303
rect 34103 33269 34112 33303
rect 34060 33260 34112 33269
rect 37464 33532 37516 33584
rect 38660 33464 38712 33516
rect 37280 33439 37332 33448
rect 37280 33405 37289 33439
rect 37289 33405 37323 33439
rect 37323 33405 37332 33439
rect 37280 33396 37332 33405
rect 36636 33328 36688 33380
rect 37372 33260 37424 33312
rect 39028 33303 39080 33312
rect 39028 33269 39037 33303
rect 39037 33269 39071 33303
rect 39071 33269 39080 33303
rect 39028 33260 39080 33269
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 18236 33099 18288 33108
rect 18236 33065 18245 33099
rect 18245 33065 18279 33099
rect 18279 33065 18288 33099
rect 18236 33056 18288 33065
rect 19800 33099 19852 33108
rect 19800 33065 19809 33099
rect 19809 33065 19843 33099
rect 19843 33065 19852 33099
rect 19800 33056 19852 33065
rect 22560 33099 22612 33108
rect 22560 33065 22569 33099
rect 22569 33065 22603 33099
rect 22603 33065 22612 33099
rect 22560 33056 22612 33065
rect 18328 33031 18380 33040
rect 18328 32997 18337 33031
rect 18337 32997 18371 33031
rect 18371 32997 18380 33031
rect 18328 32988 18380 32997
rect 13912 32852 13964 32904
rect 18972 32920 19024 32972
rect 21824 32920 21876 32972
rect 17868 32852 17920 32904
rect 18052 32852 18104 32904
rect 18144 32895 18196 32904
rect 18144 32861 18153 32895
rect 18153 32861 18187 32895
rect 18187 32861 18196 32895
rect 18144 32852 18196 32861
rect 20628 32852 20680 32904
rect 22284 32920 22336 32972
rect 23756 33056 23808 33108
rect 23572 32988 23624 33040
rect 25228 33056 25280 33108
rect 25320 33056 25372 33108
rect 26332 33056 26384 33108
rect 31116 33056 31168 33108
rect 33140 33056 33192 33108
rect 33968 33056 34020 33108
rect 37464 33056 37516 33108
rect 25688 32988 25740 33040
rect 32772 32988 32824 33040
rect 37188 32988 37240 33040
rect 23572 32852 23624 32904
rect 23848 32852 23900 32904
rect 24860 32852 24912 32904
rect 26240 32920 26292 32972
rect 27804 32963 27856 32972
rect 27804 32929 27813 32963
rect 27813 32929 27847 32963
rect 27847 32929 27856 32963
rect 27804 32920 27856 32929
rect 14648 32827 14700 32836
rect 14648 32793 14657 32827
rect 14657 32793 14691 32827
rect 14691 32793 14700 32827
rect 14648 32784 14700 32793
rect 15936 32784 15988 32836
rect 17776 32827 17828 32836
rect 17776 32793 17785 32827
rect 17785 32793 17819 32827
rect 17819 32793 17828 32827
rect 17776 32784 17828 32793
rect 16304 32716 16356 32768
rect 16488 32716 16540 32768
rect 18236 32784 18288 32836
rect 19248 32759 19300 32768
rect 19248 32725 19257 32759
rect 19257 32725 19291 32759
rect 19291 32725 19300 32759
rect 19248 32716 19300 32725
rect 22008 32716 22060 32768
rect 24584 32759 24636 32768
rect 24584 32725 24593 32759
rect 24593 32725 24627 32759
rect 24627 32725 24636 32759
rect 24584 32716 24636 32725
rect 25964 32895 26016 32904
rect 25964 32861 25973 32895
rect 25973 32861 26007 32895
rect 26007 32861 26016 32895
rect 25964 32852 26016 32861
rect 30564 32895 30616 32904
rect 30564 32861 30573 32895
rect 30573 32861 30607 32895
rect 30607 32861 30616 32895
rect 30564 32852 30616 32861
rect 30656 32895 30708 32904
rect 30656 32861 30665 32895
rect 30665 32861 30699 32895
rect 30699 32861 30708 32895
rect 30656 32852 30708 32861
rect 26792 32784 26844 32836
rect 27528 32827 27580 32836
rect 27528 32793 27537 32827
rect 27537 32793 27571 32827
rect 27571 32793 27580 32827
rect 27528 32784 27580 32793
rect 28908 32784 28960 32836
rect 32772 32852 32824 32904
rect 32588 32784 32640 32836
rect 25872 32716 25924 32768
rect 27160 32716 27212 32768
rect 30840 32759 30892 32768
rect 30840 32725 30849 32759
rect 30849 32725 30883 32759
rect 30883 32725 30892 32759
rect 30840 32716 30892 32725
rect 33508 32895 33560 32904
rect 33508 32861 33517 32895
rect 33517 32861 33551 32895
rect 33551 32861 33560 32895
rect 33508 32852 33560 32861
rect 33600 32852 33652 32904
rect 33784 32895 33836 32904
rect 33784 32861 33793 32895
rect 33793 32861 33827 32895
rect 33827 32861 33836 32895
rect 33784 32852 33836 32861
rect 34244 32852 34296 32904
rect 36820 32920 36872 32972
rect 34520 32895 34572 32904
rect 34520 32861 34529 32895
rect 34529 32861 34563 32895
rect 34563 32861 34572 32895
rect 34520 32852 34572 32861
rect 37096 32852 37148 32904
rect 35992 32784 36044 32836
rect 36084 32827 36136 32836
rect 36084 32793 36093 32827
rect 36093 32793 36127 32827
rect 36127 32793 36136 32827
rect 36084 32784 36136 32793
rect 33692 32716 33744 32768
rect 36268 32716 36320 32768
rect 36728 32716 36780 32768
rect 37556 32759 37608 32768
rect 37556 32725 37565 32759
rect 37565 32725 37599 32759
rect 37599 32725 37608 32759
rect 37556 32716 37608 32725
rect 37832 32827 37884 32836
rect 37832 32793 37841 32827
rect 37841 32793 37875 32827
rect 37875 32793 37884 32827
rect 37832 32784 37884 32793
rect 39028 32784 39080 32836
rect 38568 32716 38620 32768
rect 4874 32614 4926 32666
rect 4938 32614 4990 32666
rect 5002 32614 5054 32666
rect 5066 32614 5118 32666
rect 5130 32614 5182 32666
rect 35594 32614 35646 32666
rect 35658 32614 35710 32666
rect 35722 32614 35774 32666
rect 35786 32614 35838 32666
rect 35850 32614 35902 32666
rect 14648 32512 14700 32564
rect 26792 32512 26844 32564
rect 27252 32512 27304 32564
rect 27528 32512 27580 32564
rect 30472 32512 30524 32564
rect 13912 32444 13964 32496
rect 16304 32419 16356 32428
rect 16304 32385 16313 32419
rect 16313 32385 16347 32419
rect 16347 32385 16356 32419
rect 16304 32376 16356 32385
rect 17316 32376 17368 32428
rect 26332 32376 26384 32428
rect 17040 32308 17092 32360
rect 26516 32351 26568 32360
rect 26516 32317 26525 32351
rect 26525 32317 26559 32351
rect 26559 32317 26568 32351
rect 26516 32308 26568 32317
rect 27160 32419 27212 32428
rect 27160 32385 27169 32419
rect 27169 32385 27203 32419
rect 27203 32385 27212 32419
rect 27160 32376 27212 32385
rect 30840 32444 30892 32496
rect 30472 32419 30524 32428
rect 30472 32385 30481 32419
rect 30481 32385 30515 32419
rect 30515 32385 30524 32419
rect 30472 32376 30524 32385
rect 30564 32376 30616 32428
rect 31300 32308 31352 32360
rect 32956 32444 33008 32496
rect 34244 32512 34296 32564
rect 32864 32376 32916 32428
rect 33784 32444 33836 32496
rect 34152 32444 34204 32496
rect 35992 32512 36044 32564
rect 36084 32555 36136 32564
rect 36084 32521 36093 32555
rect 36093 32521 36127 32555
rect 36127 32521 36136 32555
rect 36084 32512 36136 32521
rect 36636 32555 36688 32564
rect 34336 32376 34388 32428
rect 34428 32376 34480 32428
rect 35440 32444 35492 32496
rect 34520 32308 34572 32360
rect 34888 32376 34940 32428
rect 36268 32419 36320 32428
rect 36268 32385 36277 32419
rect 36277 32385 36311 32419
rect 36311 32385 36320 32419
rect 36268 32376 36320 32385
rect 36636 32521 36645 32555
rect 36645 32521 36679 32555
rect 36679 32521 36688 32555
rect 36636 32512 36688 32521
rect 37556 32444 37608 32496
rect 29368 32240 29420 32292
rect 33048 32240 33100 32292
rect 17960 32215 18012 32224
rect 17960 32181 17969 32215
rect 17969 32181 18003 32215
rect 18003 32181 18012 32215
rect 17960 32172 18012 32181
rect 18328 32172 18380 32224
rect 29920 32215 29972 32224
rect 29920 32181 29929 32215
rect 29929 32181 29963 32215
rect 29963 32181 29972 32215
rect 29920 32172 29972 32181
rect 30104 32172 30156 32224
rect 33324 32215 33376 32224
rect 33324 32181 33333 32215
rect 33333 32181 33367 32215
rect 33367 32181 33376 32215
rect 33324 32172 33376 32181
rect 33600 32172 33652 32224
rect 33876 32215 33928 32224
rect 33876 32181 33885 32215
rect 33885 32181 33919 32215
rect 33919 32181 33928 32215
rect 33876 32172 33928 32181
rect 34244 32172 34296 32224
rect 35992 32240 36044 32292
rect 36728 32240 36780 32292
rect 35440 32172 35492 32224
rect 37832 32376 37884 32428
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 16488 31968 16540 32020
rect 18144 31968 18196 32020
rect 19432 32011 19484 32020
rect 19432 31977 19441 32011
rect 19441 31977 19475 32011
rect 19475 31977 19484 32011
rect 19432 31968 19484 31977
rect 22100 31968 22152 32020
rect 24584 31968 24636 32020
rect 28908 31968 28960 32020
rect 29920 31968 29972 32020
rect 31300 32011 31352 32020
rect 31300 31977 31309 32011
rect 31309 31977 31343 32011
rect 31343 31977 31352 32011
rect 31300 31968 31352 31977
rect 33784 32011 33836 32020
rect 33784 31977 33793 32011
rect 33793 31977 33827 32011
rect 33827 31977 33836 32011
rect 33784 31968 33836 31977
rect 18604 31832 18656 31884
rect 20628 31832 20680 31884
rect 15568 31807 15620 31816
rect 15568 31773 15577 31807
rect 15577 31773 15611 31807
rect 15611 31773 15620 31807
rect 15568 31764 15620 31773
rect 15844 31764 15896 31816
rect 17960 31764 18012 31816
rect 18420 31764 18472 31816
rect 19248 31807 19300 31816
rect 19248 31773 19257 31807
rect 19257 31773 19291 31807
rect 19291 31773 19300 31807
rect 19248 31764 19300 31773
rect 23664 31832 23716 31884
rect 25596 31832 25648 31884
rect 17316 31696 17368 31748
rect 25412 31807 25464 31816
rect 25412 31773 25421 31807
rect 25421 31773 25455 31807
rect 25455 31773 25464 31807
rect 25412 31764 25464 31773
rect 26240 31807 26292 31816
rect 26240 31773 26249 31807
rect 26249 31773 26283 31807
rect 26283 31773 26292 31807
rect 26240 31764 26292 31773
rect 29000 31832 29052 31884
rect 16120 31628 16172 31680
rect 18236 31671 18288 31680
rect 18236 31637 18245 31671
rect 18245 31637 18279 31671
rect 18279 31637 18288 31671
rect 18236 31628 18288 31637
rect 19708 31671 19760 31680
rect 19708 31637 19717 31671
rect 19717 31637 19751 31671
rect 19751 31637 19760 31671
rect 19708 31628 19760 31637
rect 20536 31739 20588 31748
rect 20536 31705 20545 31739
rect 20545 31705 20579 31739
rect 20579 31705 20588 31739
rect 20536 31696 20588 31705
rect 22284 31696 22336 31748
rect 22376 31739 22428 31748
rect 22376 31705 22385 31739
rect 22385 31705 22419 31739
rect 22419 31705 22428 31739
rect 22376 31696 22428 31705
rect 23756 31696 23808 31748
rect 29368 31807 29420 31816
rect 29368 31773 29377 31807
rect 29377 31773 29411 31807
rect 29411 31773 29420 31807
rect 29368 31764 29420 31773
rect 33508 31900 33560 31952
rect 33600 31900 33652 31952
rect 37372 31968 37424 32020
rect 37556 31968 37608 32020
rect 34244 31900 34296 31952
rect 36728 31900 36780 31952
rect 38752 31900 38804 31952
rect 34796 31832 34848 31884
rect 38384 31832 38436 31884
rect 32312 31807 32364 31816
rect 32312 31773 32321 31807
rect 32321 31773 32355 31807
rect 32355 31773 32364 31807
rect 32312 31764 32364 31773
rect 32956 31764 33008 31816
rect 33232 31807 33284 31816
rect 33232 31773 33241 31807
rect 33241 31773 33275 31807
rect 33275 31773 33284 31807
rect 33232 31764 33284 31773
rect 33416 31764 33468 31816
rect 33876 31764 33928 31816
rect 33968 31764 34020 31816
rect 34704 31764 34756 31816
rect 37832 31764 37884 31816
rect 30104 31696 30156 31748
rect 31576 31696 31628 31748
rect 21456 31628 21508 31680
rect 22560 31628 22612 31680
rect 24400 31671 24452 31680
rect 24400 31637 24409 31671
rect 24409 31637 24443 31671
rect 24443 31637 24452 31671
rect 24400 31628 24452 31637
rect 29368 31671 29420 31680
rect 29368 31637 29377 31671
rect 29377 31637 29411 31671
rect 29411 31637 29420 31671
rect 29368 31628 29420 31637
rect 30564 31628 30616 31680
rect 32864 31628 32916 31680
rect 33324 31739 33376 31748
rect 33324 31705 33333 31739
rect 33333 31705 33367 31739
rect 33367 31705 33376 31739
rect 33324 31696 33376 31705
rect 33508 31671 33560 31680
rect 33508 31637 33517 31671
rect 33517 31637 33551 31671
rect 33551 31637 33560 31671
rect 33508 31628 33560 31637
rect 33692 31628 33744 31680
rect 34612 31696 34664 31748
rect 37924 31739 37976 31748
rect 37924 31705 37933 31739
rect 37933 31705 37967 31739
rect 37967 31705 37976 31739
rect 37924 31696 37976 31705
rect 34520 31628 34572 31680
rect 4874 31526 4926 31578
rect 4938 31526 4990 31578
rect 5002 31526 5054 31578
rect 5066 31526 5118 31578
rect 5130 31526 5182 31578
rect 35594 31526 35646 31578
rect 35658 31526 35710 31578
rect 35722 31526 35774 31578
rect 35786 31526 35838 31578
rect 35850 31526 35902 31578
rect 15568 31424 15620 31476
rect 18144 31467 18196 31476
rect 18144 31433 18169 31467
rect 18169 31433 18196 31467
rect 18144 31424 18196 31433
rect 18420 31424 18472 31476
rect 22376 31424 22428 31476
rect 23848 31467 23900 31476
rect 23848 31433 23857 31467
rect 23857 31433 23891 31467
rect 23891 31433 23900 31467
rect 23848 31424 23900 31433
rect 15936 31356 15988 31408
rect 17868 31356 17920 31408
rect 22284 31399 22336 31408
rect 13912 31331 13964 31340
rect 13912 31297 13921 31331
rect 13921 31297 13955 31331
rect 13955 31297 13964 31331
rect 13912 31288 13964 31297
rect 16120 31331 16172 31340
rect 16120 31297 16129 31331
rect 16129 31297 16163 31331
rect 16163 31297 16172 31331
rect 16120 31288 16172 31297
rect 16488 31220 16540 31272
rect 17224 31263 17276 31272
rect 17224 31229 17233 31263
rect 17233 31229 17267 31263
rect 17267 31229 17276 31263
rect 22284 31365 22311 31399
rect 22311 31365 22336 31399
rect 22284 31356 22336 31365
rect 22560 31356 22612 31408
rect 17224 31220 17276 31229
rect 15844 31152 15896 31204
rect 15936 31084 15988 31136
rect 16488 31084 16540 31136
rect 17776 31084 17828 31136
rect 18512 31127 18564 31136
rect 18512 31093 18521 31127
rect 18521 31093 18555 31127
rect 18555 31093 18564 31127
rect 18512 31084 18564 31093
rect 21456 31331 21508 31340
rect 21456 31297 21465 31331
rect 21465 31297 21499 31331
rect 21499 31297 21508 31331
rect 21456 31288 21508 31297
rect 19432 31220 19484 31272
rect 19800 31263 19852 31272
rect 19800 31229 19809 31263
rect 19809 31229 19843 31263
rect 19843 31229 19852 31263
rect 19800 31220 19852 31229
rect 20536 31263 20588 31272
rect 20536 31229 20545 31263
rect 20545 31229 20579 31263
rect 20579 31229 20588 31263
rect 20536 31220 20588 31229
rect 22008 31331 22060 31340
rect 22008 31297 22017 31331
rect 22017 31297 22051 31331
rect 22051 31297 22060 31331
rect 22008 31288 22060 31297
rect 23388 31399 23440 31408
rect 23388 31365 23397 31399
rect 23397 31365 23431 31399
rect 23431 31365 23440 31399
rect 23388 31356 23440 31365
rect 24860 31424 24912 31476
rect 27436 31424 27488 31476
rect 24676 31331 24728 31340
rect 24676 31297 24685 31331
rect 24685 31297 24719 31331
rect 24719 31297 24728 31331
rect 24676 31288 24728 31297
rect 25688 31331 25740 31340
rect 25688 31297 25697 31331
rect 25697 31297 25731 31331
rect 25731 31297 25740 31331
rect 29000 31356 29052 31408
rect 29552 31424 29604 31476
rect 30196 31424 30248 31476
rect 36728 31467 36780 31476
rect 36728 31433 36737 31467
rect 36737 31433 36771 31467
rect 36771 31433 36780 31467
rect 36728 31424 36780 31433
rect 32036 31356 32088 31408
rect 32312 31356 32364 31408
rect 36636 31356 36688 31408
rect 37924 31424 37976 31476
rect 25688 31288 25740 31297
rect 21640 31152 21692 31204
rect 19432 31084 19484 31136
rect 21824 31152 21876 31204
rect 22192 31152 22244 31204
rect 21916 31084 21968 31136
rect 25412 31152 25464 31204
rect 26332 31263 26384 31272
rect 26332 31229 26341 31263
rect 26341 31229 26375 31263
rect 26375 31229 26384 31263
rect 30380 31288 30432 31340
rect 31576 31288 31628 31340
rect 33232 31288 33284 31340
rect 33600 31288 33652 31340
rect 33968 31288 34020 31340
rect 34336 31331 34388 31340
rect 34336 31297 34345 31331
rect 34345 31297 34379 31331
rect 34379 31297 34388 31331
rect 34336 31288 34388 31297
rect 34704 31331 34756 31340
rect 34704 31297 34713 31331
rect 34713 31297 34747 31331
rect 34747 31297 34756 31331
rect 38660 31356 38712 31408
rect 38752 31399 38804 31408
rect 38752 31365 38761 31399
rect 38761 31365 38795 31399
rect 38795 31365 38804 31399
rect 38752 31356 38804 31365
rect 34704 31288 34756 31297
rect 26332 31220 26384 31229
rect 29368 31220 29420 31272
rect 34428 31220 34480 31272
rect 36360 31220 36412 31272
rect 38660 31220 38712 31272
rect 22928 31084 22980 31136
rect 23664 31127 23716 31136
rect 23664 31093 23673 31127
rect 23673 31093 23707 31127
rect 23707 31093 23716 31127
rect 23664 31084 23716 31093
rect 25504 31084 25556 31136
rect 30564 31084 30616 31136
rect 32956 31084 33008 31136
rect 34060 31127 34112 31136
rect 34060 31093 34069 31127
rect 34069 31093 34103 31127
rect 34103 31093 34112 31127
rect 34060 31084 34112 31093
rect 34612 31127 34664 31136
rect 34612 31093 34621 31127
rect 34621 31093 34655 31127
rect 34655 31093 34664 31127
rect 34612 31084 34664 31093
rect 34704 31084 34756 31136
rect 36820 31084 36872 31136
rect 38752 31084 38804 31136
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 17224 30880 17276 30932
rect 18604 30880 18656 30932
rect 22008 30880 22060 30932
rect 25044 30923 25096 30932
rect 25044 30889 25053 30923
rect 25053 30889 25087 30923
rect 25087 30889 25096 30923
rect 25044 30880 25096 30889
rect 25688 30880 25740 30932
rect 26332 30880 26384 30932
rect 30104 30880 30156 30932
rect 33876 30880 33928 30932
rect 34060 30880 34112 30932
rect 34796 30880 34848 30932
rect 36360 30923 36412 30932
rect 36360 30889 36369 30923
rect 36369 30889 36403 30923
rect 36403 30889 36412 30923
rect 36360 30880 36412 30889
rect 37832 30880 37884 30932
rect 17316 30719 17368 30728
rect 17316 30685 17325 30719
rect 17325 30685 17359 30719
rect 17359 30685 17368 30719
rect 17316 30676 17368 30685
rect 17776 30719 17828 30728
rect 17776 30685 17785 30719
rect 17785 30685 17819 30719
rect 17819 30685 17828 30719
rect 17776 30676 17828 30685
rect 18420 30812 18472 30864
rect 21916 30812 21968 30864
rect 22744 30812 22796 30864
rect 25596 30787 25648 30796
rect 25596 30753 25605 30787
rect 25605 30753 25639 30787
rect 25639 30753 25648 30787
rect 25596 30744 25648 30753
rect 29000 30744 29052 30796
rect 32036 30744 32088 30796
rect 18512 30676 18564 30728
rect 19432 30719 19484 30728
rect 19432 30685 19441 30719
rect 19441 30685 19475 30719
rect 19475 30685 19484 30719
rect 19432 30676 19484 30685
rect 22192 30676 22244 30728
rect 22928 30719 22980 30728
rect 22928 30685 22937 30719
rect 22937 30685 22971 30719
rect 22971 30685 22980 30719
rect 22928 30676 22980 30685
rect 24400 30676 24452 30728
rect 25504 30719 25556 30728
rect 25504 30685 25513 30719
rect 25513 30685 25547 30719
rect 25547 30685 25556 30719
rect 25504 30676 25556 30685
rect 30472 30719 30524 30728
rect 30472 30685 30481 30719
rect 30481 30685 30515 30719
rect 30515 30685 30524 30719
rect 30472 30676 30524 30685
rect 30564 30719 30616 30728
rect 30564 30685 30573 30719
rect 30573 30685 30607 30719
rect 30607 30685 30616 30719
rect 30564 30676 30616 30685
rect 32772 30676 32824 30728
rect 33508 30787 33560 30796
rect 33508 30753 33517 30787
rect 33517 30753 33551 30787
rect 33551 30753 33560 30787
rect 33508 30744 33560 30753
rect 34152 30855 34204 30864
rect 34152 30821 34161 30855
rect 34161 30821 34195 30855
rect 34195 30821 34204 30855
rect 34152 30812 34204 30821
rect 34612 30744 34664 30796
rect 34704 30676 34756 30728
rect 16488 30608 16540 30660
rect 18236 30608 18288 30660
rect 24860 30651 24912 30660
rect 24860 30617 24869 30651
rect 24869 30617 24903 30651
rect 24903 30617 24912 30651
rect 24860 30608 24912 30617
rect 27436 30608 27488 30660
rect 17960 30540 18012 30592
rect 18696 30540 18748 30592
rect 22744 30540 22796 30592
rect 24676 30540 24728 30592
rect 31576 30608 31628 30660
rect 32220 30540 32272 30592
rect 33968 30608 34020 30660
rect 35348 30651 35400 30660
rect 35348 30617 35357 30651
rect 35357 30617 35391 30651
rect 35391 30617 35400 30651
rect 35348 30608 35400 30617
rect 33232 30540 33284 30592
rect 33784 30583 33836 30592
rect 33784 30549 33793 30583
rect 33793 30549 33827 30583
rect 33827 30549 33836 30583
rect 33784 30540 33836 30549
rect 33876 30540 33928 30592
rect 36636 30719 36688 30728
rect 36636 30685 36645 30719
rect 36645 30685 36679 30719
rect 36679 30685 36688 30719
rect 36636 30676 36688 30685
rect 36912 30719 36964 30728
rect 36912 30685 36921 30719
rect 36921 30685 36955 30719
rect 36955 30685 36964 30719
rect 36912 30676 36964 30685
rect 37280 30608 37332 30660
rect 38568 30608 38620 30660
rect 38752 30651 38804 30660
rect 38752 30617 38761 30651
rect 38761 30617 38795 30651
rect 38795 30617 38804 30651
rect 38752 30608 38804 30617
rect 36820 30540 36872 30592
rect 38844 30540 38896 30592
rect 4874 30438 4926 30490
rect 4938 30438 4990 30490
rect 5002 30438 5054 30490
rect 5066 30438 5118 30490
rect 5130 30438 5182 30490
rect 35594 30438 35646 30490
rect 35658 30438 35710 30490
rect 35722 30438 35774 30490
rect 35786 30438 35838 30490
rect 35850 30438 35902 30490
rect 19800 30379 19852 30388
rect 19800 30345 19809 30379
rect 19809 30345 19843 30379
rect 19843 30345 19852 30379
rect 19800 30336 19852 30345
rect 24860 30336 24912 30388
rect 25044 30379 25096 30388
rect 25044 30345 25053 30379
rect 25053 30345 25087 30379
rect 25087 30345 25096 30379
rect 25044 30336 25096 30345
rect 18420 30268 18472 30320
rect 17316 30200 17368 30252
rect 18696 30132 18748 30184
rect 22468 30311 22520 30320
rect 22468 30277 22477 30311
rect 22477 30277 22511 30311
rect 22511 30277 22520 30311
rect 27436 30336 27488 30388
rect 32220 30336 32272 30388
rect 33600 30336 33652 30388
rect 35348 30336 35400 30388
rect 22468 30268 22520 30277
rect 26240 30268 26292 30320
rect 32588 30268 32640 30320
rect 33876 30268 33928 30320
rect 22100 30200 22152 30252
rect 36636 30268 36688 30320
rect 38844 30311 38896 30320
rect 38844 30277 38853 30311
rect 38853 30277 38887 30311
rect 38887 30277 38896 30311
rect 38844 30268 38896 30277
rect 43352 30268 43404 30320
rect 22836 30175 22888 30184
rect 22836 30141 22845 30175
rect 22845 30141 22879 30175
rect 22879 30141 22888 30175
rect 22836 30132 22888 30141
rect 28264 30132 28316 30184
rect 34152 30200 34204 30252
rect 38568 30243 38620 30252
rect 38568 30209 38577 30243
rect 38577 30209 38611 30243
rect 38611 30209 38620 30243
rect 38568 30200 38620 30209
rect 42432 30243 42484 30252
rect 42432 30209 42441 30243
rect 42441 30209 42475 30243
rect 42475 30209 42484 30243
rect 42432 30200 42484 30209
rect 42524 30243 42576 30252
rect 42524 30209 42533 30243
rect 42533 30209 42567 30243
rect 42567 30209 42576 30243
rect 42524 30200 42576 30209
rect 42708 30243 42760 30252
rect 42708 30209 42717 30243
rect 42717 30209 42751 30243
rect 42751 30209 42760 30243
rect 42708 30200 42760 30209
rect 33784 30132 33836 30184
rect 36912 30132 36964 30184
rect 38752 30132 38804 30184
rect 25228 29996 25280 30048
rect 29644 29996 29696 30048
rect 36636 30064 36688 30116
rect 38568 30064 38620 30116
rect 44732 30132 44784 30184
rect 33600 29996 33652 30048
rect 33968 30039 34020 30048
rect 33968 30005 33977 30039
rect 33977 30005 34011 30039
rect 34011 30005 34020 30039
rect 33968 29996 34020 30005
rect 34612 30039 34664 30048
rect 34612 30005 34621 30039
rect 34621 30005 34655 30039
rect 34655 30005 34664 30039
rect 34612 29996 34664 30005
rect 36544 29996 36596 30048
rect 37464 29996 37516 30048
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 22836 29792 22888 29844
rect 28816 29835 28868 29844
rect 28816 29801 28825 29835
rect 28825 29801 28859 29835
rect 28859 29801 28868 29835
rect 28816 29792 28868 29801
rect 16856 29724 16908 29776
rect 25228 29724 25280 29776
rect 22744 29656 22796 29708
rect 24860 29656 24912 29708
rect 27160 29520 27212 29572
rect 32128 29792 32180 29844
rect 32956 29792 33008 29844
rect 37280 29835 37332 29844
rect 37280 29801 37289 29835
rect 37289 29801 37323 29835
rect 37323 29801 37332 29835
rect 37280 29792 37332 29801
rect 37556 29792 37608 29844
rect 29092 29724 29144 29776
rect 32496 29724 32548 29776
rect 33232 29724 33284 29776
rect 29276 29631 29328 29640
rect 29276 29597 29285 29631
rect 29285 29597 29319 29631
rect 29319 29597 29328 29631
rect 29276 29588 29328 29597
rect 29644 29656 29696 29708
rect 30012 29588 30064 29640
rect 33784 29631 33836 29640
rect 33784 29597 33793 29631
rect 33793 29597 33827 29631
rect 33827 29597 33836 29631
rect 33784 29588 33836 29597
rect 33968 29631 34020 29640
rect 33968 29597 33977 29631
rect 33977 29597 34011 29631
rect 34011 29597 34020 29631
rect 33968 29588 34020 29597
rect 30472 29520 30524 29572
rect 32496 29520 32548 29572
rect 32864 29520 32916 29572
rect 32956 29520 33008 29572
rect 34152 29520 34204 29572
rect 37832 29767 37884 29776
rect 37832 29733 37841 29767
rect 37841 29733 37875 29767
rect 37875 29733 37884 29767
rect 37832 29724 37884 29733
rect 40316 29724 40368 29776
rect 38200 29699 38252 29708
rect 38200 29665 38209 29699
rect 38209 29665 38243 29699
rect 38243 29665 38252 29699
rect 38200 29656 38252 29665
rect 42524 29792 42576 29844
rect 42708 29792 42760 29844
rect 40776 29724 40828 29776
rect 28632 29495 28684 29504
rect 28632 29461 28641 29495
rect 28641 29461 28675 29495
rect 28675 29461 28684 29495
rect 28632 29452 28684 29461
rect 32772 29495 32824 29504
rect 32772 29461 32781 29495
rect 32781 29461 32815 29495
rect 32815 29461 32824 29495
rect 32772 29452 32824 29461
rect 34980 29452 35032 29504
rect 37464 29563 37516 29572
rect 37464 29529 37473 29563
rect 37473 29529 37507 29563
rect 37507 29529 37516 29563
rect 37464 29520 37516 29529
rect 39672 29588 39724 29640
rect 40592 29631 40644 29640
rect 40592 29597 40601 29631
rect 40601 29597 40635 29631
rect 40635 29597 40644 29631
rect 40592 29588 40644 29597
rect 42524 29588 42576 29640
rect 37648 29452 37700 29504
rect 40500 29495 40552 29504
rect 40500 29461 40509 29495
rect 40509 29461 40543 29495
rect 40543 29461 40552 29495
rect 40500 29452 40552 29461
rect 41420 29520 41472 29572
rect 42800 29520 42852 29572
rect 44180 29656 44232 29708
rect 44364 29588 44416 29640
rect 49700 29588 49752 29640
rect 41144 29452 41196 29504
rect 41236 29452 41288 29504
rect 43352 29452 43404 29504
rect 43996 29563 44048 29572
rect 43996 29529 44005 29563
rect 44005 29529 44039 29563
rect 44039 29529 44048 29563
rect 43996 29520 44048 29529
rect 45376 29563 45428 29572
rect 45376 29529 45385 29563
rect 45385 29529 45419 29563
rect 45419 29529 45428 29563
rect 45376 29520 45428 29529
rect 44180 29452 44232 29504
rect 47124 29563 47176 29572
rect 47124 29529 47133 29563
rect 47133 29529 47167 29563
rect 47167 29529 47176 29563
rect 47124 29520 47176 29529
rect 47400 29452 47452 29504
rect 4874 29350 4926 29402
rect 4938 29350 4990 29402
rect 5002 29350 5054 29402
rect 5066 29350 5118 29402
rect 5130 29350 5182 29402
rect 35594 29350 35646 29402
rect 35658 29350 35710 29402
rect 35722 29350 35774 29402
rect 35786 29350 35838 29402
rect 35850 29350 35902 29402
rect 27160 29248 27212 29300
rect 29092 29180 29144 29232
rect 30472 29291 30524 29300
rect 30472 29257 30481 29291
rect 30481 29257 30515 29291
rect 30515 29257 30524 29291
rect 30472 29248 30524 29257
rect 31576 29180 31628 29232
rect 26516 29087 26568 29096
rect 26516 29053 26525 29087
rect 26525 29053 26559 29087
rect 26559 29053 26568 29087
rect 26516 29044 26568 29053
rect 32496 29180 32548 29232
rect 33968 29291 34020 29300
rect 33968 29257 33977 29291
rect 33977 29257 34011 29291
rect 34011 29257 34020 29291
rect 33968 29248 34020 29257
rect 38016 29248 38068 29300
rect 38660 29248 38712 29300
rect 37648 29223 37700 29232
rect 37648 29189 37657 29223
rect 37657 29189 37691 29223
rect 37691 29189 37700 29223
rect 37648 29180 37700 29189
rect 41144 29248 41196 29300
rect 41052 29180 41104 29232
rect 42892 29248 42944 29300
rect 45376 29248 45428 29300
rect 47124 29248 47176 29300
rect 28264 29044 28316 29096
rect 27436 28976 27488 29028
rect 28080 29019 28132 29028
rect 28080 28985 28089 29019
rect 28089 28985 28123 29019
rect 28123 28985 28132 29019
rect 28080 28976 28132 28985
rect 32036 29112 32088 29164
rect 35992 29112 36044 29164
rect 36912 29112 36964 29164
rect 39948 29112 40000 29164
rect 40224 29155 40276 29164
rect 40224 29121 40237 29155
rect 40237 29121 40276 29155
rect 25964 28908 26016 28960
rect 30656 28908 30708 28960
rect 31852 28951 31904 28960
rect 31852 28917 31861 28951
rect 31861 28917 31895 28951
rect 31895 28917 31904 28951
rect 31852 28908 31904 28917
rect 32404 29087 32456 29096
rect 32404 29053 32413 29087
rect 32413 29053 32447 29087
rect 32447 29053 32456 29087
rect 32404 29044 32456 29053
rect 34980 29044 35032 29096
rect 40224 29112 40276 29121
rect 40316 29112 40368 29164
rect 40776 29155 40828 29164
rect 40776 29121 40785 29155
rect 40785 29121 40819 29155
rect 40819 29121 40828 29155
rect 40776 29112 40828 29121
rect 42984 29223 43036 29232
rect 42984 29189 42993 29223
rect 42993 29189 43027 29223
rect 43027 29189 43036 29223
rect 42984 29180 43036 29189
rect 40408 29044 40460 29096
rect 41420 29155 41472 29164
rect 41420 29121 41429 29155
rect 41429 29121 41463 29155
rect 41463 29121 41472 29155
rect 41420 29112 41472 29121
rect 41328 29044 41380 29096
rect 43904 29180 43956 29232
rect 43720 29112 43772 29164
rect 40500 28976 40552 29028
rect 41144 28976 41196 29028
rect 43536 29087 43588 29096
rect 43536 29053 43545 29087
rect 43545 29053 43579 29087
rect 43579 29053 43588 29087
rect 44180 29155 44232 29164
rect 44180 29121 44189 29155
rect 44189 29121 44223 29155
rect 44223 29121 44232 29155
rect 44180 29112 44232 29121
rect 44732 29112 44784 29164
rect 46112 29155 46164 29164
rect 46112 29121 46121 29155
rect 46121 29121 46155 29155
rect 46155 29121 46164 29155
rect 46112 29112 46164 29121
rect 43536 29044 43588 29053
rect 44364 29044 44416 29096
rect 45928 29087 45980 29096
rect 45928 29053 45937 29087
rect 45937 29053 45971 29087
rect 45971 29053 45980 29087
rect 45928 29044 45980 29053
rect 43812 28976 43864 29028
rect 32864 28908 32916 28960
rect 33140 28908 33192 28960
rect 39672 28951 39724 28960
rect 39672 28917 39681 28951
rect 39681 28917 39715 28951
rect 39715 28917 39724 28951
rect 39672 28908 39724 28917
rect 43444 28908 43496 28960
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 26516 28704 26568 28756
rect 25872 28568 25924 28620
rect 28816 28747 28868 28756
rect 28816 28713 28825 28747
rect 28825 28713 28859 28747
rect 28859 28713 28868 28747
rect 28816 28704 28868 28713
rect 30656 28747 30708 28756
rect 30656 28713 30665 28747
rect 30665 28713 30699 28747
rect 30699 28713 30708 28747
rect 30656 28704 30708 28713
rect 31852 28704 31904 28756
rect 32404 28704 32456 28756
rect 33784 28704 33836 28756
rect 38016 28747 38068 28756
rect 38016 28713 38025 28747
rect 38025 28713 38059 28747
rect 38059 28713 38068 28747
rect 38016 28704 38068 28713
rect 38200 28704 38252 28756
rect 42432 28704 42484 28756
rect 43076 28704 43128 28756
rect 40592 28679 40644 28688
rect 40592 28645 40601 28679
rect 40601 28645 40635 28679
rect 40635 28645 40644 28679
rect 40592 28636 40644 28645
rect 41328 28636 41380 28688
rect 43168 28636 43220 28688
rect 45192 28704 45244 28756
rect 46112 28704 46164 28756
rect 44364 28636 44416 28688
rect 44824 28636 44876 28688
rect 29276 28500 29328 28552
rect 35992 28611 36044 28620
rect 35992 28577 36001 28611
rect 36001 28577 36035 28611
rect 36035 28577 36044 28611
rect 35992 28568 36044 28577
rect 25964 28432 26016 28484
rect 27436 28432 27488 28484
rect 30472 28543 30524 28552
rect 30472 28509 30481 28543
rect 30481 28509 30515 28543
rect 30515 28509 30524 28543
rect 30472 28500 30524 28509
rect 32496 28500 32548 28552
rect 32864 28543 32916 28552
rect 32864 28509 32873 28543
rect 32873 28509 32907 28543
rect 32907 28509 32916 28543
rect 32864 28500 32916 28509
rect 33140 28543 33192 28552
rect 33140 28509 33149 28543
rect 33149 28509 33183 28543
rect 33183 28509 33192 28543
rect 33140 28500 33192 28509
rect 39672 28500 39724 28552
rect 40224 28543 40276 28552
rect 40224 28509 40233 28543
rect 40233 28509 40267 28543
rect 40267 28509 40276 28543
rect 40224 28500 40276 28509
rect 40500 28500 40552 28552
rect 42800 28543 42852 28552
rect 42800 28509 42809 28543
rect 42809 28509 42843 28543
rect 42843 28509 42852 28543
rect 42800 28500 42852 28509
rect 43168 28543 43220 28552
rect 43168 28509 43177 28543
rect 43177 28509 43211 28543
rect 43211 28509 43220 28543
rect 43168 28500 43220 28509
rect 43260 28543 43312 28552
rect 43260 28509 43269 28543
rect 43269 28509 43303 28543
rect 43303 28509 43312 28543
rect 43260 28500 43312 28509
rect 43444 28543 43496 28552
rect 43444 28509 43453 28543
rect 43453 28509 43487 28543
rect 43487 28509 43496 28543
rect 43444 28500 43496 28509
rect 30564 28432 30616 28484
rect 32128 28475 32180 28484
rect 32128 28441 32137 28475
rect 32137 28441 32171 28475
rect 32171 28441 32180 28475
rect 32128 28432 32180 28441
rect 32772 28432 32824 28484
rect 36268 28475 36320 28484
rect 36268 28441 36277 28475
rect 36277 28441 36311 28475
rect 36311 28441 36320 28475
rect 36268 28432 36320 28441
rect 38016 28432 38068 28484
rect 38384 28432 38436 28484
rect 38936 28475 38988 28484
rect 38936 28441 38945 28475
rect 38945 28441 38979 28475
rect 38979 28441 38988 28475
rect 38936 28432 38988 28441
rect 41236 28432 41288 28484
rect 42248 28432 42300 28484
rect 43720 28500 43772 28552
rect 43812 28500 43864 28552
rect 43996 28500 44048 28552
rect 45192 28543 45244 28552
rect 45192 28509 45201 28543
rect 45201 28509 45235 28543
rect 45235 28509 45244 28543
rect 45192 28500 45244 28509
rect 45284 28543 45336 28552
rect 45284 28509 45293 28543
rect 45293 28509 45327 28543
rect 45327 28509 45336 28543
rect 45284 28500 45336 28509
rect 45652 28543 45704 28552
rect 45652 28509 45661 28543
rect 45661 28509 45695 28543
rect 45695 28509 45704 28543
rect 45652 28500 45704 28509
rect 50620 28500 50672 28552
rect 44180 28432 44232 28484
rect 44732 28475 44784 28484
rect 44732 28441 44741 28475
rect 44741 28441 44775 28475
rect 44775 28441 44784 28475
rect 44732 28432 44784 28441
rect 30012 28364 30064 28416
rect 37740 28407 37792 28416
rect 37740 28373 37749 28407
rect 37749 28373 37783 28407
rect 37783 28373 37792 28407
rect 37740 28364 37792 28373
rect 43904 28364 43956 28416
rect 44272 28407 44324 28416
rect 44272 28373 44281 28407
rect 44281 28373 44315 28407
rect 44315 28373 44324 28407
rect 44272 28364 44324 28373
rect 49884 28364 49936 28416
rect 4874 28262 4926 28314
rect 4938 28262 4990 28314
rect 5002 28262 5054 28314
rect 5066 28262 5118 28314
rect 5130 28262 5182 28314
rect 35594 28262 35646 28314
rect 35658 28262 35710 28314
rect 35722 28262 35774 28314
rect 35786 28262 35838 28314
rect 35850 28262 35902 28314
rect 27436 28160 27488 28212
rect 28632 28092 28684 28144
rect 30012 28203 30064 28212
rect 30012 28169 30021 28203
rect 30021 28169 30055 28203
rect 30055 28169 30064 28203
rect 30012 28160 30064 28169
rect 36268 28160 36320 28212
rect 41236 28160 41288 28212
rect 42708 28160 42760 28212
rect 43720 28160 43772 28212
rect 44180 28160 44232 28212
rect 36544 28092 36596 28144
rect 37832 28092 37884 28144
rect 40040 28092 40092 28144
rect 44916 28160 44968 28212
rect 38936 28024 38988 28076
rect 42248 28067 42300 28076
rect 42248 28033 42257 28067
rect 42257 28033 42291 28067
rect 42291 28033 42300 28067
rect 42248 28024 42300 28033
rect 42708 28067 42760 28076
rect 42708 28033 42717 28067
rect 42717 28033 42751 28067
rect 42751 28033 42760 28067
rect 42708 28024 42760 28033
rect 42800 28067 42852 28076
rect 42800 28033 42809 28067
rect 42809 28033 42843 28067
rect 42843 28033 42852 28067
rect 42800 28024 42852 28033
rect 42892 28024 42944 28076
rect 43076 28067 43128 28076
rect 43076 28033 43085 28067
rect 43085 28033 43119 28067
rect 43119 28033 43128 28067
rect 43076 28024 43128 28033
rect 43996 28024 44048 28076
rect 48136 28092 48188 28144
rect 49700 28092 49752 28144
rect 28264 27999 28316 28008
rect 28264 27965 28273 27999
rect 28273 27965 28307 27999
rect 28307 27965 28316 27999
rect 28264 27956 28316 27965
rect 37740 27999 37792 28008
rect 37740 27965 37749 27999
rect 37749 27965 37783 27999
rect 37783 27965 37792 27999
rect 37740 27956 37792 27965
rect 37832 27999 37884 28008
rect 37832 27965 37841 27999
rect 37841 27965 37875 27999
rect 37875 27965 37884 27999
rect 37832 27956 37884 27965
rect 41788 27956 41840 28008
rect 47584 28067 47636 28076
rect 47584 28033 47593 28067
rect 47593 28033 47627 28067
rect 47627 28033 47636 28067
rect 47584 28024 47636 28033
rect 49608 28067 49660 28076
rect 49608 28033 49617 28067
rect 49617 28033 49651 28067
rect 49651 28033 49660 28067
rect 49608 28024 49660 28033
rect 49884 28067 49936 28076
rect 49884 28033 49893 28067
rect 49893 28033 49927 28067
rect 49927 28033 49936 28067
rect 49884 28024 49936 28033
rect 50068 28024 50120 28076
rect 44640 27999 44692 28008
rect 44640 27965 44649 27999
rect 44649 27965 44683 27999
rect 44683 27965 44692 27999
rect 44640 27956 44692 27965
rect 44732 27999 44784 28008
rect 44732 27965 44741 27999
rect 44741 27965 44775 27999
rect 44775 27965 44784 27999
rect 44732 27956 44784 27965
rect 44824 27999 44876 28008
rect 44824 27965 44833 27999
rect 44833 27965 44867 27999
rect 44867 27965 44876 27999
rect 44824 27956 44876 27965
rect 40500 27931 40552 27940
rect 40500 27897 40509 27931
rect 40509 27897 40543 27931
rect 40543 27897 40552 27931
rect 40500 27888 40552 27897
rect 42984 27888 43036 27940
rect 40960 27820 41012 27872
rect 42616 27820 42668 27872
rect 42708 27820 42760 27872
rect 45652 27888 45704 27940
rect 45928 27888 45980 27940
rect 50896 27956 50948 28008
rect 43628 27820 43680 27872
rect 46480 27863 46532 27872
rect 46480 27829 46489 27863
rect 46489 27829 46523 27863
rect 46523 27829 46532 27863
rect 46480 27820 46532 27829
rect 49424 27863 49476 27872
rect 49424 27829 49433 27863
rect 49433 27829 49467 27863
rect 49467 27829 49476 27863
rect 49424 27820 49476 27829
rect 49792 27863 49844 27872
rect 49792 27829 49801 27863
rect 49801 27829 49835 27863
rect 49835 27829 49844 27863
rect 49792 27820 49844 27829
rect 50068 27863 50120 27872
rect 50068 27829 50077 27863
rect 50077 27829 50111 27863
rect 50111 27829 50120 27863
rect 50068 27820 50120 27829
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 43076 27659 43128 27668
rect 43076 27625 43085 27659
rect 43085 27625 43119 27659
rect 43119 27625 43128 27659
rect 43076 27616 43128 27625
rect 40960 27591 41012 27600
rect 40960 27557 40969 27591
rect 40969 27557 41003 27591
rect 41003 27557 41012 27591
rect 40960 27548 41012 27557
rect 42892 27548 42944 27600
rect 43628 27659 43680 27668
rect 43628 27625 43637 27659
rect 43637 27625 43671 27659
rect 43671 27625 43680 27659
rect 43628 27616 43680 27625
rect 43904 27616 43956 27668
rect 44272 27616 44324 27668
rect 44732 27616 44784 27668
rect 46480 27616 46532 27668
rect 47400 27616 47452 27668
rect 48136 27659 48188 27668
rect 48136 27625 48145 27659
rect 48145 27625 48179 27659
rect 48179 27625 48188 27659
rect 48136 27616 48188 27625
rect 52460 27616 52512 27668
rect 40500 27523 40552 27532
rect 40500 27489 40509 27523
rect 40509 27489 40543 27523
rect 40543 27489 40552 27523
rect 40500 27480 40552 27489
rect 41604 27480 41656 27532
rect 30564 27455 30616 27464
rect 30564 27421 30573 27455
rect 30573 27421 30607 27455
rect 30607 27421 30616 27455
rect 30564 27412 30616 27421
rect 30932 27455 30984 27464
rect 30932 27421 30941 27455
rect 30941 27421 30975 27455
rect 30975 27421 30984 27455
rect 30932 27412 30984 27421
rect 32772 27412 32824 27464
rect 37648 27455 37700 27464
rect 37648 27421 37657 27455
rect 37657 27421 37691 27455
rect 37691 27421 37700 27455
rect 37648 27412 37700 27421
rect 41420 27412 41472 27464
rect 29552 27387 29604 27396
rect 29552 27353 29561 27387
rect 29561 27353 29595 27387
rect 29595 27353 29604 27387
rect 29552 27344 29604 27353
rect 32220 27344 32272 27396
rect 32496 27276 32548 27328
rect 34704 27344 34756 27396
rect 36268 27344 36320 27396
rect 33324 27276 33376 27328
rect 34520 27276 34572 27328
rect 36728 27276 36780 27328
rect 39948 27276 40000 27328
rect 40408 27344 40460 27396
rect 41788 27387 41840 27396
rect 41788 27353 41797 27387
rect 41797 27353 41831 27387
rect 41831 27353 41840 27387
rect 41788 27344 41840 27353
rect 42800 27412 42852 27464
rect 42984 27412 43036 27464
rect 43168 27455 43220 27464
rect 43168 27421 43177 27455
rect 43177 27421 43211 27455
rect 43211 27421 43220 27455
rect 43168 27412 43220 27421
rect 43536 27480 43588 27532
rect 43720 27480 43772 27532
rect 44088 27480 44140 27532
rect 48228 27480 48280 27532
rect 49792 27480 49844 27532
rect 50988 27480 51040 27532
rect 51908 27523 51960 27532
rect 51908 27489 51917 27523
rect 51917 27489 51951 27523
rect 51951 27489 51960 27523
rect 51908 27480 51960 27489
rect 43996 27344 44048 27396
rect 46296 27412 46348 27464
rect 49700 27455 49752 27464
rect 49700 27421 49709 27455
rect 49709 27421 49743 27455
rect 49743 27421 49752 27455
rect 49700 27412 49752 27421
rect 47400 27344 47452 27396
rect 50436 27387 50488 27396
rect 50436 27353 50445 27387
rect 50445 27353 50479 27387
rect 50479 27353 50488 27387
rect 50436 27344 50488 27353
rect 50528 27344 50580 27396
rect 41236 27276 41288 27328
rect 45100 27276 45152 27328
rect 47584 27276 47636 27328
rect 52000 27319 52052 27328
rect 52000 27285 52009 27319
rect 52009 27285 52043 27319
rect 52043 27285 52052 27319
rect 52000 27276 52052 27285
rect 4874 27174 4926 27226
rect 4938 27174 4990 27226
rect 5002 27174 5054 27226
rect 5066 27174 5118 27226
rect 5130 27174 5182 27226
rect 35594 27174 35646 27226
rect 35658 27174 35710 27226
rect 35722 27174 35774 27226
rect 35786 27174 35838 27226
rect 35850 27174 35902 27226
rect 28908 27072 28960 27124
rect 30932 27072 30984 27124
rect 32772 27115 32824 27124
rect 32772 27081 32781 27115
rect 32781 27081 32815 27115
rect 32815 27081 32824 27115
rect 32772 27072 32824 27081
rect 32036 26936 32088 26988
rect 32404 26979 32456 26988
rect 32404 26945 32413 26979
rect 32413 26945 32447 26979
rect 32447 26945 32456 26979
rect 32404 26936 32456 26945
rect 32496 26936 32548 26988
rect 32864 26936 32916 26988
rect 32956 26979 33008 26988
rect 32956 26945 32965 26979
rect 32965 26945 32999 26979
rect 32999 26945 33008 26979
rect 32956 26936 33008 26945
rect 33324 26979 33376 26988
rect 33324 26945 33333 26979
rect 33333 26945 33367 26979
rect 33367 26945 33376 26979
rect 33324 26936 33376 26945
rect 22836 26868 22888 26920
rect 23480 26911 23532 26920
rect 23480 26877 23489 26911
rect 23489 26877 23523 26911
rect 23523 26877 23532 26911
rect 23480 26868 23532 26877
rect 24952 26775 25004 26784
rect 24952 26741 24961 26775
rect 24961 26741 24995 26775
rect 24995 26741 25004 26775
rect 24952 26732 25004 26741
rect 25320 26911 25372 26920
rect 25320 26877 25329 26911
rect 25329 26877 25363 26911
rect 25363 26877 25372 26911
rect 25320 26868 25372 26877
rect 25872 26868 25924 26920
rect 25872 26732 25924 26784
rect 26792 26775 26844 26784
rect 26792 26741 26801 26775
rect 26801 26741 26835 26775
rect 26835 26741 26844 26775
rect 26792 26732 26844 26741
rect 27620 26911 27672 26920
rect 27620 26877 27629 26911
rect 27629 26877 27663 26911
rect 27663 26877 27672 26911
rect 27620 26868 27672 26877
rect 33692 26979 33744 26988
rect 33692 26945 33701 26979
rect 33701 26945 33735 26979
rect 33735 26945 33744 26979
rect 33692 26936 33744 26945
rect 34520 27072 34572 27124
rect 35992 27072 36044 27124
rect 36268 27004 36320 27056
rect 36544 27072 36596 27124
rect 37832 27072 37884 27124
rect 34612 26868 34664 26920
rect 34888 26979 34940 26988
rect 34888 26945 34897 26979
rect 34897 26945 34931 26979
rect 34931 26945 34940 26979
rect 34888 26936 34940 26945
rect 34520 26800 34572 26852
rect 34888 26800 34940 26852
rect 28356 26732 28408 26784
rect 28632 26732 28684 26784
rect 32864 26732 32916 26784
rect 34796 26732 34848 26784
rect 36636 26911 36688 26920
rect 36636 26877 36645 26911
rect 36645 26877 36679 26911
rect 36679 26877 36688 26911
rect 36636 26868 36688 26877
rect 36820 26868 36872 26920
rect 37648 26936 37700 26988
rect 36084 26732 36136 26784
rect 39948 27115 40000 27124
rect 39948 27081 39957 27115
rect 39957 27081 39991 27115
rect 39991 27081 40000 27115
rect 39948 27072 40000 27081
rect 42800 27072 42852 27124
rect 43812 27115 43864 27124
rect 43812 27081 43821 27115
rect 43821 27081 43855 27115
rect 43855 27081 43864 27115
rect 43812 27072 43864 27081
rect 49884 27072 49936 27124
rect 50436 27072 50488 27124
rect 52460 27115 52512 27124
rect 52460 27081 52469 27115
rect 52469 27081 52503 27115
rect 52503 27081 52512 27115
rect 52460 27072 52512 27081
rect 40224 26936 40276 26988
rect 41052 26936 41104 26988
rect 41236 26979 41288 26988
rect 41236 26945 41245 26979
rect 41245 26945 41279 26979
rect 41279 26945 41288 26979
rect 41236 26936 41288 26945
rect 41788 26936 41840 26988
rect 40408 26868 40460 26920
rect 41604 26868 41656 26920
rect 42340 26868 42392 26920
rect 42708 26868 42760 26920
rect 43628 26979 43680 26988
rect 43628 26945 43637 26979
rect 43637 26945 43671 26979
rect 43671 26945 43680 26979
rect 43628 26936 43680 26945
rect 43904 26979 43956 26988
rect 43904 26945 43913 26979
rect 43913 26945 43947 26979
rect 43947 26945 43956 26979
rect 43904 26936 43956 26945
rect 49424 27004 49476 27056
rect 53288 27004 53340 27056
rect 48320 26868 48372 26920
rect 48688 26911 48740 26920
rect 48688 26877 48697 26911
rect 48697 26877 48731 26911
rect 48731 26877 48740 26911
rect 48688 26868 48740 26877
rect 48228 26800 48280 26852
rect 40500 26732 40552 26784
rect 42708 26732 42760 26784
rect 43628 26775 43680 26784
rect 43628 26741 43637 26775
rect 43637 26741 43671 26775
rect 43671 26741 43680 26775
rect 43628 26732 43680 26741
rect 46848 26775 46900 26784
rect 46848 26741 46857 26775
rect 46857 26741 46891 26775
rect 46891 26741 46900 26775
rect 46848 26732 46900 26741
rect 49148 26868 49200 26920
rect 50528 26936 50580 26988
rect 50804 26936 50856 26988
rect 52000 26936 52052 26988
rect 50620 26911 50672 26920
rect 50620 26877 50629 26911
rect 50629 26877 50663 26911
rect 50663 26877 50672 26911
rect 50620 26868 50672 26877
rect 49700 26732 49752 26784
rect 52184 26800 52236 26852
rect 53012 26911 53064 26920
rect 53012 26877 53021 26911
rect 53021 26877 53055 26911
rect 53055 26877 53064 26911
rect 53012 26868 53064 26877
rect 50988 26732 51040 26784
rect 54484 26775 54536 26784
rect 54484 26741 54493 26775
rect 54493 26741 54527 26775
rect 54527 26741 54536 26775
rect 54484 26732 54536 26741
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 23480 26528 23532 26580
rect 25228 26528 25280 26580
rect 25228 26392 25280 26444
rect 24768 26367 24820 26376
rect 24768 26333 24777 26367
rect 24777 26333 24811 26367
rect 24811 26333 24820 26367
rect 24768 26324 24820 26333
rect 24952 26324 25004 26376
rect 25320 26367 25372 26376
rect 25320 26333 25329 26367
rect 25329 26333 25363 26367
rect 25363 26333 25372 26367
rect 25320 26324 25372 26333
rect 27988 26460 28040 26512
rect 25504 26392 25556 26444
rect 25964 26367 26016 26376
rect 25964 26333 25973 26367
rect 25973 26333 26007 26367
rect 26007 26333 26016 26367
rect 25964 26324 26016 26333
rect 26332 26367 26384 26376
rect 26332 26333 26341 26367
rect 26341 26333 26375 26367
rect 26375 26333 26384 26367
rect 27804 26392 27856 26444
rect 26332 26324 26384 26333
rect 22744 26231 22796 26240
rect 22744 26197 22753 26231
rect 22753 26197 22787 26231
rect 22787 26197 22796 26231
rect 22744 26188 22796 26197
rect 24860 26188 24912 26240
rect 25228 26188 25280 26240
rect 26240 26256 26292 26308
rect 26792 26256 26844 26308
rect 27712 26367 27764 26376
rect 27712 26333 27721 26367
rect 27721 26333 27755 26367
rect 27755 26333 27764 26367
rect 27712 26324 27764 26333
rect 29092 26528 29144 26580
rect 30196 26528 30248 26580
rect 32404 26528 32456 26580
rect 34704 26528 34756 26580
rect 35164 26528 35216 26580
rect 35808 26528 35860 26580
rect 32864 26460 32916 26512
rect 33692 26460 33744 26512
rect 29920 26392 29972 26444
rect 30196 26435 30248 26444
rect 30196 26401 30205 26435
rect 30205 26401 30239 26435
rect 30239 26401 30248 26435
rect 30196 26392 30248 26401
rect 28816 26367 28868 26376
rect 28816 26333 28825 26367
rect 28825 26333 28859 26367
rect 28859 26333 28868 26367
rect 28816 26324 28868 26333
rect 32496 26367 32548 26376
rect 32496 26333 32505 26367
rect 32505 26333 32539 26367
rect 32539 26333 32548 26367
rect 32496 26324 32548 26333
rect 33324 26392 33376 26444
rect 34520 26392 34572 26444
rect 34704 26392 34756 26444
rect 34796 26392 34848 26444
rect 33048 26324 33100 26376
rect 33140 26324 33192 26376
rect 34428 26324 34480 26376
rect 35072 26367 35124 26376
rect 35072 26333 35081 26367
rect 35081 26333 35115 26367
rect 35115 26333 35124 26367
rect 35072 26324 35124 26333
rect 35900 26460 35952 26512
rect 36636 26528 36688 26580
rect 38936 26571 38988 26580
rect 38936 26537 38945 26571
rect 38945 26537 38979 26571
rect 38979 26537 38988 26571
rect 38936 26528 38988 26537
rect 40224 26571 40276 26580
rect 40224 26537 40233 26571
rect 40233 26537 40267 26571
rect 40267 26537 40276 26571
rect 40224 26528 40276 26537
rect 40500 26528 40552 26580
rect 44180 26528 44232 26580
rect 48688 26528 48740 26580
rect 49608 26528 49660 26580
rect 27712 26188 27764 26240
rect 28356 26256 28408 26308
rect 30564 26256 30616 26308
rect 32404 26256 32456 26308
rect 35624 26324 35676 26376
rect 35900 26367 35952 26376
rect 35900 26333 35909 26367
rect 35909 26333 35943 26367
rect 35943 26333 35952 26367
rect 35900 26324 35952 26333
rect 36728 26460 36780 26512
rect 39028 26460 39080 26512
rect 40132 26460 40184 26512
rect 36360 26367 36412 26376
rect 36360 26333 36369 26367
rect 36369 26333 36403 26367
rect 36403 26333 36412 26367
rect 36360 26324 36412 26333
rect 36452 26367 36504 26376
rect 36452 26333 36461 26367
rect 36461 26333 36495 26367
rect 36495 26333 36504 26367
rect 36452 26324 36504 26333
rect 28540 26231 28592 26240
rect 28540 26197 28549 26231
rect 28549 26197 28583 26231
rect 28583 26197 28592 26231
rect 28540 26188 28592 26197
rect 30932 26188 30984 26240
rect 33232 26188 33284 26240
rect 35256 26188 35308 26240
rect 35532 26188 35584 26240
rect 36268 26256 36320 26308
rect 36176 26188 36228 26240
rect 38660 26392 38712 26444
rect 42892 26460 42944 26512
rect 43444 26460 43496 26512
rect 45836 26460 45888 26512
rect 37188 26324 37240 26376
rect 39304 26231 39356 26240
rect 39304 26197 39313 26231
rect 39313 26197 39347 26231
rect 39347 26197 39356 26231
rect 39304 26188 39356 26197
rect 39948 26324 40000 26376
rect 40500 26324 40552 26376
rect 39488 26188 39540 26240
rect 40040 26231 40092 26240
rect 40040 26197 40049 26231
rect 40049 26197 40083 26231
rect 40083 26197 40092 26231
rect 40040 26188 40092 26197
rect 40224 26188 40276 26240
rect 42064 26392 42116 26444
rect 42432 26392 42484 26444
rect 45560 26392 45612 26444
rect 46296 26392 46348 26444
rect 46848 26435 46900 26444
rect 46848 26401 46857 26435
rect 46857 26401 46891 26435
rect 46891 26401 46900 26435
rect 46848 26392 46900 26401
rect 48044 26392 48096 26444
rect 49516 26460 49568 26512
rect 42892 26324 42944 26376
rect 43352 26256 43404 26308
rect 44916 26256 44968 26308
rect 48688 26324 48740 26376
rect 42156 26188 42208 26240
rect 43628 26188 43680 26240
rect 45928 26188 45980 26240
rect 47124 26256 47176 26308
rect 48136 26256 48188 26308
rect 48780 26256 48832 26308
rect 49148 26256 49200 26308
rect 49516 26367 49568 26376
rect 49516 26333 49520 26367
rect 49520 26333 49554 26367
rect 49554 26333 49568 26367
rect 50804 26571 50856 26580
rect 50804 26537 50813 26571
rect 50813 26537 50847 26571
rect 50847 26537 50856 26571
rect 50804 26528 50856 26537
rect 53012 26528 53064 26580
rect 50620 26460 50672 26512
rect 51908 26460 51960 26512
rect 57888 26460 57940 26512
rect 50436 26392 50488 26444
rect 49516 26324 49568 26333
rect 49976 26367 50028 26376
rect 49976 26333 49985 26367
rect 49985 26333 50019 26367
rect 50019 26333 50028 26367
rect 49976 26324 50028 26333
rect 49332 26256 49384 26308
rect 49700 26299 49752 26308
rect 49700 26265 49709 26299
rect 49709 26265 49743 26299
rect 49743 26265 49752 26299
rect 49700 26256 49752 26265
rect 49792 26256 49844 26308
rect 50528 26367 50580 26376
rect 50528 26333 50537 26367
rect 50537 26333 50571 26367
rect 50571 26333 50580 26367
rect 50528 26324 50580 26333
rect 50988 26392 51040 26444
rect 52644 26367 52696 26376
rect 52644 26333 52653 26367
rect 52653 26333 52687 26367
rect 52687 26333 52696 26367
rect 52644 26324 52696 26333
rect 48228 26188 48280 26240
rect 49056 26188 49108 26240
rect 49976 26188 50028 26240
rect 50436 26299 50488 26308
rect 50436 26265 50445 26299
rect 50445 26265 50479 26299
rect 50479 26265 50488 26299
rect 50436 26256 50488 26265
rect 54484 26324 54536 26376
rect 58256 26367 58308 26376
rect 58256 26333 58265 26367
rect 58265 26333 58299 26367
rect 58299 26333 58308 26367
rect 58256 26324 58308 26333
rect 53012 26188 53064 26240
rect 4874 26086 4926 26138
rect 4938 26086 4990 26138
rect 5002 26086 5054 26138
rect 5066 26086 5118 26138
rect 5130 26086 5182 26138
rect 35594 26086 35646 26138
rect 35658 26086 35710 26138
rect 35722 26086 35774 26138
rect 35786 26086 35838 26138
rect 35850 26086 35902 26138
rect 22284 25984 22336 26036
rect 22744 25984 22796 26036
rect 20168 25916 20220 25968
rect 19616 25848 19668 25900
rect 19800 25780 19852 25832
rect 20536 25780 20588 25832
rect 22376 25848 22428 25900
rect 22744 25848 22796 25900
rect 23296 25848 23348 25900
rect 23480 25848 23532 25900
rect 24124 25848 24176 25900
rect 25044 25848 25096 25900
rect 23020 25780 23072 25832
rect 23388 25780 23440 25832
rect 25228 25891 25280 25900
rect 25228 25857 25237 25891
rect 25237 25857 25271 25891
rect 25271 25857 25280 25891
rect 25228 25848 25280 25857
rect 26516 25916 26568 25968
rect 27804 25916 27856 25968
rect 27620 25848 27672 25900
rect 18236 25644 18288 25696
rect 21180 25644 21232 25696
rect 22008 25644 22060 25696
rect 24768 25712 24820 25764
rect 24860 25755 24912 25764
rect 24860 25721 24869 25755
rect 24869 25721 24903 25755
rect 24903 25721 24912 25755
rect 24860 25712 24912 25721
rect 26240 25780 26292 25832
rect 26976 25780 27028 25832
rect 27988 25891 28040 25900
rect 27988 25857 27997 25891
rect 27997 25857 28031 25891
rect 28031 25857 28040 25891
rect 27988 25848 28040 25857
rect 28540 25916 28592 25968
rect 28908 25916 28960 25968
rect 30196 25984 30248 26036
rect 32956 25916 33008 25968
rect 35532 25984 35584 26036
rect 35624 25916 35676 25968
rect 37648 25984 37700 26036
rect 36912 25916 36964 25968
rect 38936 25916 38988 25968
rect 40040 25984 40092 26036
rect 42524 25984 42576 26036
rect 40868 25916 40920 25968
rect 42708 25959 42760 25968
rect 42708 25925 42717 25959
rect 42717 25925 42751 25959
rect 42751 25925 42760 25959
rect 42708 25916 42760 25925
rect 42892 26027 42944 26036
rect 42892 25993 42917 26027
rect 42917 25993 42944 26027
rect 42892 25984 42944 25993
rect 43812 25959 43864 25968
rect 43812 25925 43821 25959
rect 43821 25925 43855 25959
rect 43855 25925 43864 25959
rect 43812 25916 43864 25925
rect 28356 25891 28408 25900
rect 28356 25857 28365 25891
rect 28365 25857 28399 25891
rect 28399 25857 28408 25891
rect 28356 25848 28408 25857
rect 32128 25891 32180 25900
rect 32128 25857 32137 25891
rect 32137 25857 32171 25891
rect 32171 25857 32180 25891
rect 32128 25848 32180 25857
rect 32588 25848 32640 25900
rect 35164 25848 35216 25900
rect 28632 25780 28684 25832
rect 32404 25780 32456 25832
rect 35256 25780 35308 25832
rect 35532 25780 35584 25832
rect 35808 25891 35860 25900
rect 35808 25857 35817 25891
rect 35817 25857 35851 25891
rect 35851 25857 35860 25891
rect 35808 25848 35860 25857
rect 36084 25891 36136 25900
rect 36084 25857 36093 25891
rect 36093 25857 36127 25891
rect 36127 25857 36136 25891
rect 36084 25848 36136 25857
rect 37188 25848 37240 25900
rect 39304 25848 39356 25900
rect 39672 25891 39724 25900
rect 39672 25857 39681 25891
rect 39681 25857 39715 25891
rect 39715 25857 39724 25891
rect 39672 25848 39724 25857
rect 36728 25780 36780 25832
rect 25320 25712 25372 25764
rect 39396 25780 39448 25832
rect 39488 25823 39540 25832
rect 39488 25789 39497 25823
rect 39497 25789 39531 25823
rect 39531 25789 39540 25823
rect 39488 25780 39540 25789
rect 42340 25848 42392 25900
rect 39948 25823 40000 25832
rect 39948 25789 39957 25823
rect 39957 25789 39991 25823
rect 39991 25789 40000 25823
rect 39948 25780 40000 25789
rect 40316 25780 40368 25832
rect 41972 25780 42024 25832
rect 25412 25644 25464 25696
rect 25504 25644 25556 25696
rect 26148 25644 26200 25696
rect 28724 25644 28776 25696
rect 31760 25644 31812 25696
rect 33324 25644 33376 25696
rect 35532 25687 35584 25696
rect 35532 25653 35541 25687
rect 35541 25653 35575 25687
rect 35575 25653 35584 25687
rect 35532 25644 35584 25653
rect 35624 25644 35676 25696
rect 37740 25644 37792 25696
rect 38752 25644 38804 25696
rect 39856 25712 39908 25764
rect 39396 25687 39448 25696
rect 39396 25653 39405 25687
rect 39405 25653 39439 25687
rect 39439 25653 39448 25687
rect 39396 25644 39448 25653
rect 40592 25644 40644 25696
rect 42616 25644 42668 25696
rect 43444 25823 43496 25832
rect 43444 25789 43453 25823
rect 43453 25789 43487 25823
rect 43487 25789 43496 25823
rect 44180 25891 44232 25900
rect 44180 25857 44189 25891
rect 44189 25857 44223 25891
rect 44223 25857 44232 25891
rect 45744 25984 45796 26036
rect 47124 25984 47176 26036
rect 48320 26027 48372 26036
rect 48320 25993 48329 26027
rect 48329 25993 48363 26027
rect 48363 25993 48372 26027
rect 48320 25984 48372 25993
rect 45928 25916 45980 25968
rect 47216 25916 47268 25968
rect 48136 25916 48188 25968
rect 49700 25984 49752 26036
rect 50436 25984 50488 26036
rect 44180 25848 44232 25857
rect 47952 25848 48004 25900
rect 43444 25780 43496 25789
rect 45560 25823 45612 25832
rect 45560 25789 45569 25823
rect 45569 25789 45603 25823
rect 45603 25789 45612 25823
rect 45560 25780 45612 25789
rect 47308 25823 47360 25832
rect 47308 25789 47317 25823
rect 47317 25789 47351 25823
rect 47351 25789 47360 25823
rect 47308 25780 47360 25789
rect 48688 25891 48740 25900
rect 48688 25857 48697 25891
rect 48697 25857 48731 25891
rect 48731 25857 48740 25891
rect 48688 25848 48740 25857
rect 50528 25916 50580 25968
rect 52644 25984 52696 26036
rect 51908 25959 51960 25968
rect 51908 25925 51917 25959
rect 51917 25925 51951 25959
rect 51951 25925 51960 25959
rect 51908 25916 51960 25925
rect 53012 25959 53064 25968
rect 53012 25925 53021 25959
rect 53021 25925 53055 25959
rect 53055 25925 53064 25959
rect 53012 25916 53064 25925
rect 54208 25916 54260 25968
rect 49516 25848 49568 25900
rect 50344 25848 50396 25900
rect 51356 25848 51408 25900
rect 51632 25891 51684 25900
rect 51632 25857 51642 25891
rect 51642 25857 51676 25891
rect 51676 25857 51684 25891
rect 51632 25848 51684 25857
rect 52644 25848 52696 25900
rect 49148 25780 49200 25832
rect 49792 25780 49844 25832
rect 50160 25823 50212 25832
rect 50160 25789 50169 25823
rect 50169 25789 50203 25823
rect 50203 25789 50212 25823
rect 50160 25780 50212 25789
rect 50712 25780 50764 25832
rect 53472 25848 53524 25900
rect 53748 25848 53800 25900
rect 56692 25891 56744 25900
rect 56692 25857 56701 25891
rect 56701 25857 56735 25891
rect 56735 25857 56744 25891
rect 56692 25848 56744 25857
rect 56876 25891 56928 25900
rect 56876 25857 56885 25891
rect 56885 25857 56919 25891
rect 56919 25857 56928 25891
rect 56876 25848 56928 25857
rect 55312 25780 55364 25832
rect 55956 25823 56008 25832
rect 55956 25789 55965 25823
rect 55965 25789 55999 25823
rect 55999 25789 56008 25823
rect 55956 25780 56008 25789
rect 56232 25823 56284 25832
rect 56232 25789 56241 25823
rect 56241 25789 56275 25823
rect 56275 25789 56284 25823
rect 56232 25780 56284 25789
rect 43812 25644 43864 25696
rect 44272 25644 44324 25696
rect 44456 25644 44508 25696
rect 49608 25712 49660 25764
rect 50436 25755 50488 25764
rect 50436 25721 50445 25755
rect 50445 25721 50479 25755
rect 50479 25721 50488 25755
rect 50436 25712 50488 25721
rect 58256 25780 58308 25832
rect 49976 25687 50028 25696
rect 49976 25653 49985 25687
rect 49985 25653 50019 25687
rect 50019 25653 50028 25687
rect 49976 25644 50028 25653
rect 51356 25687 51408 25696
rect 51356 25653 51365 25687
rect 51365 25653 51399 25687
rect 51399 25653 51408 25687
rect 51356 25644 51408 25653
rect 51816 25644 51868 25696
rect 56508 25687 56560 25696
rect 56508 25653 56517 25687
rect 56517 25653 56551 25687
rect 56551 25653 56560 25687
rect 56508 25644 56560 25653
rect 57520 25687 57572 25696
rect 57520 25653 57529 25687
rect 57529 25653 57563 25687
rect 57563 25653 57572 25687
rect 57520 25644 57572 25653
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 21548 25440 21600 25492
rect 22192 25440 22244 25492
rect 22376 25440 22428 25492
rect 23296 25483 23348 25492
rect 23296 25449 23305 25483
rect 23305 25449 23339 25483
rect 23339 25449 23348 25483
rect 23296 25440 23348 25449
rect 17960 25304 18012 25356
rect 19524 25279 19576 25288
rect 19524 25245 19533 25279
rect 19533 25245 19567 25279
rect 19567 25245 19576 25279
rect 19524 25236 19576 25245
rect 19432 25168 19484 25220
rect 19616 25211 19668 25220
rect 19616 25177 19625 25211
rect 19625 25177 19659 25211
rect 19659 25177 19668 25211
rect 19616 25168 19668 25177
rect 19708 25211 19760 25220
rect 19708 25177 19717 25211
rect 19717 25177 19751 25211
rect 19751 25177 19760 25211
rect 19708 25168 19760 25177
rect 20168 25279 20220 25288
rect 20168 25245 20177 25279
rect 20177 25245 20211 25279
rect 20211 25245 20220 25279
rect 20168 25236 20220 25245
rect 21824 25304 21876 25356
rect 23388 25304 23440 25356
rect 20536 25279 20588 25288
rect 20536 25245 20545 25279
rect 20545 25245 20579 25279
rect 20579 25245 20588 25279
rect 20536 25236 20588 25245
rect 20904 25279 20956 25288
rect 20904 25245 20913 25279
rect 20913 25245 20947 25279
rect 20947 25245 20956 25279
rect 20904 25236 20956 25245
rect 21180 25279 21232 25288
rect 21180 25245 21189 25279
rect 21189 25245 21223 25279
rect 21223 25245 21232 25279
rect 21180 25236 21232 25245
rect 23296 25236 23348 25288
rect 23480 25279 23532 25288
rect 23480 25245 23484 25279
rect 23484 25245 23518 25279
rect 23518 25245 23532 25279
rect 23480 25236 23532 25245
rect 22008 25168 22060 25220
rect 23020 25168 23072 25220
rect 23572 25211 23624 25220
rect 23572 25177 23581 25211
rect 23581 25177 23615 25211
rect 23615 25177 23624 25211
rect 23572 25168 23624 25177
rect 25044 25372 25096 25424
rect 25228 25372 25280 25424
rect 24952 25304 25004 25356
rect 25688 25304 25740 25356
rect 22376 25100 22428 25152
rect 23296 25100 23348 25152
rect 25228 25236 25280 25288
rect 26240 25372 26292 25424
rect 28816 25440 28868 25492
rect 31852 25440 31904 25492
rect 34336 25440 34388 25492
rect 36268 25440 36320 25492
rect 30196 25372 30248 25424
rect 32864 25372 32916 25424
rect 25412 25168 25464 25220
rect 28356 25279 28408 25288
rect 28356 25245 28365 25279
rect 28365 25245 28399 25279
rect 28399 25245 28408 25279
rect 28356 25236 28408 25245
rect 28448 25236 28500 25288
rect 28816 25236 28868 25288
rect 24216 25100 24268 25152
rect 26056 25100 26108 25152
rect 27712 25168 27764 25220
rect 28632 25211 28684 25220
rect 28632 25177 28641 25211
rect 28641 25177 28675 25211
rect 28675 25177 28684 25211
rect 28632 25168 28684 25177
rect 27344 25100 27396 25152
rect 28172 25100 28224 25152
rect 30564 25304 30616 25356
rect 34980 25304 35032 25356
rect 36820 25304 36872 25356
rect 37464 25372 37516 25424
rect 33232 25279 33284 25288
rect 33232 25245 33241 25279
rect 33241 25245 33275 25279
rect 33275 25245 33284 25279
rect 33232 25236 33284 25245
rect 33324 25279 33376 25288
rect 33324 25245 33333 25279
rect 33333 25245 33367 25279
rect 33367 25245 33376 25279
rect 33324 25236 33376 25245
rect 32220 25168 32272 25220
rect 33048 25168 33100 25220
rect 35072 25279 35124 25288
rect 35072 25245 35081 25279
rect 35081 25245 35115 25279
rect 35115 25245 35124 25279
rect 35072 25236 35124 25245
rect 35992 25236 36044 25288
rect 37096 25304 37148 25356
rect 37740 25347 37792 25356
rect 37740 25313 37749 25347
rect 37749 25313 37783 25347
rect 37783 25313 37792 25347
rect 37740 25304 37792 25313
rect 37004 25279 37056 25288
rect 37004 25245 37013 25279
rect 37013 25245 37047 25279
rect 37047 25245 37056 25279
rect 37004 25236 37056 25245
rect 37188 25236 37240 25288
rect 36084 25168 36136 25220
rect 36544 25168 36596 25220
rect 36820 25211 36872 25220
rect 36820 25177 36829 25211
rect 36829 25177 36863 25211
rect 36863 25177 36872 25211
rect 36820 25168 36872 25177
rect 37648 25168 37700 25220
rect 38936 25440 38988 25492
rect 40224 25440 40276 25492
rect 41512 25440 41564 25492
rect 42708 25440 42760 25492
rect 38844 25372 38896 25424
rect 39488 25304 39540 25356
rect 38660 25279 38712 25288
rect 38660 25245 38664 25279
rect 38664 25245 38698 25279
rect 38698 25245 38712 25279
rect 38660 25236 38712 25245
rect 38752 25279 38804 25288
rect 38752 25245 38761 25279
rect 38761 25245 38795 25279
rect 38795 25245 38804 25279
rect 38752 25236 38804 25245
rect 39028 25279 39080 25288
rect 39028 25245 39036 25279
rect 39036 25245 39070 25279
rect 39070 25245 39080 25279
rect 39028 25236 39080 25245
rect 39120 25279 39172 25288
rect 39120 25245 39129 25279
rect 39129 25245 39163 25279
rect 39163 25245 39172 25279
rect 39120 25236 39172 25245
rect 31760 25100 31812 25152
rect 32036 25100 32088 25152
rect 33232 25100 33284 25152
rect 37004 25100 37056 25152
rect 37556 25100 37608 25152
rect 38476 25143 38528 25152
rect 38476 25109 38485 25143
rect 38485 25109 38519 25143
rect 38519 25109 38528 25143
rect 38476 25100 38528 25109
rect 38844 25211 38896 25220
rect 38844 25177 38853 25211
rect 38853 25177 38887 25211
rect 38887 25177 38896 25211
rect 38844 25168 38896 25177
rect 39396 25236 39448 25288
rect 39856 25236 39908 25288
rect 40040 25279 40092 25288
rect 40040 25245 40058 25279
rect 40058 25245 40092 25279
rect 40040 25236 40092 25245
rect 40316 25304 40368 25356
rect 41236 25304 41288 25356
rect 41972 25347 42024 25356
rect 41972 25313 41981 25347
rect 41981 25313 42015 25347
rect 42015 25313 42024 25347
rect 41972 25304 42024 25313
rect 42064 25347 42116 25356
rect 42064 25313 42073 25347
rect 42073 25313 42107 25347
rect 42107 25313 42116 25347
rect 42064 25304 42116 25313
rect 42340 25304 42392 25356
rect 42800 25372 42852 25424
rect 43352 25483 43404 25492
rect 43352 25449 43361 25483
rect 43361 25449 43395 25483
rect 43395 25449 43404 25483
rect 43352 25440 43404 25449
rect 43812 25483 43864 25492
rect 43812 25449 43821 25483
rect 43821 25449 43855 25483
rect 43855 25449 43864 25483
rect 43812 25440 43864 25449
rect 43996 25440 44048 25492
rect 44456 25372 44508 25424
rect 48228 25483 48280 25492
rect 48228 25449 48237 25483
rect 48237 25449 48271 25483
rect 48271 25449 48280 25483
rect 48228 25440 48280 25449
rect 50160 25483 50212 25492
rect 50160 25449 50169 25483
rect 50169 25449 50203 25483
rect 50203 25449 50212 25483
rect 50160 25440 50212 25449
rect 52644 25440 52696 25492
rect 39672 25168 39724 25220
rect 39304 25100 39356 25152
rect 40960 25100 41012 25152
rect 41420 25211 41472 25220
rect 41420 25177 41429 25211
rect 41429 25177 41463 25211
rect 41463 25177 41472 25211
rect 41420 25168 41472 25177
rect 42524 25236 42576 25288
rect 42892 25236 42944 25288
rect 43812 25304 43864 25356
rect 43628 25279 43680 25288
rect 43628 25245 43637 25279
rect 43637 25245 43671 25279
rect 43671 25245 43680 25279
rect 43628 25236 43680 25245
rect 42616 25168 42668 25220
rect 42708 25211 42760 25220
rect 42708 25177 42717 25211
rect 42717 25177 42751 25211
rect 42751 25177 42760 25211
rect 42708 25168 42760 25177
rect 41512 25100 41564 25152
rect 43996 25100 44048 25152
rect 46480 25304 46532 25356
rect 47952 25304 48004 25356
rect 50252 25372 50304 25424
rect 45652 25279 45704 25288
rect 45652 25245 45661 25279
rect 45661 25245 45695 25279
rect 45695 25245 45704 25279
rect 45652 25236 45704 25245
rect 45928 25211 45980 25220
rect 45928 25177 45937 25211
rect 45937 25177 45971 25211
rect 45971 25177 45980 25211
rect 45928 25168 45980 25177
rect 47216 25168 47268 25220
rect 47492 25168 47544 25220
rect 48964 25236 49016 25288
rect 49148 25236 49200 25288
rect 49332 25279 49384 25288
rect 49332 25245 49341 25279
rect 49341 25245 49375 25279
rect 49375 25245 49384 25279
rect 49332 25236 49384 25245
rect 49424 25279 49476 25288
rect 49424 25245 49433 25279
rect 49433 25245 49467 25279
rect 49467 25245 49476 25279
rect 49424 25236 49476 25245
rect 50160 25236 50212 25288
rect 50620 25236 50672 25288
rect 50712 25279 50764 25288
rect 50712 25245 50720 25279
rect 50720 25245 50754 25279
rect 50754 25245 50764 25279
rect 50712 25236 50764 25245
rect 52184 25347 52236 25356
rect 52184 25313 52193 25347
rect 52193 25313 52227 25347
rect 52227 25313 52236 25347
rect 52184 25304 52236 25313
rect 52828 25304 52880 25356
rect 53472 25304 53524 25356
rect 51816 25279 51868 25288
rect 51816 25245 51825 25279
rect 51825 25245 51859 25279
rect 51859 25245 51868 25279
rect 51816 25236 51868 25245
rect 52000 25279 52052 25288
rect 52000 25245 52009 25279
rect 52009 25245 52043 25279
rect 52043 25245 52052 25279
rect 52000 25236 52052 25245
rect 55956 25440 56008 25492
rect 58256 25483 58308 25492
rect 58256 25449 58265 25483
rect 58265 25449 58299 25483
rect 58299 25449 58308 25483
rect 58256 25440 58308 25449
rect 56232 25372 56284 25424
rect 48596 25211 48648 25220
rect 48596 25177 48605 25211
rect 48605 25177 48639 25211
rect 48639 25177 48648 25211
rect 48596 25168 48648 25177
rect 46940 25100 46992 25152
rect 47768 25100 47820 25152
rect 48780 25100 48832 25152
rect 49792 25100 49844 25152
rect 53748 25168 53800 25220
rect 53840 25168 53892 25220
rect 54208 25168 54260 25220
rect 55312 25279 55364 25288
rect 55312 25245 55321 25279
rect 55321 25245 55355 25279
rect 55355 25245 55364 25279
rect 55312 25236 55364 25245
rect 56416 25279 56468 25288
rect 56416 25245 56425 25279
rect 56425 25245 56459 25279
rect 56459 25245 56468 25279
rect 56416 25236 56468 25245
rect 50804 25100 50856 25152
rect 53380 25100 53432 25152
rect 55680 25168 55732 25220
rect 57520 25236 57572 25288
rect 4874 24998 4926 25050
rect 4938 24998 4990 25050
rect 5002 24998 5054 25050
rect 5066 24998 5118 25050
rect 5130 24998 5182 25050
rect 35594 24998 35646 25050
rect 35658 24998 35710 25050
rect 35722 24998 35774 25050
rect 35786 24998 35838 25050
rect 35850 24998 35902 25050
rect 19800 24939 19852 24948
rect 19800 24905 19809 24939
rect 19809 24905 19843 24939
rect 19843 24905 19852 24939
rect 19800 24896 19852 24905
rect 20904 24896 20956 24948
rect 23572 24896 23624 24948
rect 18236 24871 18288 24880
rect 18236 24837 18245 24871
rect 18245 24837 18279 24871
rect 18279 24837 18288 24871
rect 18236 24828 18288 24837
rect 19708 24828 19760 24880
rect 19892 24828 19944 24880
rect 22376 24828 22428 24880
rect 22560 24828 22612 24880
rect 17960 24803 18012 24812
rect 17960 24769 17969 24803
rect 17969 24769 18003 24803
rect 18003 24769 18012 24803
rect 17960 24760 18012 24769
rect 20076 24803 20128 24812
rect 20076 24769 20085 24803
rect 20085 24769 20119 24803
rect 20119 24769 20128 24803
rect 20076 24760 20128 24769
rect 20536 24760 20588 24812
rect 26332 24896 26384 24948
rect 25596 24828 25648 24880
rect 25688 24828 25740 24880
rect 21732 24692 21784 24744
rect 21824 24735 21876 24744
rect 21824 24701 21833 24735
rect 21833 24701 21867 24735
rect 21867 24701 21876 24735
rect 21824 24692 21876 24701
rect 22836 24692 22888 24744
rect 19616 24624 19668 24676
rect 20628 24624 20680 24676
rect 20812 24624 20864 24676
rect 20444 24599 20496 24608
rect 20444 24565 20453 24599
rect 20453 24565 20487 24599
rect 20487 24565 20496 24599
rect 20444 24556 20496 24565
rect 23112 24624 23164 24676
rect 25320 24803 25372 24812
rect 25320 24769 25329 24803
rect 25329 24769 25363 24803
rect 25363 24769 25372 24803
rect 25320 24760 25372 24769
rect 30196 24896 30248 24948
rect 31852 24896 31904 24948
rect 31484 24828 31536 24880
rect 25412 24624 25464 24676
rect 23296 24556 23348 24608
rect 23572 24599 23624 24608
rect 23572 24565 23581 24599
rect 23581 24565 23615 24599
rect 23615 24565 23624 24599
rect 23572 24556 23624 24565
rect 25320 24556 25372 24608
rect 25504 24599 25556 24608
rect 25504 24565 25513 24599
rect 25513 24565 25547 24599
rect 25547 24565 25556 24599
rect 25504 24556 25556 24565
rect 25964 24760 26016 24812
rect 26056 24803 26108 24812
rect 26056 24769 26065 24803
rect 26065 24769 26099 24803
rect 26099 24769 26108 24803
rect 26056 24760 26108 24769
rect 27436 24760 27488 24812
rect 28908 24760 28960 24812
rect 32036 24828 32088 24880
rect 27528 24735 27580 24744
rect 27528 24701 27537 24735
rect 27537 24701 27571 24735
rect 27571 24701 27580 24735
rect 27528 24692 27580 24701
rect 27804 24735 27856 24744
rect 27804 24701 27813 24735
rect 27813 24701 27847 24735
rect 27847 24701 27856 24735
rect 27804 24692 27856 24701
rect 28356 24692 28408 24744
rect 31852 24760 31904 24812
rect 33048 24828 33100 24880
rect 33140 24828 33192 24880
rect 35440 24828 35492 24880
rect 32496 24803 32548 24812
rect 32496 24769 32505 24803
rect 32505 24769 32539 24803
rect 32539 24769 32548 24803
rect 32496 24760 32548 24769
rect 32680 24803 32732 24812
rect 32680 24769 32689 24803
rect 32689 24769 32723 24803
rect 32723 24769 32732 24803
rect 32680 24760 32732 24769
rect 32588 24692 32640 24744
rect 33416 24760 33468 24812
rect 34980 24803 35032 24812
rect 34980 24769 34989 24803
rect 34989 24769 35023 24803
rect 35023 24769 35032 24803
rect 34980 24760 35032 24769
rect 35072 24760 35124 24812
rect 33232 24692 33284 24744
rect 34428 24692 34480 24744
rect 35716 24760 35768 24812
rect 38016 24871 38068 24880
rect 38016 24837 38043 24871
rect 38043 24837 38068 24871
rect 38016 24828 38068 24837
rect 42432 24896 42484 24948
rect 42708 24896 42760 24948
rect 45836 24939 45888 24948
rect 45836 24905 45845 24939
rect 45845 24905 45879 24939
rect 45879 24905 45888 24939
rect 45836 24896 45888 24905
rect 45928 24939 45980 24948
rect 45928 24905 45937 24939
rect 45937 24905 45971 24939
rect 45971 24905 45980 24939
rect 45928 24896 45980 24905
rect 47400 24896 47452 24948
rect 49424 24896 49476 24948
rect 49976 24896 50028 24948
rect 50528 24896 50580 24948
rect 52000 24896 52052 24948
rect 54116 24896 54168 24948
rect 55312 24896 55364 24948
rect 40040 24828 40092 24880
rect 36268 24760 36320 24812
rect 37556 24760 37608 24812
rect 38476 24760 38528 24812
rect 39948 24760 40000 24812
rect 36084 24692 36136 24744
rect 25964 24624 26016 24676
rect 26332 24599 26384 24608
rect 26332 24565 26341 24599
rect 26341 24565 26375 24599
rect 26375 24565 26384 24599
rect 26332 24556 26384 24565
rect 32312 24624 32364 24676
rect 29000 24556 29052 24608
rect 29368 24599 29420 24608
rect 29368 24565 29377 24599
rect 29377 24565 29411 24599
rect 29411 24565 29420 24599
rect 29368 24556 29420 24565
rect 31392 24599 31444 24608
rect 31392 24565 31401 24599
rect 31401 24565 31435 24599
rect 31435 24565 31444 24599
rect 31392 24556 31444 24565
rect 31760 24556 31812 24608
rect 32772 24556 32824 24608
rect 34520 24556 34572 24608
rect 37464 24599 37516 24608
rect 37464 24565 37473 24599
rect 37473 24565 37507 24599
rect 37507 24565 37516 24599
rect 37464 24556 37516 24565
rect 38752 24624 38804 24676
rect 39856 24624 39908 24676
rect 40960 24803 41012 24812
rect 40960 24769 40969 24803
rect 40969 24769 41003 24803
rect 41003 24769 41012 24803
rect 40960 24760 41012 24769
rect 41420 24760 41472 24812
rect 41788 24803 41840 24812
rect 41788 24769 41797 24803
rect 41797 24769 41831 24803
rect 41831 24769 41840 24803
rect 41788 24760 41840 24769
rect 41328 24692 41380 24744
rect 42156 24760 42208 24812
rect 42708 24803 42760 24812
rect 42708 24769 42717 24803
rect 42717 24769 42751 24803
rect 42751 24769 42760 24803
rect 42708 24760 42760 24769
rect 46112 24803 46164 24812
rect 46112 24769 46121 24803
rect 46121 24769 46155 24803
rect 46155 24769 46164 24803
rect 46112 24760 46164 24769
rect 48780 24871 48832 24880
rect 48780 24837 48789 24871
rect 48789 24837 48823 24871
rect 48823 24837 48832 24871
rect 48780 24828 48832 24837
rect 48964 24828 49016 24880
rect 50160 24828 50212 24880
rect 50712 24871 50764 24880
rect 46480 24760 46532 24812
rect 38292 24556 38344 24608
rect 39580 24599 39632 24608
rect 39580 24565 39589 24599
rect 39589 24565 39623 24599
rect 39623 24565 39632 24599
rect 39580 24556 39632 24565
rect 39672 24556 39724 24608
rect 40132 24556 40184 24608
rect 40500 24599 40552 24608
rect 40500 24565 40509 24599
rect 40509 24565 40543 24599
rect 40543 24565 40552 24599
rect 40500 24556 40552 24565
rect 41788 24556 41840 24608
rect 42892 24692 42944 24744
rect 42984 24692 43036 24744
rect 43812 24735 43864 24744
rect 43812 24701 43821 24735
rect 43821 24701 43855 24735
rect 43855 24701 43864 24735
rect 43812 24692 43864 24701
rect 42800 24624 42852 24676
rect 43628 24624 43680 24676
rect 42432 24599 42484 24608
rect 42432 24565 42441 24599
rect 42441 24565 42475 24599
rect 42475 24565 42484 24599
rect 42432 24556 42484 24565
rect 42984 24556 43036 24608
rect 43720 24599 43772 24608
rect 43720 24565 43729 24599
rect 43729 24565 43763 24599
rect 43763 24565 43772 24599
rect 43720 24556 43772 24565
rect 46388 24556 46440 24608
rect 47032 24556 47084 24608
rect 47216 24556 47268 24608
rect 49240 24735 49292 24744
rect 49240 24701 49249 24735
rect 49249 24701 49283 24735
rect 49283 24701 49292 24735
rect 49240 24692 49292 24701
rect 49976 24803 50028 24812
rect 49976 24769 49985 24803
rect 49985 24769 50019 24803
rect 50019 24769 50028 24803
rect 49976 24760 50028 24769
rect 50252 24803 50304 24812
rect 50252 24769 50261 24803
rect 50261 24769 50295 24803
rect 50295 24769 50304 24803
rect 50252 24760 50304 24769
rect 50712 24837 50721 24871
rect 50721 24837 50755 24871
rect 50755 24837 50764 24871
rect 50712 24828 50764 24837
rect 50620 24760 50672 24812
rect 51356 24760 51408 24812
rect 52828 24803 52880 24812
rect 52828 24769 52837 24803
rect 52837 24769 52871 24803
rect 52871 24769 52880 24803
rect 52828 24760 52880 24769
rect 53472 24760 53524 24812
rect 55404 24803 55456 24812
rect 55404 24769 55411 24803
rect 55411 24769 55456 24803
rect 55404 24760 55456 24769
rect 51632 24692 51684 24744
rect 53380 24735 53432 24744
rect 53380 24701 53389 24735
rect 53389 24701 53423 24735
rect 53423 24701 53432 24735
rect 53380 24692 53432 24701
rect 49608 24624 49660 24676
rect 50896 24624 50948 24676
rect 55312 24624 55364 24676
rect 48964 24556 49016 24608
rect 49424 24599 49476 24608
rect 49424 24565 49433 24599
rect 49433 24565 49467 24599
rect 49467 24565 49476 24599
rect 49424 24556 49476 24565
rect 54208 24556 54260 24608
rect 55680 24803 55732 24812
rect 55680 24769 55694 24803
rect 55694 24769 55728 24803
rect 55728 24769 55732 24803
rect 55680 24760 55732 24769
rect 56232 24828 56284 24880
rect 56508 24828 56560 24880
rect 56232 24735 56284 24744
rect 56232 24701 56241 24735
rect 56241 24701 56275 24735
rect 56275 24701 56284 24735
rect 56232 24692 56284 24701
rect 55588 24624 55640 24676
rect 56324 24556 56376 24608
rect 57704 24599 57756 24608
rect 57704 24565 57713 24599
rect 57713 24565 57747 24599
rect 57747 24565 57756 24599
rect 57704 24556 57756 24565
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 20444 24352 20496 24404
rect 22560 24352 22612 24404
rect 22928 24352 22980 24404
rect 23112 24352 23164 24404
rect 25136 24352 25188 24404
rect 26516 24395 26568 24404
rect 26516 24361 26525 24395
rect 26525 24361 26559 24395
rect 26559 24361 26568 24395
rect 26516 24352 26568 24361
rect 27804 24352 27856 24404
rect 31760 24352 31812 24404
rect 31852 24352 31904 24404
rect 32128 24352 32180 24404
rect 32588 24352 32640 24404
rect 33140 24352 33192 24404
rect 34060 24395 34112 24404
rect 34060 24361 34069 24395
rect 34069 24361 34103 24395
rect 34103 24361 34112 24395
rect 34060 24352 34112 24361
rect 34520 24395 34572 24404
rect 34520 24361 34529 24395
rect 34529 24361 34563 24395
rect 34563 24361 34572 24395
rect 34520 24352 34572 24361
rect 35992 24352 36044 24404
rect 36084 24352 36136 24404
rect 21824 24284 21876 24336
rect 21548 24216 21600 24268
rect 22560 24216 22612 24268
rect 18512 24012 18564 24064
rect 19524 24191 19576 24200
rect 19524 24157 19533 24191
rect 19533 24157 19567 24191
rect 19567 24157 19576 24191
rect 19524 24148 19576 24157
rect 19984 24148 20036 24200
rect 22284 24148 22336 24200
rect 22468 24191 22520 24200
rect 22468 24157 22477 24191
rect 22477 24157 22511 24191
rect 22511 24157 22520 24191
rect 22468 24148 22520 24157
rect 23296 24327 23348 24336
rect 23296 24293 23305 24327
rect 23305 24293 23339 24327
rect 23339 24293 23348 24327
rect 23296 24284 23348 24293
rect 25320 24284 25372 24336
rect 26056 24284 26108 24336
rect 23572 24216 23624 24268
rect 26424 24216 26476 24268
rect 23664 24148 23716 24200
rect 25044 24148 25096 24200
rect 25228 24191 25280 24200
rect 25228 24157 25237 24191
rect 25237 24157 25271 24191
rect 25271 24157 25280 24191
rect 25228 24148 25280 24157
rect 25412 24191 25464 24200
rect 25412 24157 25421 24191
rect 25421 24157 25455 24191
rect 25455 24157 25464 24191
rect 25412 24148 25464 24157
rect 25504 24191 25556 24200
rect 25504 24157 25513 24191
rect 25513 24157 25547 24191
rect 25547 24157 25556 24191
rect 25504 24148 25556 24157
rect 22100 24080 22152 24132
rect 22928 24080 22980 24132
rect 25780 24191 25832 24200
rect 25780 24157 25789 24191
rect 25789 24157 25823 24191
rect 25823 24157 25832 24191
rect 25780 24148 25832 24157
rect 25872 24123 25924 24132
rect 25872 24089 25881 24123
rect 25881 24089 25915 24123
rect 25915 24089 25924 24123
rect 25872 24080 25924 24089
rect 26332 24123 26384 24132
rect 26332 24089 26341 24123
rect 26341 24089 26375 24123
rect 26375 24089 26384 24123
rect 26332 24080 26384 24089
rect 20260 24012 20312 24064
rect 21824 24012 21876 24064
rect 22192 24055 22244 24064
rect 22192 24021 22201 24055
rect 22201 24021 22235 24055
rect 22235 24021 22244 24055
rect 22192 24012 22244 24021
rect 24952 24012 25004 24064
rect 25596 24012 25648 24064
rect 25688 24012 25740 24064
rect 27436 24284 27488 24336
rect 28080 24216 28132 24268
rect 28356 24216 28408 24268
rect 26976 24148 27028 24200
rect 28172 24191 28224 24200
rect 28172 24157 28181 24191
rect 28181 24157 28215 24191
rect 28215 24157 28224 24191
rect 28172 24148 28224 24157
rect 29368 24216 29420 24268
rect 28816 24191 28868 24200
rect 28816 24157 28825 24191
rect 28825 24157 28859 24191
rect 28859 24157 28868 24191
rect 28816 24148 28868 24157
rect 29092 24148 29144 24200
rect 31392 24259 31444 24268
rect 31392 24225 31401 24259
rect 31401 24225 31435 24259
rect 31435 24225 31444 24259
rect 31392 24216 31444 24225
rect 33048 24216 33100 24268
rect 27896 24012 27948 24064
rect 30012 24012 30064 24064
rect 30380 24191 30432 24200
rect 30380 24157 30425 24191
rect 30425 24157 30432 24191
rect 30380 24148 30432 24157
rect 30932 24148 30984 24200
rect 31024 24191 31076 24200
rect 31024 24157 31033 24191
rect 31033 24157 31067 24191
rect 31067 24157 31076 24191
rect 31024 24148 31076 24157
rect 33140 24191 33192 24200
rect 33140 24157 33149 24191
rect 33149 24157 33183 24191
rect 33183 24157 33192 24191
rect 33140 24148 33192 24157
rect 32220 24080 32272 24132
rect 32680 24080 32732 24132
rect 33048 24080 33100 24132
rect 33968 24148 34020 24200
rect 34980 24284 35032 24336
rect 35256 24284 35308 24336
rect 39948 24352 40000 24404
rect 42708 24352 42760 24404
rect 47400 24352 47452 24404
rect 34796 24216 34848 24268
rect 35348 24216 35400 24268
rect 35900 24259 35952 24268
rect 35900 24225 35909 24259
rect 35909 24225 35943 24259
rect 35943 24225 35952 24259
rect 35900 24216 35952 24225
rect 36360 24327 36412 24336
rect 36360 24293 36369 24327
rect 36369 24293 36403 24327
rect 36403 24293 36412 24327
rect 36360 24284 36412 24293
rect 38292 24284 38344 24336
rect 39764 24284 39816 24336
rect 41512 24284 41564 24336
rect 42524 24284 42576 24336
rect 48688 24352 48740 24404
rect 48780 24352 48832 24404
rect 49516 24352 49568 24404
rect 49700 24352 49752 24404
rect 50528 24352 50580 24404
rect 50988 24395 51040 24404
rect 50988 24361 50997 24395
rect 50997 24361 51031 24395
rect 51031 24361 51040 24395
rect 50988 24352 51040 24361
rect 34520 24191 34572 24200
rect 34520 24157 34529 24191
rect 34529 24157 34563 24191
rect 34563 24157 34572 24191
rect 34520 24148 34572 24157
rect 35624 24148 35676 24200
rect 36820 24216 36872 24268
rect 39672 24216 39724 24268
rect 30656 24055 30708 24064
rect 30656 24021 30665 24055
rect 30665 24021 30699 24055
rect 30699 24021 30708 24055
rect 30656 24012 30708 24021
rect 30840 24055 30892 24064
rect 30840 24021 30849 24055
rect 30849 24021 30883 24055
rect 30883 24021 30892 24055
rect 30840 24012 30892 24021
rect 31484 24012 31536 24064
rect 35716 24080 35768 24132
rect 35900 24080 35952 24132
rect 36084 24157 36093 24166
rect 36093 24157 36127 24166
rect 36127 24157 36136 24166
rect 36084 24114 36136 24157
rect 36544 24148 36596 24200
rect 36728 24191 36780 24200
rect 36728 24157 36737 24191
rect 36737 24157 36771 24191
rect 36771 24157 36780 24191
rect 36728 24148 36780 24157
rect 36912 24191 36964 24200
rect 36912 24157 36921 24191
rect 36921 24157 36955 24191
rect 36955 24157 36964 24191
rect 36912 24148 36964 24157
rect 37096 24191 37148 24200
rect 37096 24157 37105 24191
rect 37105 24157 37139 24191
rect 37139 24157 37148 24191
rect 37096 24148 37148 24157
rect 39580 24148 39632 24200
rect 39948 24148 40000 24200
rect 45652 24216 45704 24268
rect 41328 24148 41380 24200
rect 42156 24148 42208 24200
rect 33968 24055 34020 24064
rect 33968 24021 33977 24055
rect 33977 24021 34011 24055
rect 34011 24021 34020 24055
rect 33968 24012 34020 24021
rect 37004 24080 37056 24132
rect 39488 24080 39540 24132
rect 40040 24080 40092 24132
rect 40776 24123 40828 24132
rect 40776 24089 40785 24123
rect 40785 24089 40819 24123
rect 40819 24089 40828 24123
rect 40776 24080 40828 24089
rect 41420 24080 41472 24132
rect 43720 24148 43772 24200
rect 46848 24216 46900 24268
rect 48412 24216 48464 24268
rect 48688 24216 48740 24268
rect 48964 24216 49016 24268
rect 50712 24284 50764 24336
rect 54392 24352 54444 24404
rect 56232 24352 56284 24404
rect 53840 24284 53892 24336
rect 49884 24216 49936 24268
rect 52368 24216 52420 24268
rect 42432 24123 42484 24132
rect 42432 24089 42441 24123
rect 42441 24089 42475 24123
rect 42475 24089 42484 24123
rect 42432 24080 42484 24089
rect 42984 24123 43036 24132
rect 42984 24089 42993 24123
rect 42993 24089 43027 24123
rect 43027 24089 43036 24123
rect 42984 24080 43036 24089
rect 43260 24123 43312 24132
rect 43260 24089 43269 24123
rect 43269 24089 43303 24123
rect 43303 24089 43312 24123
rect 43260 24080 43312 24089
rect 45284 24080 45336 24132
rect 46388 24123 46440 24132
rect 46388 24089 46397 24123
rect 46397 24089 46431 24123
rect 46431 24089 46440 24123
rect 46388 24080 46440 24089
rect 46940 24080 46992 24132
rect 47308 24080 47360 24132
rect 47584 24080 47636 24132
rect 47768 24123 47820 24132
rect 47768 24089 47777 24123
rect 47777 24089 47811 24123
rect 47811 24089 47820 24123
rect 47768 24080 47820 24089
rect 38752 24055 38804 24064
rect 38752 24021 38761 24055
rect 38761 24021 38795 24055
rect 38795 24021 38804 24055
rect 38752 24012 38804 24021
rect 39120 24012 39172 24064
rect 39948 24012 40000 24064
rect 43168 24012 43220 24064
rect 44824 24055 44876 24064
rect 44824 24021 44833 24055
rect 44833 24021 44867 24055
rect 44867 24021 44876 24055
rect 44824 24012 44876 24021
rect 47124 24012 47176 24064
rect 49424 24148 49476 24200
rect 54116 24259 54168 24268
rect 54116 24225 54125 24259
rect 54125 24225 54159 24259
rect 54159 24225 54168 24259
rect 54116 24216 54168 24225
rect 55220 24216 55272 24268
rect 56416 24216 56468 24268
rect 57704 24284 57756 24336
rect 50712 24191 50764 24200
rect 50712 24157 50721 24191
rect 50721 24157 50755 24191
rect 50755 24157 50764 24191
rect 50712 24148 50764 24157
rect 50804 24191 50856 24200
rect 50804 24157 50813 24191
rect 50813 24157 50847 24191
rect 50847 24157 50856 24191
rect 50804 24148 50856 24157
rect 52184 24191 52236 24200
rect 52184 24157 52193 24191
rect 52193 24157 52227 24191
rect 52227 24157 52236 24191
rect 52184 24148 52236 24157
rect 53564 24191 53616 24200
rect 53564 24157 53573 24191
rect 53573 24157 53607 24191
rect 53607 24157 53616 24191
rect 53564 24148 53616 24157
rect 49976 24080 50028 24132
rect 48136 24055 48188 24064
rect 48136 24021 48145 24055
rect 48145 24021 48179 24055
rect 48179 24021 48188 24055
rect 48136 24012 48188 24021
rect 48320 24012 48372 24064
rect 48596 24012 48648 24064
rect 50712 24012 50764 24064
rect 53380 24123 53432 24132
rect 53380 24089 53389 24123
rect 53389 24089 53423 24123
rect 53423 24089 53432 24123
rect 53380 24080 53432 24089
rect 53840 24148 53892 24200
rect 54024 24191 54076 24200
rect 54024 24157 54033 24191
rect 54033 24157 54067 24191
rect 54067 24157 54076 24191
rect 54024 24148 54076 24157
rect 54392 24191 54444 24200
rect 54392 24157 54401 24191
rect 54401 24157 54435 24191
rect 54435 24157 54444 24191
rect 54392 24148 54444 24157
rect 54852 24148 54904 24200
rect 56324 24191 56376 24200
rect 56324 24157 56333 24191
rect 56333 24157 56367 24191
rect 56367 24157 56376 24191
rect 56324 24148 56376 24157
rect 57428 24191 57480 24200
rect 57428 24157 57437 24191
rect 57437 24157 57471 24191
rect 57471 24157 57480 24191
rect 57428 24148 57480 24157
rect 54300 24012 54352 24064
rect 54760 24012 54812 24064
rect 56508 24012 56560 24064
rect 58256 24012 58308 24064
rect 4874 23910 4926 23962
rect 4938 23910 4990 23962
rect 5002 23910 5054 23962
rect 5066 23910 5118 23962
rect 5130 23910 5182 23962
rect 35594 23910 35646 23962
rect 35658 23910 35710 23962
rect 35722 23910 35774 23962
rect 35786 23910 35838 23962
rect 35850 23910 35902 23962
rect 19524 23808 19576 23860
rect 18512 23783 18564 23792
rect 18512 23749 18521 23783
rect 18521 23749 18555 23783
rect 18555 23749 18564 23783
rect 18512 23740 18564 23749
rect 20996 23808 21048 23860
rect 20812 23740 20864 23792
rect 19524 23672 19576 23724
rect 19800 23672 19852 23724
rect 20628 23715 20680 23724
rect 20628 23681 20637 23715
rect 20637 23681 20671 23715
rect 20671 23681 20680 23715
rect 22928 23808 22980 23860
rect 23112 23808 23164 23860
rect 25044 23851 25096 23860
rect 25044 23817 25053 23851
rect 25053 23817 25087 23851
rect 25087 23817 25096 23851
rect 25044 23808 25096 23817
rect 25228 23808 25280 23860
rect 22100 23740 22152 23792
rect 22836 23783 22888 23792
rect 22836 23749 22845 23783
rect 22845 23749 22879 23783
rect 22879 23749 22888 23783
rect 22836 23740 22888 23749
rect 25596 23740 25648 23792
rect 20628 23672 20680 23681
rect 19248 23604 19300 23656
rect 22008 23715 22060 23724
rect 22008 23681 22017 23715
rect 22017 23681 22051 23715
rect 22051 23681 22060 23715
rect 22008 23672 22060 23681
rect 23572 23672 23624 23724
rect 23756 23715 23808 23724
rect 23756 23681 23765 23715
rect 23765 23681 23799 23715
rect 23799 23681 23808 23715
rect 23756 23672 23808 23681
rect 23848 23715 23900 23724
rect 23848 23681 23857 23715
rect 23857 23681 23891 23715
rect 23891 23681 23900 23715
rect 23848 23672 23900 23681
rect 24032 23715 24084 23724
rect 24032 23681 24041 23715
rect 24041 23681 24075 23715
rect 24075 23681 24084 23715
rect 24032 23672 24084 23681
rect 22284 23604 22336 23656
rect 19248 23468 19300 23520
rect 19984 23511 20036 23520
rect 19984 23477 19993 23511
rect 19993 23477 20027 23511
rect 20027 23477 20036 23511
rect 25320 23672 25372 23724
rect 25688 23715 25740 23724
rect 25688 23681 25697 23715
rect 25697 23681 25731 23715
rect 25731 23681 25740 23715
rect 25688 23672 25740 23681
rect 26608 23808 26660 23860
rect 31668 23808 31720 23860
rect 31760 23808 31812 23860
rect 32220 23808 32272 23860
rect 33140 23808 33192 23860
rect 26424 23783 26476 23792
rect 26424 23749 26433 23783
rect 26433 23749 26467 23783
rect 26467 23749 26476 23783
rect 26424 23740 26476 23749
rect 27068 23783 27120 23792
rect 27068 23749 27077 23783
rect 27077 23749 27111 23783
rect 27111 23749 27120 23783
rect 27068 23740 27120 23749
rect 19984 23468 20036 23477
rect 25320 23468 25372 23520
rect 26700 23715 26752 23724
rect 26700 23681 26709 23715
rect 26709 23681 26743 23715
rect 26743 23681 26752 23715
rect 26700 23672 26752 23681
rect 27436 23672 27488 23724
rect 27712 23715 27764 23724
rect 27712 23681 27721 23715
rect 27721 23681 27755 23715
rect 27755 23681 27764 23715
rect 27712 23672 27764 23681
rect 27804 23715 27856 23724
rect 27804 23681 27813 23715
rect 27813 23681 27847 23715
rect 27847 23681 27856 23715
rect 27804 23672 27856 23681
rect 28080 23740 28132 23792
rect 28264 23672 28316 23724
rect 27988 23604 28040 23656
rect 28448 23715 28500 23724
rect 28448 23681 28457 23715
rect 28457 23681 28491 23715
rect 28491 23681 28500 23715
rect 28448 23672 28500 23681
rect 32588 23740 32640 23792
rect 32956 23740 33008 23792
rect 33692 23740 33744 23792
rect 32128 23715 32180 23724
rect 32128 23681 32137 23715
rect 32137 23681 32171 23715
rect 32171 23681 32180 23715
rect 32128 23672 32180 23681
rect 32220 23672 32272 23724
rect 33140 23672 33192 23724
rect 33416 23672 33468 23724
rect 34336 23740 34388 23792
rect 34980 23851 35032 23860
rect 34980 23817 34989 23851
rect 34989 23817 35023 23851
rect 35023 23817 35032 23851
rect 34980 23808 35032 23817
rect 35440 23808 35492 23860
rect 37924 23808 37976 23860
rect 38016 23808 38068 23860
rect 25964 23468 26016 23520
rect 28356 23536 28408 23588
rect 28908 23579 28960 23588
rect 28908 23545 28917 23579
rect 28917 23545 28951 23579
rect 28951 23545 28960 23579
rect 28908 23536 28960 23545
rect 30012 23536 30064 23588
rect 34888 23672 34940 23724
rect 35164 23715 35216 23724
rect 35164 23681 35168 23715
rect 35168 23681 35202 23715
rect 35202 23681 35216 23715
rect 35164 23672 35216 23681
rect 35256 23715 35308 23724
rect 35256 23681 35265 23715
rect 35265 23681 35299 23715
rect 35299 23681 35308 23715
rect 35256 23672 35308 23681
rect 35440 23672 35492 23724
rect 36636 23783 36688 23792
rect 36636 23749 36645 23783
rect 36645 23749 36679 23783
rect 36679 23749 36688 23783
rect 36636 23740 36688 23749
rect 36820 23783 36872 23792
rect 36820 23749 36829 23783
rect 36829 23749 36863 23783
rect 36863 23749 36872 23783
rect 36820 23740 36872 23749
rect 34796 23604 34848 23656
rect 38108 23715 38160 23724
rect 38108 23681 38117 23715
rect 38117 23681 38151 23715
rect 38151 23681 38160 23715
rect 38108 23672 38160 23681
rect 38384 23808 38436 23860
rect 39856 23808 39908 23860
rect 40040 23808 40092 23860
rect 38660 23740 38712 23792
rect 38292 23672 38344 23724
rect 39672 23740 39724 23792
rect 39764 23783 39816 23792
rect 39764 23749 39773 23783
rect 39773 23749 39807 23783
rect 39807 23749 39816 23783
rect 39764 23740 39816 23749
rect 40500 23783 40552 23792
rect 40500 23749 40509 23783
rect 40509 23749 40543 23783
rect 40543 23749 40552 23783
rect 40500 23740 40552 23749
rect 42524 23740 42576 23792
rect 42892 23740 42944 23792
rect 43168 23783 43220 23792
rect 43168 23749 43177 23783
rect 43177 23749 43211 23783
rect 43211 23749 43220 23783
rect 43168 23740 43220 23749
rect 39212 23672 39264 23724
rect 42708 23715 42760 23724
rect 42708 23681 42717 23715
rect 42717 23681 42751 23715
rect 42751 23681 42760 23715
rect 42708 23672 42760 23681
rect 42800 23672 42852 23724
rect 45284 23851 45336 23860
rect 45284 23817 45293 23851
rect 45293 23817 45327 23851
rect 45327 23817 45336 23851
rect 45284 23808 45336 23817
rect 46112 23808 46164 23860
rect 47860 23808 47912 23860
rect 44824 23740 44876 23792
rect 45376 23740 45428 23792
rect 46664 23783 46716 23792
rect 46664 23749 46673 23783
rect 46673 23749 46707 23783
rect 46707 23749 46716 23783
rect 48780 23851 48832 23860
rect 48780 23817 48789 23851
rect 48789 23817 48823 23851
rect 48823 23817 48832 23851
rect 48780 23808 48832 23817
rect 49148 23808 49200 23860
rect 52184 23851 52236 23860
rect 46664 23740 46716 23749
rect 45192 23672 45244 23724
rect 46756 23715 46808 23724
rect 46756 23681 46765 23715
rect 46765 23681 46799 23715
rect 46799 23681 46808 23715
rect 46756 23672 46808 23681
rect 46940 23715 46992 23724
rect 46940 23681 46948 23715
rect 46948 23681 46982 23715
rect 46982 23681 46992 23715
rect 46940 23672 46992 23681
rect 47032 23715 47084 23724
rect 47032 23681 47041 23715
rect 47041 23681 47075 23715
rect 47075 23681 47084 23715
rect 47032 23672 47084 23681
rect 47676 23672 47728 23724
rect 47768 23715 47820 23724
rect 47768 23681 47777 23715
rect 47777 23681 47811 23715
rect 47811 23681 47820 23715
rect 47768 23672 47820 23681
rect 47860 23715 47912 23724
rect 47860 23681 47869 23715
rect 47869 23681 47903 23715
rect 47903 23681 47912 23715
rect 47860 23672 47912 23681
rect 47952 23715 48004 23724
rect 47952 23681 47961 23715
rect 47961 23681 47995 23715
rect 47995 23681 48004 23715
rect 47952 23672 48004 23681
rect 49976 23783 50028 23792
rect 49976 23749 49985 23783
rect 49985 23749 50019 23783
rect 50019 23749 50028 23783
rect 49976 23740 50028 23749
rect 52184 23817 52193 23851
rect 52193 23817 52227 23851
rect 52227 23817 52236 23851
rect 52184 23808 52236 23817
rect 53380 23808 53432 23860
rect 54208 23808 54260 23860
rect 54668 23808 54720 23860
rect 55312 23808 55364 23860
rect 50712 23783 50764 23792
rect 50712 23749 50721 23783
rect 50721 23749 50755 23783
rect 50755 23749 50764 23783
rect 50712 23740 50764 23749
rect 51448 23740 51500 23792
rect 35808 23604 35860 23656
rect 36176 23604 36228 23656
rect 36912 23604 36964 23656
rect 28448 23468 28500 23520
rect 28632 23468 28684 23520
rect 28816 23468 28868 23520
rect 29000 23511 29052 23520
rect 29000 23477 29009 23511
rect 29009 23477 29043 23511
rect 29043 23477 29052 23511
rect 29000 23468 29052 23477
rect 32220 23468 32272 23520
rect 32496 23468 32548 23520
rect 32680 23511 32732 23520
rect 32680 23477 32689 23511
rect 32689 23477 32723 23511
rect 32723 23477 32732 23511
rect 32680 23468 32732 23477
rect 33600 23511 33652 23520
rect 33600 23477 33609 23511
rect 33609 23477 33643 23511
rect 33643 23477 33652 23511
rect 33600 23468 33652 23477
rect 37924 23536 37976 23588
rect 40132 23536 40184 23588
rect 41512 23604 41564 23656
rect 43260 23647 43312 23656
rect 43260 23613 43269 23647
rect 43269 23613 43303 23647
rect 43303 23613 43312 23647
rect 43260 23604 43312 23613
rect 34888 23468 34940 23520
rect 36544 23468 36596 23520
rect 38568 23468 38620 23520
rect 38936 23468 38988 23520
rect 40224 23468 40276 23520
rect 43812 23536 43864 23588
rect 44456 23468 44508 23520
rect 45652 23536 45704 23588
rect 47492 23604 47544 23656
rect 48136 23604 48188 23656
rect 48596 23715 48648 23724
rect 48596 23681 48605 23715
rect 48605 23681 48639 23715
rect 48639 23681 48648 23715
rect 48596 23672 48648 23681
rect 49700 23715 49752 23724
rect 49700 23681 49709 23715
rect 49709 23681 49743 23715
rect 49743 23681 49752 23715
rect 49700 23672 49752 23681
rect 49884 23715 49936 23724
rect 49884 23681 49891 23715
rect 49891 23681 49936 23715
rect 49884 23672 49936 23681
rect 48964 23647 49016 23656
rect 48964 23613 48973 23647
rect 48973 23613 49007 23647
rect 49007 23613 49016 23647
rect 48964 23604 49016 23613
rect 45100 23511 45152 23520
rect 45100 23477 45109 23511
rect 45109 23477 45143 23511
rect 45143 23477 45152 23511
rect 45100 23468 45152 23477
rect 47124 23468 47176 23520
rect 48136 23511 48188 23520
rect 48136 23477 48145 23511
rect 48145 23477 48179 23511
rect 48179 23477 48188 23511
rect 48136 23468 48188 23477
rect 48320 23536 48372 23588
rect 53288 23740 53340 23792
rect 54760 23740 54812 23792
rect 50344 23579 50396 23588
rect 50344 23545 50353 23579
rect 50353 23545 50387 23579
rect 50387 23545 50396 23579
rect 50344 23536 50396 23545
rect 49148 23468 49200 23520
rect 49240 23468 49292 23520
rect 52644 23604 52696 23656
rect 53564 23672 53616 23724
rect 58256 23715 58308 23724
rect 58256 23681 58265 23715
rect 58265 23681 58299 23715
rect 58299 23681 58308 23715
rect 58256 23672 58308 23681
rect 53932 23604 53984 23656
rect 54300 23647 54352 23656
rect 54300 23613 54309 23647
rect 54309 23613 54343 23647
rect 54343 23613 54352 23647
rect 54300 23604 54352 23613
rect 56692 23647 56744 23656
rect 56692 23613 56701 23647
rect 56701 23613 56735 23647
rect 56735 23613 56744 23647
rect 56692 23604 56744 23613
rect 57428 23604 57480 23656
rect 53748 23468 53800 23520
rect 54024 23468 54076 23520
rect 55404 23468 55456 23520
rect 55956 23468 56008 23520
rect 58440 23511 58492 23520
rect 58440 23477 58449 23511
rect 58449 23477 58483 23511
rect 58483 23477 58492 23511
rect 58440 23468 58492 23477
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 20996 23307 21048 23316
rect 20996 23273 21005 23307
rect 21005 23273 21039 23307
rect 21039 23273 21048 23307
rect 20996 23264 21048 23273
rect 22192 23264 22244 23316
rect 22468 23264 22520 23316
rect 23664 23264 23716 23316
rect 19248 23171 19300 23180
rect 19248 23137 19257 23171
rect 19257 23137 19291 23171
rect 19291 23137 19300 23171
rect 19248 23128 19300 23137
rect 21548 23171 21600 23180
rect 21548 23137 21557 23171
rect 21557 23137 21591 23171
rect 21591 23137 21600 23171
rect 21548 23128 21600 23137
rect 17960 23060 18012 23112
rect 22100 23171 22152 23180
rect 22100 23137 22109 23171
rect 22109 23137 22143 23171
rect 22143 23137 22152 23171
rect 22100 23128 22152 23137
rect 22376 23171 22428 23180
rect 22376 23137 22385 23171
rect 22385 23137 22419 23171
rect 22419 23137 22428 23171
rect 22376 23128 22428 23137
rect 18604 22992 18656 23044
rect 19616 22992 19668 23044
rect 19892 22924 19944 22976
rect 21824 23103 21876 23112
rect 21824 23069 21833 23103
rect 21833 23069 21867 23103
rect 21867 23069 21876 23103
rect 21824 23060 21876 23069
rect 28816 23264 28868 23316
rect 30380 23264 30432 23316
rect 34796 23264 34848 23316
rect 26700 23196 26752 23248
rect 28816 23128 28868 23180
rect 31024 23128 31076 23180
rect 32864 23171 32916 23180
rect 32864 23137 32873 23171
rect 32873 23137 32907 23171
rect 32907 23137 32916 23171
rect 32864 23128 32916 23137
rect 22192 22924 22244 22976
rect 22836 22992 22888 23044
rect 24860 22992 24912 23044
rect 23664 22924 23716 22976
rect 24032 22924 24084 22976
rect 26056 22924 26108 22976
rect 26332 22967 26384 22976
rect 26332 22933 26341 22967
rect 26341 22933 26375 22967
rect 26375 22933 26384 22967
rect 26332 22924 26384 22933
rect 27528 23103 27580 23112
rect 27528 23069 27537 23103
rect 27537 23069 27571 23103
rect 27571 23069 27580 23103
rect 27528 23060 27580 23069
rect 32588 23103 32640 23112
rect 32588 23069 32597 23103
rect 32597 23069 32631 23103
rect 32631 23069 32640 23103
rect 32588 23060 32640 23069
rect 32680 23103 32732 23112
rect 32680 23069 32689 23103
rect 32689 23069 32723 23103
rect 32723 23069 32732 23103
rect 32680 23060 32732 23069
rect 28080 22992 28132 23044
rect 28448 22992 28500 23044
rect 31576 22992 31628 23044
rect 33048 23060 33100 23112
rect 33692 23128 33744 23180
rect 35348 23128 35400 23180
rect 37464 23128 37516 23180
rect 36268 23060 36320 23112
rect 36452 23060 36504 23112
rect 36636 23060 36688 23112
rect 39212 23307 39264 23316
rect 39212 23273 39221 23307
rect 39221 23273 39255 23307
rect 39255 23273 39264 23307
rect 39212 23264 39264 23273
rect 39580 23264 39632 23316
rect 40132 23307 40184 23316
rect 40132 23273 40141 23307
rect 40141 23273 40175 23307
rect 40175 23273 40184 23307
rect 40132 23264 40184 23273
rect 40592 23264 40644 23316
rect 43444 23264 43496 23316
rect 44180 23264 44232 23316
rect 45468 23264 45520 23316
rect 45836 23264 45888 23316
rect 46664 23307 46716 23316
rect 46664 23273 46673 23307
rect 46673 23273 46707 23307
rect 46707 23273 46716 23307
rect 46664 23264 46716 23273
rect 47768 23264 47820 23316
rect 48504 23264 48556 23316
rect 38936 23196 38988 23248
rect 38292 23171 38344 23180
rect 38292 23137 38301 23171
rect 38301 23137 38335 23171
rect 38335 23137 38344 23171
rect 38292 23128 38344 23137
rect 39120 23060 39172 23112
rect 35624 22992 35676 23044
rect 39396 23060 39448 23112
rect 41604 23196 41656 23248
rect 46020 23196 46072 23248
rect 39764 23128 39816 23180
rect 40132 23128 40184 23180
rect 41696 23128 41748 23180
rect 39948 23103 40000 23112
rect 39948 23069 39957 23103
rect 39957 23069 39991 23103
rect 39991 23069 40000 23103
rect 39948 23060 40000 23069
rect 41420 23103 41472 23112
rect 41420 23069 41429 23103
rect 41429 23069 41463 23103
rect 41463 23069 41472 23103
rect 41420 23060 41472 23069
rect 41604 23103 41656 23112
rect 41604 23069 41613 23103
rect 41613 23069 41647 23103
rect 41647 23069 41656 23103
rect 41604 23060 41656 23069
rect 42432 23128 42484 23180
rect 47492 23128 47544 23180
rect 48412 23171 48464 23180
rect 48412 23137 48421 23171
rect 48421 23137 48455 23171
rect 48455 23137 48464 23171
rect 49240 23264 49292 23316
rect 49700 23264 49752 23316
rect 49884 23264 49936 23316
rect 50804 23264 50856 23316
rect 53840 23264 53892 23316
rect 48412 23128 48464 23137
rect 27988 22924 28040 22976
rect 32312 22924 32364 22976
rect 33968 22924 34020 22976
rect 36820 22924 36872 22976
rect 38660 22967 38712 22976
rect 38660 22933 38669 22967
rect 38669 22933 38703 22967
rect 38703 22933 38712 22967
rect 38660 22924 38712 22933
rect 39580 22924 39632 22976
rect 39764 22924 39816 22976
rect 42800 23060 42852 23112
rect 43444 23103 43496 23112
rect 43444 23069 43453 23103
rect 43453 23069 43487 23103
rect 43487 23069 43496 23103
rect 43444 23060 43496 23069
rect 45192 23103 45244 23112
rect 45192 23069 45196 23103
rect 45196 23069 45230 23103
rect 45230 23069 45244 23103
rect 42156 23035 42208 23044
rect 42156 23001 42165 23035
rect 42165 23001 42199 23035
rect 42199 23001 42208 23035
rect 42156 22992 42208 23001
rect 42340 22992 42392 23044
rect 45192 23060 45244 23069
rect 42248 22924 42300 22976
rect 43904 22967 43956 22976
rect 43904 22933 43913 22967
rect 43913 22933 43947 22967
rect 43947 22933 43956 22967
rect 43904 22924 43956 22933
rect 44364 22967 44416 22976
rect 44364 22933 44373 22967
rect 44373 22933 44407 22967
rect 44407 22933 44416 22967
rect 44364 22924 44416 22933
rect 45284 23035 45336 23044
rect 45284 23001 45293 23035
rect 45293 23001 45327 23035
rect 45327 23001 45336 23035
rect 45284 22992 45336 23001
rect 45652 23103 45704 23112
rect 45652 23069 45661 23103
rect 45661 23069 45695 23103
rect 45695 23069 45704 23103
rect 45652 23060 45704 23069
rect 46296 23103 46348 23112
rect 46296 23069 46305 23103
rect 46305 23069 46339 23103
rect 46339 23069 46348 23103
rect 46296 23060 46348 23069
rect 49884 23060 49936 23112
rect 52368 23196 52420 23248
rect 46664 22992 46716 23044
rect 47584 22992 47636 23044
rect 48872 22992 48924 23044
rect 48964 23035 49016 23044
rect 48964 23001 48973 23035
rect 48973 23001 49007 23035
rect 49007 23001 49016 23035
rect 48964 22992 49016 23001
rect 45560 22924 45612 22976
rect 46756 22924 46808 22976
rect 47216 22924 47268 22976
rect 50712 23103 50764 23112
rect 50712 23069 50721 23103
rect 50721 23069 50755 23103
rect 50755 23069 50764 23103
rect 50712 23060 50764 23069
rect 50804 22992 50856 23044
rect 52920 22992 52972 23044
rect 53380 23035 53432 23044
rect 53380 23001 53389 23035
rect 53389 23001 53423 23035
rect 53423 23001 53432 23035
rect 53380 22992 53432 23001
rect 53932 23060 53984 23112
rect 57428 23307 57480 23316
rect 57428 23273 57437 23307
rect 57437 23273 57471 23307
rect 57471 23273 57480 23307
rect 57428 23264 57480 23273
rect 55956 23171 56008 23180
rect 55956 23137 55965 23171
rect 55965 23137 55999 23171
rect 55999 23137 56008 23171
rect 55956 23128 56008 23137
rect 55588 23060 55640 23112
rect 51908 22967 51960 22976
rect 51908 22933 51917 22967
rect 51917 22933 51951 22967
rect 51951 22933 51960 22967
rect 51908 22924 51960 22933
rect 52460 22924 52512 22976
rect 53656 22924 53708 22976
rect 56600 22924 56652 22976
rect 4874 22822 4926 22874
rect 4938 22822 4990 22874
rect 5002 22822 5054 22874
rect 5066 22822 5118 22874
rect 5130 22822 5182 22874
rect 35594 22822 35646 22874
rect 35658 22822 35710 22874
rect 35722 22822 35774 22874
rect 35786 22822 35838 22874
rect 35850 22822 35902 22874
rect 17960 22652 18012 22704
rect 19248 22652 19300 22704
rect 18328 22627 18380 22636
rect 18328 22593 18337 22627
rect 18337 22593 18371 22627
rect 18371 22593 18380 22627
rect 22008 22720 22060 22772
rect 19800 22627 19852 22636
rect 18328 22584 18380 22593
rect 19800 22593 19804 22627
rect 19804 22593 19838 22627
rect 19838 22593 19852 22627
rect 19800 22584 19852 22593
rect 19892 22627 19944 22636
rect 19892 22593 19901 22627
rect 19901 22593 19935 22627
rect 19935 22593 19944 22627
rect 19892 22584 19944 22593
rect 19984 22627 20036 22636
rect 19984 22593 19993 22627
rect 19993 22593 20027 22627
rect 20027 22593 20036 22627
rect 19984 22584 20036 22593
rect 20076 22627 20128 22636
rect 22100 22652 22152 22704
rect 22836 22720 22888 22772
rect 23664 22720 23716 22772
rect 22560 22652 22612 22704
rect 20076 22593 20121 22627
rect 20121 22593 20128 22627
rect 20076 22584 20128 22593
rect 20352 22516 20404 22568
rect 23756 22584 23808 22636
rect 25596 22584 25648 22636
rect 27436 22720 27488 22772
rect 28080 22763 28132 22772
rect 28080 22729 28089 22763
rect 28089 22729 28123 22763
rect 28123 22729 28132 22763
rect 28080 22720 28132 22729
rect 34612 22720 34664 22772
rect 35992 22720 36044 22772
rect 26332 22652 26384 22704
rect 28540 22652 28592 22704
rect 32128 22652 32180 22704
rect 34796 22652 34848 22704
rect 22192 22516 22244 22568
rect 26976 22584 27028 22636
rect 28264 22627 28316 22636
rect 28264 22593 28273 22627
rect 28273 22593 28307 22627
rect 28307 22593 28316 22627
rect 28264 22584 28316 22593
rect 28356 22627 28408 22636
rect 28356 22593 28365 22627
rect 28365 22593 28399 22627
rect 28399 22593 28408 22627
rect 28356 22584 28408 22593
rect 28448 22584 28500 22636
rect 28816 22584 28868 22636
rect 19616 22423 19668 22432
rect 19616 22389 19625 22423
rect 19625 22389 19659 22423
rect 19659 22389 19668 22423
rect 19616 22380 19668 22389
rect 20444 22423 20496 22432
rect 20444 22389 20453 22423
rect 20453 22389 20487 22423
rect 20487 22389 20496 22423
rect 20444 22380 20496 22389
rect 21824 22380 21876 22432
rect 31576 22516 31628 22568
rect 32404 22627 32456 22636
rect 32404 22593 32413 22627
rect 32413 22593 32447 22627
rect 32447 22593 32456 22627
rect 32404 22584 32456 22593
rect 32680 22627 32732 22636
rect 32680 22593 32689 22627
rect 32689 22593 32723 22627
rect 32723 22593 32732 22627
rect 32680 22584 32732 22593
rect 34704 22584 34756 22636
rect 33232 22516 33284 22568
rect 25872 22491 25924 22500
rect 25872 22457 25881 22491
rect 25881 22457 25915 22491
rect 25915 22457 25924 22491
rect 25872 22448 25924 22457
rect 26240 22448 26292 22500
rect 30012 22448 30064 22500
rect 32772 22448 32824 22500
rect 34428 22448 34480 22500
rect 35348 22584 35400 22636
rect 35808 22695 35860 22704
rect 35808 22661 35817 22695
rect 35817 22661 35851 22695
rect 35851 22661 35860 22695
rect 35808 22652 35860 22661
rect 35900 22516 35952 22568
rect 36084 22584 36136 22636
rect 36452 22584 36504 22636
rect 37832 22763 37884 22772
rect 37832 22729 37841 22763
rect 37841 22729 37875 22763
rect 37875 22729 37884 22763
rect 37832 22720 37884 22729
rect 38660 22720 38712 22772
rect 39396 22763 39448 22772
rect 39396 22729 39405 22763
rect 39405 22729 39439 22763
rect 39439 22729 39448 22763
rect 39396 22720 39448 22729
rect 36636 22627 36688 22636
rect 36636 22593 36645 22627
rect 36645 22593 36679 22627
rect 36679 22593 36688 22627
rect 36636 22584 36688 22593
rect 37556 22584 37608 22636
rect 38384 22627 38436 22636
rect 38384 22593 38393 22627
rect 38393 22593 38427 22627
rect 38427 22593 38436 22627
rect 38384 22584 38436 22593
rect 39120 22584 39172 22636
rect 36360 22559 36412 22568
rect 36360 22525 36369 22559
rect 36369 22525 36403 22559
rect 36403 22525 36412 22559
rect 36360 22516 36412 22525
rect 36820 22516 36872 22568
rect 42340 22720 42392 22772
rect 42708 22720 42760 22772
rect 39580 22627 39632 22636
rect 39580 22593 39589 22627
rect 39589 22593 39623 22627
rect 39623 22593 39632 22627
rect 39580 22584 39632 22593
rect 39948 22584 40000 22636
rect 43536 22652 43588 22704
rect 44364 22695 44416 22704
rect 44364 22661 44373 22695
rect 44373 22661 44407 22695
rect 44407 22661 44416 22695
rect 44364 22652 44416 22661
rect 48872 22763 48924 22772
rect 48872 22729 48881 22763
rect 48881 22729 48915 22763
rect 48915 22729 48924 22763
rect 48872 22720 48924 22729
rect 49056 22763 49108 22772
rect 49056 22729 49065 22763
rect 49065 22729 49099 22763
rect 49099 22729 49108 22763
rect 49056 22720 49108 22729
rect 49700 22720 49752 22772
rect 53288 22720 53340 22772
rect 53380 22720 53432 22772
rect 48136 22652 48188 22704
rect 41604 22584 41656 22636
rect 42248 22584 42300 22636
rect 42616 22627 42668 22636
rect 42616 22593 42625 22627
rect 42625 22593 42659 22627
rect 42659 22593 42668 22627
rect 42616 22584 42668 22593
rect 41512 22516 41564 22568
rect 42524 22516 42576 22568
rect 42984 22627 43036 22636
rect 42984 22593 42993 22627
rect 42993 22593 43027 22627
rect 43027 22593 43036 22627
rect 42984 22584 43036 22593
rect 46664 22584 46716 22636
rect 53656 22652 53708 22704
rect 55588 22652 55640 22704
rect 43996 22516 44048 22568
rect 26332 22423 26384 22432
rect 26332 22389 26341 22423
rect 26341 22389 26375 22423
rect 26375 22389 26384 22423
rect 26332 22380 26384 22389
rect 32128 22423 32180 22432
rect 32128 22389 32137 22423
rect 32137 22389 32171 22423
rect 32171 22389 32180 22423
rect 32128 22380 32180 22389
rect 32864 22380 32916 22432
rect 33140 22380 33192 22432
rect 33600 22380 33652 22432
rect 35348 22380 35400 22432
rect 37648 22380 37700 22432
rect 37832 22380 37884 22432
rect 39764 22423 39816 22432
rect 39764 22389 39773 22423
rect 39773 22389 39807 22423
rect 39807 22389 39816 22423
rect 39764 22380 39816 22389
rect 41144 22423 41196 22432
rect 41144 22389 41153 22423
rect 41153 22389 41187 22423
rect 41187 22389 41196 22423
rect 41144 22380 41196 22389
rect 47216 22516 47268 22568
rect 47676 22516 47728 22568
rect 49240 22627 49292 22636
rect 49240 22593 49249 22627
rect 49249 22593 49283 22627
rect 49283 22593 49292 22627
rect 49240 22584 49292 22593
rect 51908 22584 51960 22636
rect 53748 22627 53800 22636
rect 53748 22593 53757 22627
rect 53757 22593 53791 22627
rect 53791 22593 53800 22627
rect 53748 22584 53800 22593
rect 56140 22627 56192 22636
rect 56140 22593 56149 22627
rect 56149 22593 56183 22627
rect 56183 22593 56192 22627
rect 56140 22584 56192 22593
rect 58256 22627 58308 22636
rect 58256 22593 58265 22627
rect 58265 22593 58299 22627
rect 58299 22593 58308 22627
rect 58256 22584 58308 22593
rect 55864 22559 55916 22568
rect 55864 22525 55873 22559
rect 55873 22525 55907 22559
rect 55907 22525 55916 22559
rect 55864 22516 55916 22525
rect 42156 22380 42208 22432
rect 42984 22380 43036 22432
rect 46296 22380 46348 22432
rect 48044 22380 48096 22432
rect 50988 22448 51040 22500
rect 58440 22491 58492 22500
rect 58440 22457 58449 22491
rect 58449 22457 58483 22491
rect 58483 22457 58492 22491
rect 58440 22448 58492 22457
rect 48688 22380 48740 22432
rect 48872 22380 48924 22432
rect 53564 22423 53616 22432
rect 53564 22389 53573 22423
rect 53573 22389 53607 22423
rect 53607 22389 53616 22423
rect 53564 22380 53616 22389
rect 54392 22423 54444 22432
rect 54392 22389 54401 22423
rect 54401 22389 54435 22423
rect 54435 22389 54444 22423
rect 54392 22380 54444 22389
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 18604 22219 18656 22228
rect 18604 22185 18613 22219
rect 18613 22185 18647 22219
rect 18647 22185 18656 22219
rect 18604 22176 18656 22185
rect 20444 22176 20496 22228
rect 22744 22176 22796 22228
rect 24860 22176 24912 22228
rect 25596 22219 25648 22228
rect 25596 22185 25605 22219
rect 25605 22185 25639 22219
rect 25639 22185 25648 22219
rect 25596 22176 25648 22185
rect 25872 22176 25924 22228
rect 26332 22176 26384 22228
rect 28172 22176 28224 22228
rect 29000 22176 29052 22228
rect 30288 22176 30340 22228
rect 32680 22176 32732 22228
rect 19616 22040 19668 22092
rect 20996 22040 21048 22092
rect 19892 22015 19944 22024
rect 19892 21981 19901 22015
rect 19901 21981 19935 22015
rect 19935 21981 19944 22015
rect 19892 21972 19944 21981
rect 27988 22108 28040 22160
rect 27528 22040 27580 22092
rect 29092 22040 29144 22092
rect 19340 21904 19392 21956
rect 19432 21836 19484 21888
rect 20536 21904 20588 21956
rect 20904 21904 20956 21956
rect 24216 21904 24268 21956
rect 28540 21972 28592 22024
rect 32128 22040 32180 22092
rect 34428 22176 34480 22228
rect 35624 22219 35676 22228
rect 35624 22185 35633 22219
rect 35633 22185 35667 22219
rect 35667 22185 35676 22219
rect 35624 22176 35676 22185
rect 35716 22176 35768 22228
rect 35992 22176 36044 22228
rect 36268 22176 36320 22228
rect 36452 22176 36504 22228
rect 41144 22176 41196 22228
rect 43536 22176 43588 22228
rect 45560 22176 45612 22228
rect 47860 22176 47912 22228
rect 48320 22176 48372 22228
rect 49700 22219 49752 22228
rect 49700 22185 49709 22219
rect 49709 22185 49743 22219
rect 49743 22185 49752 22219
rect 49700 22176 49752 22185
rect 33140 22151 33192 22160
rect 33140 22117 33149 22151
rect 33149 22117 33183 22151
rect 33183 22117 33192 22151
rect 33140 22108 33192 22117
rect 42248 22108 42300 22160
rect 45284 22108 45336 22160
rect 48044 22108 48096 22160
rect 52920 22108 52972 22160
rect 53656 22108 53708 22160
rect 31208 22015 31260 22024
rect 31208 21981 31217 22015
rect 31217 21981 31251 22015
rect 31251 21981 31260 22015
rect 31208 21972 31260 21981
rect 27436 21904 27488 21956
rect 27988 21947 28040 21956
rect 27988 21913 27997 21947
rect 27997 21913 28031 21947
rect 28031 21913 28040 21947
rect 27988 21904 28040 21913
rect 20076 21879 20128 21888
rect 20076 21845 20085 21879
rect 20085 21845 20119 21879
rect 20119 21845 20128 21879
rect 20352 21879 20404 21888
rect 20076 21836 20128 21845
rect 20352 21845 20361 21879
rect 20361 21845 20395 21879
rect 20395 21845 20404 21879
rect 20352 21836 20404 21845
rect 21548 21836 21600 21888
rect 22284 21836 22336 21888
rect 23296 21836 23348 21888
rect 24032 21836 24084 21888
rect 28724 21836 28776 21888
rect 31024 21836 31076 21888
rect 31668 21836 31720 21888
rect 31944 21904 31996 21956
rect 33600 22015 33652 22024
rect 33600 21981 33609 22015
rect 33609 21981 33643 22015
rect 33643 21981 33652 22015
rect 33600 21972 33652 21981
rect 34612 21972 34664 22024
rect 35348 22015 35400 22024
rect 35348 21981 35357 22015
rect 35357 21981 35391 22015
rect 35391 21981 35400 22015
rect 35348 21972 35400 21981
rect 32220 21836 32272 21888
rect 34704 21904 34756 21956
rect 35072 21879 35124 21888
rect 35072 21845 35081 21879
rect 35081 21845 35115 21879
rect 35115 21845 35124 21879
rect 35072 21836 35124 21845
rect 35164 21879 35216 21888
rect 35164 21845 35173 21879
rect 35173 21845 35207 21879
rect 35207 21845 35216 21879
rect 35164 21836 35216 21845
rect 35348 21836 35400 21888
rect 37464 22040 37516 22092
rect 44180 22040 44232 22092
rect 46848 22040 46900 22092
rect 50252 22083 50304 22092
rect 35716 22015 35768 22024
rect 35716 21981 35725 22015
rect 35725 21981 35759 22015
rect 35759 21981 35768 22015
rect 35716 21972 35768 21981
rect 35808 22015 35860 22024
rect 35808 21981 35817 22015
rect 35817 21981 35851 22015
rect 35851 21981 35860 22015
rect 35808 21972 35860 21981
rect 37648 22015 37700 22024
rect 37648 21981 37657 22015
rect 37657 21981 37691 22015
rect 37691 21981 37700 22015
rect 37648 21972 37700 21981
rect 40408 22015 40460 22024
rect 40408 21981 40417 22015
rect 40417 21981 40451 22015
rect 40451 21981 40460 22015
rect 40408 21972 40460 21981
rect 44456 21972 44508 22024
rect 45192 22015 45244 22024
rect 37280 21904 37332 21956
rect 42708 21904 42760 21956
rect 44824 21904 44876 21956
rect 45192 21981 45201 22015
rect 45201 21981 45235 22015
rect 45235 21981 45244 22015
rect 45192 21972 45244 21981
rect 47216 21972 47268 22024
rect 47952 21972 48004 22024
rect 38476 21836 38528 21888
rect 41604 21836 41656 21888
rect 43904 21836 43956 21888
rect 45284 21836 45336 21888
rect 45560 21904 45612 21956
rect 46480 21904 46532 21956
rect 47860 21904 47912 21956
rect 47308 21836 47360 21888
rect 47768 21836 47820 21888
rect 48320 22015 48372 22024
rect 48320 21981 48329 22015
rect 48329 21981 48363 22015
rect 48363 21981 48372 22015
rect 48320 21972 48372 21981
rect 50252 22049 50261 22083
rect 50261 22049 50295 22083
rect 50295 22049 50304 22083
rect 50252 22040 50304 22049
rect 48688 21972 48740 22024
rect 49056 21972 49108 22024
rect 49332 21972 49384 22024
rect 55680 22040 55732 22092
rect 54484 21972 54536 22024
rect 56140 21972 56192 22024
rect 55404 21947 55456 21956
rect 55404 21913 55413 21947
rect 55413 21913 55447 21947
rect 55447 21913 55456 21947
rect 55404 21904 55456 21913
rect 57520 21904 57572 21956
rect 48504 21836 48556 21888
rect 48872 21879 48924 21888
rect 48872 21845 48881 21879
rect 48881 21845 48915 21879
rect 48915 21845 48924 21879
rect 48872 21836 48924 21845
rect 49056 21836 49108 21888
rect 49792 21836 49844 21888
rect 51356 21836 51408 21888
rect 52092 21836 52144 21888
rect 52644 21879 52696 21888
rect 52644 21845 52653 21879
rect 52653 21845 52687 21879
rect 52687 21845 52696 21879
rect 52644 21836 52696 21845
rect 53380 21879 53432 21888
rect 53380 21845 53389 21879
rect 53389 21845 53423 21879
rect 53423 21845 53432 21879
rect 53380 21836 53432 21845
rect 55312 21836 55364 21888
rect 58256 21879 58308 21888
rect 58256 21845 58265 21879
rect 58265 21845 58299 21879
rect 58299 21845 58308 21879
rect 58256 21836 58308 21845
rect 58440 21836 58492 21888
rect 4874 21734 4926 21786
rect 4938 21734 4990 21786
rect 5002 21734 5054 21786
rect 5066 21734 5118 21786
rect 5130 21734 5182 21786
rect 35594 21734 35646 21786
rect 35658 21734 35710 21786
rect 35722 21734 35774 21786
rect 35786 21734 35838 21786
rect 35850 21734 35902 21786
rect 19984 21632 20036 21684
rect 20168 21675 20220 21684
rect 20168 21641 20177 21675
rect 20177 21641 20211 21675
rect 20211 21641 20220 21675
rect 20168 21632 20220 21641
rect 20444 21632 20496 21684
rect 20904 21675 20956 21684
rect 19432 21428 19484 21480
rect 19708 21539 19760 21548
rect 19708 21505 19717 21539
rect 19717 21505 19751 21539
rect 19751 21505 19760 21539
rect 19708 21496 19760 21505
rect 19984 21539 20036 21548
rect 19984 21505 19992 21539
rect 19992 21505 20026 21539
rect 20026 21505 20036 21539
rect 19984 21496 20036 21505
rect 20260 21496 20312 21548
rect 20444 21539 20496 21548
rect 20444 21505 20453 21539
rect 20453 21505 20487 21539
rect 20487 21505 20496 21539
rect 20444 21496 20496 21505
rect 20904 21641 20913 21675
rect 20913 21641 20947 21675
rect 20947 21641 20956 21675
rect 20904 21632 20956 21641
rect 23572 21632 23624 21684
rect 26056 21675 26108 21684
rect 22376 21496 22428 21548
rect 20260 21360 20312 21412
rect 23664 21428 23716 21480
rect 23848 21496 23900 21548
rect 24400 21564 24452 21616
rect 24124 21539 24176 21548
rect 24124 21505 24133 21539
rect 24133 21505 24167 21539
rect 24167 21505 24176 21539
rect 24124 21496 24176 21505
rect 26056 21641 26065 21675
rect 26065 21641 26099 21675
rect 26099 21641 26108 21675
rect 26056 21632 26108 21641
rect 27988 21632 28040 21684
rect 24584 21564 24636 21616
rect 24860 21539 24912 21548
rect 24860 21505 24869 21539
rect 24869 21505 24903 21539
rect 24903 21505 24912 21539
rect 24860 21496 24912 21505
rect 25872 21428 25924 21480
rect 18788 21292 18840 21344
rect 18972 21292 19024 21344
rect 19340 21292 19392 21344
rect 21548 21292 21600 21344
rect 23848 21292 23900 21344
rect 23940 21292 23992 21344
rect 24584 21292 24636 21344
rect 25596 21292 25648 21344
rect 26608 21539 26660 21548
rect 26608 21505 26617 21539
rect 26617 21505 26651 21539
rect 26651 21505 26660 21539
rect 26608 21496 26660 21505
rect 27528 21564 27580 21616
rect 28632 21564 28684 21616
rect 29276 21564 29328 21616
rect 29920 21539 29972 21548
rect 29920 21505 29929 21539
rect 29929 21505 29963 21539
rect 29963 21505 29972 21539
rect 29920 21496 29972 21505
rect 31024 21675 31076 21684
rect 31024 21641 31033 21675
rect 31033 21641 31067 21675
rect 31067 21641 31076 21675
rect 31024 21632 31076 21641
rect 32312 21632 32364 21684
rect 32496 21632 32548 21684
rect 32864 21632 32916 21684
rect 34520 21632 34572 21684
rect 36728 21632 36780 21684
rect 42892 21632 42944 21684
rect 43996 21632 44048 21684
rect 44640 21632 44692 21684
rect 45560 21632 45612 21684
rect 26240 21360 26292 21412
rect 26332 21292 26384 21344
rect 27712 21428 27764 21480
rect 31576 21539 31628 21548
rect 31576 21505 31585 21539
rect 31585 21505 31619 21539
rect 31619 21505 31628 21539
rect 31576 21496 31628 21505
rect 31208 21428 31260 21480
rect 28540 21292 28592 21344
rect 30012 21360 30064 21412
rect 32220 21496 32272 21548
rect 33600 21564 33652 21616
rect 36176 21564 36228 21616
rect 37280 21564 37332 21616
rect 39304 21564 39356 21616
rect 48688 21632 48740 21684
rect 48872 21632 48924 21684
rect 32772 21539 32824 21548
rect 32772 21505 32781 21539
rect 32781 21505 32815 21539
rect 32815 21505 32824 21539
rect 32772 21496 32824 21505
rect 34060 21539 34112 21548
rect 34060 21505 34069 21539
rect 34069 21505 34103 21539
rect 34103 21505 34112 21539
rect 34060 21496 34112 21505
rect 34152 21539 34204 21548
rect 34152 21505 34162 21539
rect 34162 21505 34196 21539
rect 34196 21505 34204 21539
rect 34152 21496 34204 21505
rect 34428 21539 34480 21548
rect 34428 21505 34437 21539
rect 34437 21505 34471 21539
rect 34471 21505 34480 21539
rect 34428 21496 34480 21505
rect 34520 21539 34572 21548
rect 34520 21505 34534 21539
rect 34534 21505 34568 21539
rect 34568 21505 34572 21539
rect 34520 21496 34572 21505
rect 35164 21539 35216 21548
rect 35164 21505 35173 21539
rect 35173 21505 35207 21539
rect 35207 21505 35216 21539
rect 35164 21496 35216 21505
rect 41512 21496 41564 21548
rect 41880 21539 41932 21548
rect 41880 21505 41889 21539
rect 41889 21505 41923 21539
rect 41923 21505 41932 21539
rect 41880 21496 41932 21505
rect 35440 21428 35492 21480
rect 35900 21428 35952 21480
rect 36084 21428 36136 21480
rect 42984 21496 43036 21548
rect 47952 21564 48004 21616
rect 50804 21632 50856 21684
rect 52000 21632 52052 21684
rect 46848 21496 46900 21548
rect 49332 21564 49384 21616
rect 51448 21564 51500 21616
rect 53380 21632 53432 21684
rect 54392 21632 54444 21684
rect 55036 21632 55088 21684
rect 55864 21632 55916 21684
rect 57520 21675 57572 21684
rect 57520 21641 57529 21675
rect 57529 21641 57563 21675
rect 57563 21641 57572 21675
rect 57520 21632 57572 21641
rect 53656 21564 53708 21616
rect 54668 21564 54720 21616
rect 55128 21564 55180 21616
rect 56692 21607 56744 21616
rect 56692 21573 56701 21607
rect 56701 21573 56735 21607
rect 56735 21573 56744 21607
rect 56692 21564 56744 21573
rect 56968 21564 57020 21616
rect 43076 21428 43128 21480
rect 44180 21428 44232 21480
rect 45008 21428 45060 21480
rect 47492 21428 47544 21480
rect 47952 21428 48004 21480
rect 48872 21428 48924 21480
rect 30104 21335 30156 21344
rect 30104 21301 30113 21335
rect 30113 21301 30147 21335
rect 30147 21301 30156 21335
rect 30104 21292 30156 21301
rect 31576 21292 31628 21344
rect 33140 21360 33192 21412
rect 34336 21360 34388 21412
rect 32864 21292 32916 21344
rect 35072 21292 35124 21344
rect 39672 21360 39724 21412
rect 40316 21360 40368 21412
rect 41236 21360 41288 21412
rect 42156 21403 42208 21412
rect 42156 21369 42165 21403
rect 42165 21369 42199 21403
rect 42199 21369 42208 21403
rect 42156 21360 42208 21369
rect 36084 21292 36136 21344
rect 41696 21335 41748 21344
rect 41696 21301 41705 21335
rect 41705 21301 41739 21335
rect 41739 21301 41748 21335
rect 41696 21292 41748 21301
rect 44548 21292 44600 21344
rect 46112 21335 46164 21344
rect 46112 21301 46121 21335
rect 46121 21301 46155 21335
rect 46155 21301 46164 21335
rect 46112 21292 46164 21301
rect 49424 21428 49476 21480
rect 50252 21471 50304 21480
rect 50252 21437 50261 21471
rect 50261 21437 50295 21471
rect 50295 21437 50304 21471
rect 50252 21428 50304 21437
rect 49056 21360 49108 21412
rect 52460 21496 52512 21548
rect 54484 21496 54536 21548
rect 50988 21428 51040 21480
rect 54944 21539 54996 21548
rect 54944 21505 54953 21539
rect 54953 21505 54987 21539
rect 54987 21505 54996 21539
rect 54944 21496 54996 21505
rect 55036 21496 55088 21548
rect 55588 21539 55640 21548
rect 55588 21505 55597 21539
rect 55597 21505 55631 21539
rect 55631 21505 55640 21539
rect 55588 21496 55640 21505
rect 51540 21292 51592 21344
rect 51724 21292 51776 21344
rect 52368 21360 52420 21412
rect 54576 21360 54628 21412
rect 52184 21335 52236 21344
rect 52184 21301 52193 21335
rect 52193 21301 52227 21335
rect 52227 21301 52236 21335
rect 52184 21292 52236 21301
rect 53564 21292 53616 21344
rect 54484 21335 54536 21344
rect 54484 21301 54493 21335
rect 54493 21301 54527 21335
rect 54527 21301 54536 21335
rect 54484 21292 54536 21301
rect 55312 21335 55364 21344
rect 55312 21301 55321 21335
rect 55321 21301 55355 21335
rect 55355 21301 55364 21335
rect 55312 21292 55364 21301
rect 55680 21292 55732 21344
rect 56876 21539 56928 21548
rect 56876 21505 56885 21539
rect 56885 21505 56919 21539
rect 56919 21505 56928 21539
rect 56876 21496 56928 21505
rect 56692 21428 56744 21480
rect 58440 21539 58492 21548
rect 58440 21505 58449 21539
rect 58449 21505 58483 21539
rect 58483 21505 58492 21539
rect 58440 21496 58492 21505
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 20168 21088 20220 21140
rect 18972 21063 19024 21072
rect 18972 21029 18981 21063
rect 18981 21029 19015 21063
rect 19015 21029 19024 21063
rect 18972 21020 19024 21029
rect 19248 20995 19300 21004
rect 19248 20961 19257 20995
rect 19257 20961 19291 20995
rect 19291 20961 19300 20995
rect 19248 20952 19300 20961
rect 19984 20952 20036 21004
rect 25872 21131 25924 21140
rect 25872 21097 25881 21131
rect 25881 21097 25915 21131
rect 25915 21097 25924 21131
rect 25872 21088 25924 21097
rect 26608 21088 26660 21140
rect 30104 21088 30156 21140
rect 30288 21088 30340 21140
rect 22100 21020 22152 21072
rect 19800 20816 19852 20868
rect 21824 20884 21876 20936
rect 22284 20995 22336 21004
rect 22284 20961 22293 20995
rect 22293 20961 22327 20995
rect 22327 20961 22336 20995
rect 22284 20952 22336 20961
rect 24124 21020 24176 21072
rect 25504 20952 25556 21004
rect 22376 20927 22428 20936
rect 22376 20893 22385 20927
rect 22385 20893 22419 20927
rect 22419 20893 22428 20927
rect 22376 20884 22428 20893
rect 24584 20884 24636 20936
rect 26240 21020 26292 21072
rect 26056 20952 26108 21004
rect 20996 20791 21048 20800
rect 20996 20757 21005 20791
rect 21005 20757 21039 20791
rect 21039 20757 21048 20791
rect 20996 20748 21048 20757
rect 22192 20748 22244 20800
rect 23204 20816 23256 20868
rect 24124 20816 24176 20868
rect 24860 20816 24912 20868
rect 25596 20816 25648 20868
rect 23664 20748 23716 20800
rect 25872 20748 25924 20800
rect 27528 20952 27580 21004
rect 27160 20884 27212 20936
rect 30012 20995 30064 21004
rect 30012 20961 30021 20995
rect 30021 20961 30055 20995
rect 30055 20961 30064 20995
rect 30012 20952 30064 20961
rect 31576 20995 31628 21004
rect 31576 20961 31585 20995
rect 31585 20961 31619 20995
rect 31619 20961 31628 20995
rect 31576 20952 31628 20961
rect 34152 21088 34204 21140
rect 34428 21088 34480 21140
rect 35164 21088 35216 21140
rect 35348 21088 35400 21140
rect 36728 21088 36780 21140
rect 38660 21088 38712 21140
rect 34336 20952 34388 21004
rect 34704 20952 34756 21004
rect 29644 20884 29696 20936
rect 29736 20927 29788 20936
rect 29736 20893 29745 20927
rect 29745 20893 29779 20927
rect 29779 20893 29788 20927
rect 29736 20884 29788 20893
rect 29828 20927 29880 20936
rect 29828 20893 29837 20927
rect 29837 20893 29871 20927
rect 29871 20893 29880 20927
rect 29828 20884 29880 20893
rect 27804 20816 27856 20868
rect 28632 20816 28684 20868
rect 28816 20816 28868 20868
rect 31208 20927 31260 20936
rect 31208 20893 31217 20927
rect 31217 20893 31251 20927
rect 31251 20893 31260 20927
rect 31208 20884 31260 20893
rect 31116 20816 31168 20868
rect 27712 20748 27764 20800
rect 29920 20748 29972 20800
rect 31300 20748 31352 20800
rect 31944 20816 31996 20868
rect 36268 20952 36320 21004
rect 36360 20952 36412 21004
rect 40592 21020 40644 21072
rect 40868 21020 40920 21072
rect 42892 21088 42944 21140
rect 44088 21088 44140 21140
rect 45008 21131 45060 21140
rect 45008 21097 45017 21131
rect 45017 21097 45051 21131
rect 45051 21097 45060 21131
rect 45008 21088 45060 21097
rect 45468 21131 45520 21140
rect 45468 21097 45477 21131
rect 45477 21097 45511 21131
rect 45511 21097 45520 21131
rect 45468 21088 45520 21097
rect 47492 21131 47544 21140
rect 47492 21097 47501 21131
rect 47501 21097 47535 21131
rect 47535 21097 47544 21131
rect 47492 21088 47544 21097
rect 47952 21131 48004 21140
rect 47952 21097 47961 21131
rect 47961 21097 47995 21131
rect 47995 21097 48004 21131
rect 47952 21088 48004 21097
rect 48320 21088 48372 21140
rect 49332 21088 49384 21140
rect 43996 21063 44048 21072
rect 43996 21029 44005 21063
rect 44005 21029 44039 21063
rect 44039 21029 44048 21063
rect 43996 21020 44048 21029
rect 40040 20952 40092 21004
rect 41696 20952 41748 21004
rect 41880 20952 41932 21004
rect 35164 20884 35216 20936
rect 35808 20884 35860 20936
rect 37924 20927 37976 20936
rect 37924 20893 37933 20927
rect 37933 20893 37967 20927
rect 37967 20893 37976 20927
rect 37924 20884 37976 20893
rect 39304 20884 39356 20936
rect 40500 20884 40552 20936
rect 42892 20927 42944 20936
rect 42892 20893 42901 20927
rect 42901 20893 42935 20927
rect 42935 20893 42944 20927
rect 42892 20884 42944 20893
rect 36820 20859 36872 20868
rect 36820 20825 36829 20859
rect 36829 20825 36863 20859
rect 36863 20825 36872 20859
rect 36820 20816 36872 20825
rect 38200 20859 38252 20868
rect 38200 20825 38209 20859
rect 38209 20825 38243 20859
rect 38243 20825 38252 20859
rect 38200 20816 38252 20825
rect 34520 20748 34572 20800
rect 34704 20748 34756 20800
rect 38476 20748 38528 20800
rect 42708 20859 42760 20868
rect 42708 20825 42717 20859
rect 42717 20825 42751 20859
rect 42751 20825 42760 20859
rect 42708 20816 42760 20825
rect 39856 20791 39908 20800
rect 39856 20757 39865 20791
rect 39865 20757 39899 20791
rect 39899 20757 39908 20791
rect 39856 20748 39908 20757
rect 42984 20748 43036 20800
rect 44272 21020 44324 21072
rect 47584 21020 47636 21072
rect 48412 21020 48464 21072
rect 44272 20927 44324 20936
rect 44272 20893 44279 20927
rect 44279 20893 44324 20927
rect 44272 20884 44324 20893
rect 44456 20927 44508 20936
rect 44456 20893 44465 20927
rect 44465 20893 44499 20927
rect 44499 20893 44508 20927
rect 44456 20884 44508 20893
rect 44640 20884 44692 20936
rect 44732 20884 44784 20936
rect 45284 20927 45336 20936
rect 45284 20893 45293 20927
rect 45293 20893 45327 20927
rect 45327 20893 45336 20927
rect 45284 20884 45336 20893
rect 46112 20884 46164 20936
rect 46848 20927 46900 20936
rect 46848 20893 46857 20927
rect 46857 20893 46891 20927
rect 46891 20893 46900 20927
rect 46848 20884 46900 20893
rect 44364 20859 44416 20868
rect 44364 20825 44373 20859
rect 44373 20825 44407 20859
rect 44407 20825 44416 20859
rect 44364 20816 44416 20825
rect 44732 20748 44784 20800
rect 44916 20816 44968 20868
rect 47492 20884 47544 20936
rect 47676 20927 47728 20936
rect 47676 20893 47685 20927
rect 47685 20893 47719 20927
rect 47719 20893 47728 20927
rect 47676 20884 47728 20893
rect 47768 20927 47820 20936
rect 47768 20893 47777 20927
rect 47777 20893 47811 20927
rect 47811 20893 47820 20927
rect 47768 20884 47820 20893
rect 48872 20952 48924 21004
rect 48596 20927 48648 20936
rect 48596 20893 48600 20927
rect 48600 20893 48634 20927
rect 48634 20893 48648 20927
rect 48596 20884 48648 20893
rect 48688 20927 48740 20936
rect 48688 20893 48697 20927
rect 48697 20893 48731 20927
rect 48731 20893 48740 20927
rect 48688 20884 48740 20893
rect 48780 20927 48832 20936
rect 48780 20893 48789 20927
rect 48789 20893 48823 20927
rect 48823 20893 48832 20927
rect 48780 20884 48832 20893
rect 48964 20927 49016 20936
rect 48964 20893 48972 20927
rect 48972 20893 49006 20927
rect 49006 20893 49016 20927
rect 48964 20884 49016 20893
rect 49056 20927 49108 20936
rect 49056 20893 49065 20927
rect 49065 20893 49099 20927
rect 49099 20893 49108 20927
rect 49056 20884 49108 20893
rect 49148 20927 49200 20936
rect 49148 20893 49157 20927
rect 49157 20893 49191 20927
rect 49191 20893 49200 20927
rect 49148 20884 49200 20893
rect 49332 20927 49384 20936
rect 49332 20893 49339 20927
rect 49339 20893 49384 20927
rect 49332 20884 49384 20893
rect 49516 21020 49568 21072
rect 50988 21088 51040 21140
rect 51264 21131 51316 21140
rect 51264 21097 51273 21131
rect 51273 21097 51307 21131
rect 51307 21097 51316 21131
rect 51264 21088 51316 21097
rect 52184 21088 52236 21140
rect 52460 21131 52512 21140
rect 52460 21097 52469 21131
rect 52469 21097 52503 21131
rect 52503 21097 52512 21131
rect 52460 21088 52512 21097
rect 49792 20884 49844 20936
rect 49976 20884 50028 20936
rect 50528 20927 50580 20936
rect 50528 20893 50537 20927
rect 50537 20893 50571 20927
rect 50571 20893 50580 20927
rect 50528 20884 50580 20893
rect 46296 20748 46348 20800
rect 47308 20816 47360 20868
rect 50160 20816 50212 20868
rect 50804 20927 50856 20936
rect 50804 20893 50813 20927
rect 50813 20893 50847 20927
rect 50847 20893 50856 20927
rect 50804 20884 50856 20893
rect 51356 20995 51408 21004
rect 51356 20961 51365 20995
rect 51365 20961 51399 20995
rect 51399 20961 51408 20995
rect 51356 20952 51408 20961
rect 54484 20952 54536 21004
rect 54944 20952 54996 21004
rect 47492 20748 47544 20800
rect 48872 20748 48924 20800
rect 49240 20748 49292 20800
rect 49792 20748 49844 20800
rect 50252 20748 50304 20800
rect 51264 20816 51316 20868
rect 51908 20927 51960 20936
rect 51908 20893 51918 20927
rect 51918 20893 51952 20927
rect 51952 20893 51960 20927
rect 51908 20884 51960 20893
rect 52092 20927 52144 20936
rect 52092 20893 52101 20927
rect 52101 20893 52135 20927
rect 52135 20893 52144 20927
rect 52092 20884 52144 20893
rect 52184 20927 52236 20936
rect 52184 20893 52193 20927
rect 52193 20893 52227 20927
rect 52227 20893 52236 20927
rect 52184 20884 52236 20893
rect 52460 20884 52512 20936
rect 52644 20884 52696 20936
rect 56140 20952 56192 21004
rect 56692 20884 56744 20936
rect 51816 20748 51868 20800
rect 54392 20816 54444 20868
rect 55128 20816 55180 20868
rect 55956 20859 56008 20868
rect 55956 20825 55965 20859
rect 55965 20825 55999 20859
rect 55999 20825 56008 20859
rect 55956 20816 56008 20825
rect 57796 20859 57848 20868
rect 57796 20825 57805 20859
rect 57805 20825 57839 20859
rect 57839 20825 57848 20859
rect 57796 20816 57848 20825
rect 53472 20748 53524 20800
rect 54484 20748 54536 20800
rect 54760 20748 54812 20800
rect 55588 20748 55640 20800
rect 56048 20748 56100 20800
rect 56232 20791 56284 20800
rect 56232 20757 56241 20791
rect 56241 20757 56275 20791
rect 56275 20757 56284 20791
rect 56232 20748 56284 20757
rect 56324 20791 56376 20800
rect 56324 20757 56333 20791
rect 56333 20757 56367 20791
rect 56367 20757 56376 20791
rect 56324 20748 56376 20757
rect 4874 20646 4926 20698
rect 4938 20646 4990 20698
rect 5002 20646 5054 20698
rect 5066 20646 5118 20698
rect 5130 20646 5182 20698
rect 35594 20646 35646 20698
rect 35658 20646 35710 20698
rect 35722 20646 35774 20698
rect 35786 20646 35838 20698
rect 35850 20646 35902 20698
rect 19156 20544 19208 20596
rect 19800 20408 19852 20460
rect 20536 20544 20588 20596
rect 20352 20476 20404 20528
rect 22100 20476 22152 20528
rect 22560 20476 22612 20528
rect 23664 20587 23716 20596
rect 23664 20553 23673 20587
rect 23673 20553 23707 20587
rect 23707 20553 23716 20587
rect 23664 20544 23716 20553
rect 23848 20451 23900 20460
rect 23848 20417 23857 20451
rect 23857 20417 23891 20451
rect 23891 20417 23900 20451
rect 23848 20408 23900 20417
rect 24032 20451 24084 20460
rect 24032 20417 24041 20451
rect 24041 20417 24075 20451
rect 24075 20417 24084 20451
rect 24032 20408 24084 20417
rect 24124 20451 24176 20460
rect 24124 20417 24133 20451
rect 24133 20417 24167 20451
rect 24167 20417 24176 20451
rect 24124 20408 24176 20417
rect 18788 20383 18840 20392
rect 18788 20349 18797 20383
rect 18797 20349 18831 20383
rect 18831 20349 18840 20383
rect 18788 20340 18840 20349
rect 20444 20340 20496 20392
rect 22192 20340 22244 20392
rect 23572 20383 23624 20392
rect 23572 20349 23581 20383
rect 23581 20349 23615 20383
rect 23615 20349 23624 20383
rect 25228 20408 25280 20460
rect 23572 20340 23624 20349
rect 25136 20340 25188 20392
rect 25412 20544 25464 20596
rect 26700 20544 26752 20596
rect 27344 20544 27396 20596
rect 26332 20476 26384 20528
rect 26976 20476 27028 20528
rect 28540 20519 28592 20528
rect 28540 20485 28549 20519
rect 28549 20485 28583 20519
rect 28583 20485 28592 20519
rect 28540 20476 28592 20485
rect 29828 20544 29880 20596
rect 30932 20544 30984 20596
rect 25412 20451 25464 20460
rect 25412 20417 25421 20451
rect 25421 20417 25455 20451
rect 25455 20417 25464 20451
rect 25412 20408 25464 20417
rect 25504 20451 25556 20460
rect 25504 20417 25514 20451
rect 25514 20417 25548 20451
rect 25548 20417 25556 20451
rect 25504 20408 25556 20417
rect 26148 20451 26200 20460
rect 26148 20417 26157 20451
rect 26157 20417 26191 20451
rect 26191 20417 26200 20451
rect 26148 20408 26200 20417
rect 27712 20408 27764 20460
rect 28724 20408 28776 20460
rect 29092 20451 29144 20460
rect 29092 20417 29101 20451
rect 29101 20417 29135 20451
rect 29135 20417 29144 20451
rect 29092 20408 29144 20417
rect 29276 20519 29328 20528
rect 29276 20485 29285 20519
rect 29285 20485 29319 20519
rect 29319 20485 29328 20519
rect 29276 20476 29328 20485
rect 29920 20519 29972 20528
rect 29920 20485 29929 20519
rect 29929 20485 29963 20519
rect 29963 20485 29972 20519
rect 29920 20476 29972 20485
rect 31300 20476 31352 20528
rect 34796 20544 34848 20596
rect 29368 20451 29420 20460
rect 29368 20417 29377 20451
rect 29377 20417 29411 20451
rect 29411 20417 29420 20451
rect 29368 20408 29420 20417
rect 34796 20408 34848 20460
rect 27804 20340 27856 20392
rect 28816 20340 28868 20392
rect 29644 20383 29696 20392
rect 29644 20349 29653 20383
rect 29653 20349 29687 20383
rect 29687 20349 29696 20383
rect 29644 20340 29696 20349
rect 19524 20204 19576 20256
rect 24768 20247 24820 20256
rect 24768 20213 24777 20247
rect 24777 20213 24811 20247
rect 24811 20213 24820 20247
rect 24768 20204 24820 20213
rect 25228 20204 25280 20256
rect 25596 20204 25648 20256
rect 26516 20272 26568 20324
rect 28632 20272 28684 20324
rect 30932 20340 30984 20392
rect 31116 20340 31168 20392
rect 31392 20383 31444 20392
rect 31392 20349 31401 20383
rect 31401 20349 31435 20383
rect 31435 20349 31444 20383
rect 31392 20340 31444 20349
rect 33600 20383 33652 20392
rect 33600 20349 33609 20383
rect 33609 20349 33643 20383
rect 33643 20349 33652 20383
rect 33600 20340 33652 20349
rect 34704 20340 34756 20392
rect 35164 20340 35216 20392
rect 35348 20340 35400 20392
rect 35716 20408 35768 20460
rect 36452 20544 36504 20596
rect 38200 20544 38252 20596
rect 36268 20408 36320 20460
rect 39028 20544 39080 20596
rect 40224 20544 40276 20596
rect 39856 20476 39908 20528
rect 39304 20451 39356 20460
rect 39304 20417 39313 20451
rect 39313 20417 39347 20451
rect 39347 20417 39356 20451
rect 42616 20544 42668 20596
rect 42708 20544 42760 20596
rect 43076 20587 43128 20596
rect 43076 20553 43085 20587
rect 43085 20553 43119 20587
rect 43119 20553 43128 20587
rect 43076 20544 43128 20553
rect 43168 20544 43220 20596
rect 42800 20519 42852 20528
rect 42800 20485 42809 20519
rect 42809 20485 42843 20519
rect 42843 20485 42852 20519
rect 42800 20476 42852 20485
rect 39304 20408 39356 20417
rect 42616 20451 42668 20460
rect 42616 20417 42625 20451
rect 42625 20417 42659 20451
rect 42659 20417 42668 20451
rect 42616 20408 42668 20417
rect 42892 20408 42944 20460
rect 42984 20451 43036 20460
rect 42984 20417 42993 20451
rect 42993 20417 43027 20451
rect 43027 20417 43036 20451
rect 42984 20408 43036 20417
rect 44272 20544 44324 20596
rect 44916 20519 44968 20528
rect 44916 20485 44925 20519
rect 44925 20485 44959 20519
rect 44959 20485 44968 20519
rect 44916 20476 44968 20485
rect 45100 20544 45152 20596
rect 47124 20587 47176 20596
rect 47124 20553 47133 20587
rect 47133 20553 47167 20587
rect 47167 20553 47176 20587
rect 47124 20544 47176 20553
rect 47860 20544 47912 20596
rect 48044 20544 48096 20596
rect 48228 20544 48280 20596
rect 48872 20544 48924 20596
rect 49332 20544 49384 20596
rect 49608 20587 49660 20596
rect 49608 20553 49617 20587
rect 49617 20553 49651 20587
rect 49651 20553 49660 20587
rect 49608 20544 49660 20553
rect 26056 20247 26108 20256
rect 26056 20213 26065 20247
rect 26065 20213 26099 20247
rect 26099 20213 26108 20247
rect 26056 20204 26108 20213
rect 26608 20204 26660 20256
rect 27068 20204 27120 20256
rect 29368 20204 29420 20256
rect 39120 20340 39172 20392
rect 39488 20383 39540 20392
rect 39488 20349 39497 20383
rect 39497 20349 39531 20383
rect 39531 20349 39540 20383
rect 39488 20340 39540 20349
rect 40500 20383 40552 20392
rect 40500 20349 40509 20383
rect 40509 20349 40543 20383
rect 40543 20349 40552 20383
rect 40500 20340 40552 20349
rect 41328 20340 41380 20392
rect 43536 20408 43588 20460
rect 44364 20408 44416 20460
rect 44824 20408 44876 20460
rect 46756 20476 46808 20528
rect 41880 20272 41932 20324
rect 43168 20272 43220 20324
rect 47584 20451 47636 20460
rect 47584 20417 47593 20451
rect 47593 20417 47627 20451
rect 47627 20417 47636 20451
rect 47584 20408 47636 20417
rect 47768 20451 47820 20460
rect 47768 20417 47775 20451
rect 47775 20417 47820 20451
rect 47768 20408 47820 20417
rect 47860 20451 47912 20460
rect 47860 20417 47869 20451
rect 47869 20417 47903 20451
rect 47903 20417 47912 20451
rect 47860 20408 47912 20417
rect 47124 20340 47176 20392
rect 48136 20340 48188 20392
rect 45652 20272 45704 20324
rect 47032 20272 47084 20324
rect 47676 20272 47728 20324
rect 49884 20519 49936 20528
rect 49884 20485 49893 20519
rect 49893 20485 49927 20519
rect 49927 20485 49936 20519
rect 49884 20476 49936 20485
rect 49976 20476 50028 20528
rect 52460 20476 52512 20528
rect 48320 20272 48372 20324
rect 48688 20451 48740 20460
rect 48688 20417 48697 20451
rect 48697 20417 48731 20451
rect 48731 20417 48740 20451
rect 48688 20408 48740 20417
rect 48780 20451 48832 20460
rect 48780 20417 48813 20451
rect 48813 20417 48832 20451
rect 48780 20408 48832 20417
rect 49332 20451 49384 20460
rect 49332 20417 49341 20451
rect 49341 20417 49375 20451
rect 49375 20417 49384 20451
rect 49332 20408 49384 20417
rect 50068 20451 50120 20460
rect 50068 20417 50077 20451
rect 50077 20417 50111 20451
rect 50111 20417 50120 20451
rect 50068 20408 50120 20417
rect 50528 20408 50580 20460
rect 53840 20408 53892 20460
rect 54576 20476 54628 20528
rect 56324 20544 56376 20596
rect 57796 20544 57848 20596
rect 54944 20408 54996 20460
rect 55404 20451 55456 20460
rect 55404 20417 55413 20451
rect 55413 20417 55447 20451
rect 55447 20417 55456 20451
rect 55404 20408 55456 20417
rect 56324 20408 56376 20460
rect 49424 20340 49476 20392
rect 50896 20340 50948 20392
rect 54852 20340 54904 20392
rect 48596 20272 48648 20324
rect 37188 20204 37240 20256
rect 41236 20204 41288 20256
rect 42432 20247 42484 20256
rect 42432 20213 42441 20247
rect 42441 20213 42475 20247
rect 42475 20213 42484 20247
rect 42432 20204 42484 20213
rect 42800 20204 42852 20256
rect 43536 20204 43588 20256
rect 45192 20204 45244 20256
rect 45560 20247 45612 20256
rect 45560 20213 45569 20247
rect 45569 20213 45603 20247
rect 45603 20213 45612 20247
rect 45560 20204 45612 20213
rect 47768 20204 47820 20256
rect 48872 20272 48924 20324
rect 49516 20315 49568 20324
rect 49516 20281 49525 20315
rect 49525 20281 49559 20315
rect 49559 20281 49568 20315
rect 49516 20272 49568 20281
rect 53380 20272 53432 20324
rect 55956 20340 56008 20392
rect 55312 20272 55364 20324
rect 50436 20204 50488 20256
rect 53288 20204 53340 20256
rect 53656 20204 53708 20256
rect 53932 20204 53984 20256
rect 55220 20247 55272 20256
rect 55220 20213 55229 20247
rect 55229 20213 55263 20247
rect 55263 20213 55272 20247
rect 55220 20204 55272 20213
rect 55588 20247 55640 20256
rect 55588 20213 55597 20247
rect 55597 20213 55631 20247
rect 55631 20213 55640 20247
rect 55588 20204 55640 20213
rect 56048 20247 56100 20256
rect 56048 20213 56057 20247
rect 56057 20213 56091 20247
rect 56091 20213 56100 20247
rect 56048 20204 56100 20213
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 25412 20043 25464 20052
rect 25412 20009 25421 20043
rect 25421 20009 25455 20043
rect 25455 20009 25464 20043
rect 25412 20000 25464 20009
rect 25688 20000 25740 20052
rect 26056 20000 26108 20052
rect 27068 20000 27120 20052
rect 29184 20000 29236 20052
rect 22652 19932 22704 19984
rect 26424 19932 26476 19984
rect 25504 19864 25556 19916
rect 15200 19796 15252 19848
rect 24860 19839 24912 19848
rect 24860 19805 24869 19839
rect 24869 19805 24903 19839
rect 24903 19805 24912 19839
rect 24860 19796 24912 19805
rect 25044 19839 25096 19848
rect 25044 19805 25053 19839
rect 25053 19805 25087 19839
rect 25087 19805 25096 19839
rect 25044 19796 25096 19805
rect 25136 19771 25188 19780
rect 25136 19737 25145 19771
rect 25145 19737 25179 19771
rect 25179 19737 25188 19771
rect 25136 19728 25188 19737
rect 25320 19796 25372 19848
rect 26608 19864 26660 19916
rect 28724 19932 28776 19984
rect 25688 19728 25740 19780
rect 848 19660 900 19712
rect 26332 19839 26384 19848
rect 26332 19805 26346 19839
rect 26346 19805 26380 19839
rect 26380 19805 26384 19839
rect 27712 19864 27764 19916
rect 29644 19864 29696 19916
rect 31208 19932 31260 19984
rect 31576 19932 31628 19984
rect 34060 20000 34112 20052
rect 34704 20043 34756 20052
rect 34704 20009 34713 20043
rect 34713 20009 34747 20043
rect 34747 20009 34756 20043
rect 34704 20000 34756 20009
rect 34796 20000 34848 20052
rect 36452 20000 36504 20052
rect 36636 20000 36688 20052
rect 41236 20043 41288 20052
rect 41236 20009 41245 20043
rect 41245 20009 41279 20043
rect 41279 20009 41288 20043
rect 41236 20000 41288 20009
rect 41328 20043 41380 20052
rect 41328 20009 41337 20043
rect 41337 20009 41371 20043
rect 41371 20009 41380 20043
rect 41328 20000 41380 20009
rect 48320 20000 48372 20052
rect 49056 20000 49108 20052
rect 49240 20000 49292 20052
rect 49884 20000 49936 20052
rect 50436 20000 50488 20052
rect 26332 19796 26384 19805
rect 28816 19796 28868 19848
rect 30656 19796 30708 19848
rect 32036 19864 32088 19916
rect 31392 19839 31444 19848
rect 31392 19805 31401 19839
rect 31401 19805 31435 19839
rect 31435 19805 31444 19839
rect 31392 19796 31444 19805
rect 31576 19839 31628 19848
rect 31576 19805 31621 19839
rect 31621 19805 31628 19839
rect 31576 19796 31628 19805
rect 31760 19839 31812 19848
rect 31760 19805 31769 19839
rect 31769 19805 31803 19839
rect 31803 19805 31812 19839
rect 31760 19796 31812 19805
rect 34796 19864 34848 19916
rect 26608 19771 26660 19780
rect 26608 19737 26617 19771
rect 26617 19737 26651 19771
rect 26651 19737 26660 19771
rect 26608 19728 26660 19737
rect 27896 19728 27948 19780
rect 28724 19728 28776 19780
rect 29552 19728 29604 19780
rect 30840 19728 30892 19780
rect 26332 19660 26384 19712
rect 26424 19660 26476 19712
rect 28540 19660 28592 19712
rect 28908 19660 28960 19712
rect 29828 19703 29880 19712
rect 29828 19669 29837 19703
rect 29837 19669 29871 19703
rect 29871 19669 29880 19703
rect 29828 19660 29880 19669
rect 30380 19660 30432 19712
rect 34244 19771 34296 19780
rect 34244 19737 34253 19771
rect 34253 19737 34287 19771
rect 34287 19737 34296 19771
rect 34244 19728 34296 19737
rect 32220 19660 32272 19712
rect 34520 19839 34572 19848
rect 34520 19805 34529 19839
rect 34529 19805 34563 19839
rect 34563 19805 34572 19839
rect 34520 19796 34572 19805
rect 34612 19796 34664 19848
rect 34704 19796 34756 19848
rect 35440 19932 35492 19984
rect 51264 20000 51316 20052
rect 42064 19932 42116 19984
rect 48228 19932 48280 19984
rect 50988 19932 51040 19984
rect 35348 19796 35400 19848
rect 35716 19839 35768 19848
rect 35716 19805 35725 19839
rect 35725 19805 35759 19839
rect 35759 19805 35768 19839
rect 35716 19796 35768 19805
rect 36084 19796 36136 19848
rect 37924 19864 37976 19916
rect 44180 19864 44232 19916
rect 46388 19864 46440 19916
rect 46848 19864 46900 19916
rect 35624 19771 35676 19780
rect 35624 19737 35633 19771
rect 35633 19737 35667 19771
rect 35667 19737 35676 19771
rect 35624 19728 35676 19737
rect 34612 19660 34664 19712
rect 36084 19660 36136 19712
rect 36912 19839 36964 19848
rect 36912 19805 36921 19839
rect 36921 19805 36955 19839
rect 36955 19805 36964 19839
rect 36912 19796 36964 19805
rect 38476 19796 38528 19848
rect 39488 19839 39540 19848
rect 36268 19771 36320 19780
rect 36268 19737 36277 19771
rect 36277 19737 36311 19771
rect 36311 19737 36320 19771
rect 36268 19728 36320 19737
rect 36452 19728 36504 19780
rect 37372 19771 37424 19780
rect 37372 19737 37381 19771
rect 37381 19737 37415 19771
rect 37415 19737 37424 19771
rect 37372 19728 37424 19737
rect 39488 19805 39497 19839
rect 39497 19805 39531 19839
rect 39531 19805 39540 19839
rect 39488 19796 39540 19805
rect 41512 19839 41564 19848
rect 39120 19728 39172 19780
rect 41052 19728 41104 19780
rect 41512 19805 41521 19839
rect 41521 19805 41555 19839
rect 41555 19805 41564 19839
rect 41512 19796 41564 19805
rect 41696 19796 41748 19848
rect 41880 19839 41932 19848
rect 41880 19805 41889 19839
rect 41889 19805 41923 19839
rect 41923 19805 41932 19839
rect 41880 19796 41932 19805
rect 45192 19839 45244 19848
rect 45192 19805 45201 19839
rect 45201 19805 45235 19839
rect 45235 19805 45244 19839
rect 45192 19796 45244 19805
rect 45376 19839 45428 19848
rect 45376 19805 45385 19839
rect 45385 19805 45419 19839
rect 45419 19805 45428 19839
rect 45376 19796 45428 19805
rect 45468 19839 45520 19848
rect 45468 19805 45477 19839
rect 45477 19805 45511 19839
rect 45511 19805 45520 19839
rect 45468 19796 45520 19805
rect 46664 19796 46716 19848
rect 47768 19839 47820 19848
rect 47768 19805 47777 19839
rect 47777 19805 47811 19839
rect 47811 19805 47820 19839
rect 47768 19796 47820 19805
rect 42432 19728 42484 19780
rect 42708 19728 42760 19780
rect 45560 19771 45612 19780
rect 45560 19737 45569 19771
rect 45569 19737 45603 19771
rect 45603 19737 45612 19771
rect 45560 19728 45612 19737
rect 47492 19728 47544 19780
rect 48136 19796 48188 19848
rect 48412 19839 48464 19848
rect 48412 19805 48421 19839
rect 48421 19805 48455 19839
rect 48455 19805 48464 19839
rect 48412 19796 48464 19805
rect 36728 19660 36780 19712
rect 38844 19703 38896 19712
rect 38844 19669 38853 19703
rect 38853 19669 38887 19703
rect 38887 19669 38896 19703
rect 38844 19660 38896 19669
rect 38936 19703 38988 19712
rect 38936 19669 38945 19703
rect 38945 19669 38979 19703
rect 38979 19669 38988 19703
rect 38936 19660 38988 19669
rect 44364 19660 44416 19712
rect 46664 19660 46716 19712
rect 46848 19703 46900 19712
rect 46848 19669 46857 19703
rect 46857 19669 46891 19703
rect 46891 19669 46900 19703
rect 46848 19660 46900 19669
rect 47952 19660 48004 19712
rect 48228 19771 48280 19780
rect 48228 19737 48237 19771
rect 48237 19737 48271 19771
rect 48271 19737 48280 19771
rect 48228 19728 48280 19737
rect 49056 19839 49108 19848
rect 49056 19805 49065 19839
rect 49065 19805 49099 19839
rect 49099 19805 49108 19839
rect 49056 19796 49108 19805
rect 49424 19839 49476 19848
rect 49424 19805 49433 19839
rect 49433 19805 49467 19839
rect 49467 19805 49476 19839
rect 49424 19796 49476 19805
rect 50436 19796 50488 19848
rect 50712 19839 50764 19848
rect 50712 19805 50721 19839
rect 50721 19805 50755 19839
rect 50755 19805 50764 19839
rect 50712 19796 50764 19805
rect 50896 19796 50948 19848
rect 50988 19839 51040 19848
rect 50988 19805 50997 19839
rect 50997 19805 51031 19839
rect 51031 19805 51040 19839
rect 50988 19796 51040 19805
rect 51724 19864 51776 19916
rect 52920 19864 52972 19916
rect 48780 19660 48832 19712
rect 51080 19771 51132 19780
rect 51080 19737 51089 19771
rect 51089 19737 51123 19771
rect 51123 19737 51132 19771
rect 51080 19728 51132 19737
rect 49516 19703 49568 19712
rect 49516 19669 49525 19703
rect 49525 19669 49559 19703
rect 49559 19669 49568 19703
rect 49516 19660 49568 19669
rect 49792 19703 49844 19712
rect 49792 19669 49801 19703
rect 49801 19669 49835 19703
rect 49835 19669 49844 19703
rect 49792 19660 49844 19669
rect 50436 19660 50488 19712
rect 51724 19771 51776 19780
rect 51724 19737 51733 19771
rect 51733 19737 51767 19771
rect 51767 19737 51776 19771
rect 51724 19728 51776 19737
rect 53840 20000 53892 20052
rect 55404 20000 55456 20052
rect 55956 20000 56008 20052
rect 53472 19864 53524 19916
rect 53288 19839 53340 19848
rect 53288 19805 53297 19839
rect 53297 19805 53331 19839
rect 53331 19805 53340 19839
rect 53288 19796 53340 19805
rect 53380 19839 53432 19848
rect 53380 19805 53390 19839
rect 53390 19805 53424 19839
rect 53424 19805 53432 19839
rect 56140 19864 56192 19916
rect 53380 19796 53432 19805
rect 53748 19839 53800 19848
rect 53748 19805 53762 19839
rect 53762 19805 53796 19839
rect 53796 19805 53800 19839
rect 53748 19796 53800 19805
rect 54484 19839 54536 19848
rect 54484 19805 54493 19839
rect 54493 19805 54527 19839
rect 54527 19805 54536 19839
rect 54484 19796 54536 19805
rect 54576 19839 54628 19848
rect 54576 19805 54586 19839
rect 54586 19805 54620 19839
rect 54620 19805 54628 19839
rect 54576 19796 54628 19805
rect 54944 19839 54996 19848
rect 54944 19805 54958 19839
rect 54958 19805 54992 19839
rect 54992 19805 54996 19839
rect 54944 19796 54996 19805
rect 56692 19796 56744 19848
rect 58164 19796 58216 19848
rect 58256 19839 58308 19848
rect 58256 19805 58265 19839
rect 58265 19805 58299 19839
rect 58299 19805 58308 19839
rect 58256 19796 58308 19805
rect 51816 19660 51868 19712
rect 52092 19660 52144 19712
rect 53472 19660 53524 19712
rect 54852 19771 54904 19780
rect 54852 19737 54861 19771
rect 54861 19737 54895 19771
rect 54895 19737 54904 19771
rect 54852 19728 54904 19737
rect 55588 19771 55640 19780
rect 55588 19737 55597 19771
rect 55597 19737 55631 19771
rect 55631 19737 55640 19771
rect 55588 19728 55640 19737
rect 55956 19660 56008 19712
rect 57888 19660 57940 19712
rect 58440 19703 58492 19712
rect 58440 19669 58449 19703
rect 58449 19669 58483 19703
rect 58483 19669 58492 19703
rect 58440 19660 58492 19669
rect 4874 19558 4926 19610
rect 4938 19558 4990 19610
rect 5002 19558 5054 19610
rect 5066 19558 5118 19610
rect 5130 19558 5182 19610
rect 35594 19558 35646 19610
rect 35658 19558 35710 19610
rect 35722 19558 35774 19610
rect 35786 19558 35838 19610
rect 35850 19558 35902 19610
rect 15200 19456 15252 19508
rect 16120 19363 16172 19372
rect 16120 19329 16138 19363
rect 16138 19329 16172 19363
rect 16120 19320 16172 19329
rect 16672 19320 16724 19372
rect 19340 19456 19392 19508
rect 20076 19456 20128 19508
rect 19892 19388 19944 19440
rect 19524 19320 19576 19372
rect 19616 19363 19668 19372
rect 19616 19329 19625 19363
rect 19625 19329 19659 19363
rect 19659 19329 19668 19363
rect 19616 19320 19668 19329
rect 19800 19363 19852 19372
rect 19800 19329 19809 19363
rect 19809 19329 19843 19363
rect 19843 19329 19852 19363
rect 19800 19320 19852 19329
rect 20444 19388 20496 19440
rect 22192 19363 22244 19372
rect 22192 19329 22203 19363
rect 22203 19329 22244 19363
rect 22192 19320 22244 19329
rect 22376 19363 22428 19372
rect 22376 19329 22385 19363
rect 22385 19329 22419 19363
rect 22419 19329 22428 19363
rect 22376 19320 22428 19329
rect 25688 19456 25740 19508
rect 26148 19456 26200 19508
rect 26240 19456 26292 19508
rect 26884 19456 26936 19508
rect 28172 19456 28224 19508
rect 24768 19388 24820 19440
rect 28540 19456 28592 19508
rect 28816 19456 28868 19508
rect 28908 19499 28960 19508
rect 28908 19465 28917 19499
rect 28917 19465 28951 19499
rect 28951 19465 28960 19499
rect 28908 19456 28960 19465
rect 23020 19363 23072 19372
rect 23020 19329 23029 19363
rect 23029 19329 23063 19363
rect 23063 19329 23072 19363
rect 23020 19320 23072 19329
rect 23112 19363 23164 19372
rect 23112 19329 23121 19363
rect 23121 19329 23155 19363
rect 23155 19329 23164 19363
rect 23112 19320 23164 19329
rect 23296 19320 23348 19372
rect 18144 19252 18196 19304
rect 24584 19295 24636 19304
rect 24584 19261 24593 19295
rect 24593 19261 24627 19295
rect 24627 19261 24636 19295
rect 24584 19252 24636 19261
rect 19340 19184 19392 19236
rect 20076 19227 20128 19236
rect 20076 19193 20085 19227
rect 20085 19193 20119 19227
rect 20119 19193 20128 19227
rect 20076 19184 20128 19193
rect 17592 19116 17644 19168
rect 19248 19159 19300 19168
rect 19248 19125 19257 19159
rect 19257 19125 19291 19159
rect 19291 19125 19300 19159
rect 19248 19116 19300 19125
rect 21916 19116 21968 19168
rect 22100 19116 22152 19168
rect 22560 19116 22612 19168
rect 23020 19116 23072 19168
rect 25872 19184 25924 19236
rect 26516 19363 26568 19372
rect 26516 19329 26525 19363
rect 26525 19329 26559 19363
rect 26559 19329 26568 19363
rect 26516 19320 26568 19329
rect 30288 19388 30340 19440
rect 28724 19363 28776 19372
rect 26608 19252 26660 19304
rect 27252 19252 27304 19304
rect 28724 19329 28733 19363
rect 28733 19329 28767 19363
rect 28767 19329 28776 19363
rect 28724 19320 28776 19329
rect 29736 19320 29788 19372
rect 30196 19320 30248 19372
rect 34244 19456 34296 19508
rect 36268 19456 36320 19508
rect 28632 19252 28684 19304
rect 30564 19252 30616 19304
rect 31484 19363 31536 19372
rect 31484 19329 31493 19363
rect 31493 19329 31527 19363
rect 31527 19329 31536 19363
rect 31484 19320 31536 19329
rect 31668 19320 31720 19372
rect 33600 19320 33652 19372
rect 35348 19388 35400 19440
rect 34428 19320 34480 19372
rect 36084 19320 36136 19372
rect 36360 19320 36412 19372
rect 38108 19363 38160 19372
rect 38108 19329 38117 19363
rect 38117 19329 38151 19363
rect 38151 19329 38160 19363
rect 38108 19320 38160 19329
rect 40500 19456 40552 19508
rect 34520 19295 34572 19304
rect 34520 19261 34529 19295
rect 34529 19261 34563 19295
rect 34563 19261 34572 19295
rect 34520 19252 34572 19261
rect 34704 19252 34756 19304
rect 35440 19252 35492 19304
rect 37372 19252 37424 19304
rect 38016 19252 38068 19304
rect 38936 19320 38988 19372
rect 39120 19363 39172 19372
rect 39120 19329 39129 19363
rect 39129 19329 39163 19363
rect 39163 19329 39172 19363
rect 39120 19320 39172 19329
rect 39212 19363 39264 19372
rect 39212 19329 39221 19363
rect 39221 19329 39255 19363
rect 39255 19329 39264 19363
rect 39212 19320 39264 19329
rect 40040 19320 40092 19372
rect 40224 19320 40276 19372
rect 40684 19388 40736 19440
rect 25044 19116 25096 19168
rect 25964 19116 26016 19168
rect 28264 19184 28316 19236
rect 35532 19184 35584 19236
rect 40408 19184 40460 19236
rect 26976 19159 27028 19168
rect 26976 19125 26985 19159
rect 26985 19125 27019 19159
rect 27019 19125 27028 19159
rect 26976 19116 27028 19125
rect 31024 19116 31076 19168
rect 32496 19116 32548 19168
rect 34888 19116 34940 19168
rect 39488 19116 39540 19168
rect 45468 19456 45520 19508
rect 41328 19388 41380 19440
rect 40960 19320 41012 19372
rect 42156 19320 42208 19372
rect 42892 19320 42944 19372
rect 43720 19320 43772 19372
rect 41236 19252 41288 19304
rect 44364 19295 44416 19304
rect 44364 19261 44373 19295
rect 44373 19261 44407 19295
rect 44407 19261 44416 19295
rect 44364 19252 44416 19261
rect 46664 19431 46716 19440
rect 46664 19397 46673 19431
rect 46673 19397 46707 19431
rect 46707 19397 46716 19431
rect 46664 19388 46716 19397
rect 46940 19456 46992 19508
rect 48044 19456 48096 19508
rect 49332 19456 49384 19508
rect 49516 19456 49568 19508
rect 49884 19456 49936 19508
rect 50068 19456 50120 19508
rect 52920 19499 52972 19508
rect 52920 19465 52929 19499
rect 52929 19465 52963 19499
rect 52963 19465 52972 19499
rect 52920 19456 52972 19465
rect 54944 19456 54996 19508
rect 56784 19456 56836 19508
rect 45468 19295 45520 19304
rect 45468 19261 45477 19295
rect 45477 19261 45511 19295
rect 45511 19261 45520 19295
rect 45468 19252 45520 19261
rect 46388 19320 46440 19372
rect 47032 19363 47084 19372
rect 47032 19329 47041 19363
rect 47041 19329 47075 19363
rect 47075 19329 47084 19363
rect 47032 19320 47084 19329
rect 48780 19320 48832 19372
rect 50252 19388 50304 19440
rect 51356 19388 51408 19440
rect 51448 19388 51500 19440
rect 53932 19388 53984 19440
rect 54116 19388 54168 19440
rect 56600 19320 56652 19372
rect 41144 19184 41196 19236
rect 47124 19252 47176 19304
rect 49424 19252 49476 19304
rect 49700 19295 49752 19304
rect 49700 19261 49709 19295
rect 49709 19261 49743 19295
rect 49743 19261 49752 19295
rect 49700 19252 49752 19261
rect 49976 19295 50028 19304
rect 49976 19261 49985 19295
rect 49985 19261 50019 19295
rect 50019 19261 50028 19295
rect 49976 19252 50028 19261
rect 51172 19252 51224 19304
rect 53656 19295 53708 19304
rect 53656 19261 53665 19295
rect 53665 19261 53699 19295
rect 53699 19261 53708 19295
rect 53656 19252 53708 19261
rect 58256 19252 58308 19304
rect 46848 19184 46900 19236
rect 47400 19184 47452 19236
rect 47768 19227 47820 19236
rect 47768 19193 47777 19227
rect 47777 19193 47811 19227
rect 47811 19193 47820 19227
rect 47768 19184 47820 19193
rect 49608 19184 49660 19236
rect 57060 19184 57112 19236
rect 40960 19116 41012 19168
rect 45284 19116 45336 19168
rect 47032 19116 47084 19168
rect 47492 19116 47544 19168
rect 49148 19116 49200 19168
rect 49240 19159 49292 19168
rect 49240 19125 49249 19159
rect 49249 19125 49283 19159
rect 49283 19125 49292 19159
rect 49240 19116 49292 19125
rect 51540 19159 51592 19168
rect 51540 19125 51549 19159
rect 51549 19125 51583 19159
rect 51583 19125 51592 19159
rect 51540 19116 51592 19125
rect 57428 19159 57480 19168
rect 57428 19125 57437 19159
rect 57437 19125 57471 19159
rect 57471 19125 57480 19159
rect 57428 19116 57480 19125
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 16120 18955 16172 18964
rect 16120 18921 16129 18955
rect 16129 18921 16163 18955
rect 16163 18921 16172 18955
rect 16120 18912 16172 18921
rect 16856 18955 16908 18964
rect 16856 18921 16865 18955
rect 16865 18921 16899 18955
rect 16899 18921 16908 18955
rect 16856 18912 16908 18921
rect 25320 18912 25372 18964
rect 26976 18912 27028 18964
rect 15200 18776 15252 18828
rect 19616 18844 19668 18896
rect 20076 18844 20128 18896
rect 17592 18819 17644 18828
rect 17592 18785 17601 18819
rect 17601 18785 17635 18819
rect 17635 18785 17644 18819
rect 17592 18776 17644 18785
rect 19524 18776 19576 18828
rect 16764 18751 16816 18760
rect 16764 18717 16773 18751
rect 16773 18717 16807 18751
rect 16807 18717 16816 18751
rect 16764 18708 16816 18717
rect 17316 18751 17368 18760
rect 17316 18717 17325 18751
rect 17325 18717 17359 18751
rect 17359 18717 17368 18751
rect 17316 18708 17368 18717
rect 21916 18819 21968 18828
rect 21916 18785 21925 18819
rect 21925 18785 21959 18819
rect 21959 18785 21968 18819
rect 21916 18776 21968 18785
rect 22560 18819 22612 18828
rect 22560 18785 22569 18819
rect 22569 18785 22603 18819
rect 22603 18785 22612 18819
rect 22560 18776 22612 18785
rect 23020 18776 23072 18828
rect 23296 18776 23348 18828
rect 25136 18844 25188 18896
rect 30380 18912 30432 18964
rect 30564 18955 30616 18964
rect 30564 18921 30573 18955
rect 30573 18921 30607 18955
rect 30607 18921 30616 18955
rect 30564 18912 30616 18921
rect 34520 18955 34572 18964
rect 34520 18921 34529 18955
rect 34529 18921 34563 18955
rect 34563 18921 34572 18955
rect 34520 18912 34572 18921
rect 35532 18912 35584 18964
rect 39212 18912 39264 18964
rect 39764 18912 39816 18964
rect 39856 18912 39908 18964
rect 22192 18751 22244 18760
rect 22192 18717 22201 18751
rect 22201 18717 22235 18751
rect 22235 18717 22244 18751
rect 22192 18708 22244 18717
rect 24400 18708 24452 18760
rect 24952 18776 25004 18828
rect 17960 18572 18012 18624
rect 19524 18640 19576 18692
rect 19616 18572 19668 18624
rect 19708 18572 19760 18624
rect 20260 18615 20312 18624
rect 20260 18581 20269 18615
rect 20269 18581 20303 18615
rect 20303 18581 20312 18615
rect 20260 18572 20312 18581
rect 21916 18640 21968 18692
rect 24768 18683 24820 18692
rect 24768 18649 24777 18683
rect 24777 18649 24811 18683
rect 24811 18649 24820 18683
rect 24768 18640 24820 18649
rect 22376 18572 22428 18624
rect 23848 18572 23900 18624
rect 24584 18572 24636 18624
rect 25044 18708 25096 18760
rect 25136 18640 25188 18692
rect 25412 18708 25464 18760
rect 25044 18572 25096 18624
rect 25872 18708 25924 18760
rect 26608 18776 26660 18828
rect 26424 18751 26476 18760
rect 27620 18819 27672 18828
rect 27620 18785 27629 18819
rect 27629 18785 27663 18819
rect 27663 18785 27672 18819
rect 27620 18776 27672 18785
rect 28632 18776 28684 18828
rect 26424 18717 26438 18751
rect 26438 18717 26472 18751
rect 26472 18717 26476 18751
rect 26424 18708 26476 18717
rect 25964 18572 26016 18624
rect 26148 18572 26200 18624
rect 26332 18683 26384 18692
rect 26332 18649 26341 18683
rect 26341 18649 26375 18683
rect 26375 18649 26384 18683
rect 26332 18640 26384 18649
rect 27344 18751 27396 18760
rect 27344 18717 27353 18751
rect 27353 18717 27387 18751
rect 27387 18717 27396 18751
rect 27344 18708 27396 18717
rect 30564 18776 30616 18828
rect 31668 18776 31720 18828
rect 34060 18819 34112 18828
rect 34060 18785 34069 18819
rect 34069 18785 34103 18819
rect 34103 18785 34112 18819
rect 34060 18776 34112 18785
rect 26424 18572 26476 18624
rect 26608 18615 26660 18624
rect 26608 18581 26617 18615
rect 26617 18581 26651 18615
rect 26651 18581 26660 18615
rect 26608 18572 26660 18581
rect 26792 18615 26844 18624
rect 26792 18581 26801 18615
rect 26801 18581 26835 18615
rect 26835 18581 26844 18615
rect 26792 18572 26844 18581
rect 26976 18572 27028 18624
rect 27988 18640 28040 18692
rect 28908 18640 28960 18692
rect 27344 18572 27396 18624
rect 28264 18572 28316 18624
rect 29368 18615 29420 18624
rect 29368 18581 29377 18615
rect 29377 18581 29411 18615
rect 29411 18581 29420 18615
rect 29368 18572 29420 18581
rect 30288 18751 30340 18760
rect 30288 18717 30297 18751
rect 30297 18717 30331 18751
rect 30331 18717 30340 18751
rect 30288 18708 30340 18717
rect 30748 18708 30800 18760
rect 34336 18844 34388 18896
rect 39488 18844 39540 18896
rect 41328 18844 41380 18896
rect 46756 18955 46808 18964
rect 46756 18921 46765 18955
rect 46765 18921 46799 18955
rect 46799 18921 46808 18955
rect 46756 18912 46808 18921
rect 47124 18955 47176 18964
rect 47124 18921 47133 18955
rect 47133 18921 47167 18955
rect 47167 18921 47176 18955
rect 47124 18912 47176 18921
rect 48412 18912 48464 18964
rect 49056 18912 49108 18964
rect 47400 18844 47452 18896
rect 34612 18776 34664 18828
rect 37924 18819 37976 18828
rect 37924 18785 37933 18819
rect 37933 18785 37967 18819
rect 37967 18785 37976 18819
rect 37924 18776 37976 18785
rect 45284 18819 45336 18828
rect 45284 18785 45293 18819
rect 45293 18785 45327 18819
rect 45327 18785 45336 18819
rect 45284 18776 45336 18785
rect 49240 18844 49292 18896
rect 49700 18912 49752 18964
rect 49976 18912 50028 18964
rect 51724 18912 51776 18964
rect 52552 18912 52604 18964
rect 53288 18912 53340 18964
rect 54116 18912 54168 18964
rect 58256 18955 58308 18964
rect 58256 18921 58265 18955
rect 58265 18921 58299 18955
rect 58299 18921 58308 18955
rect 58256 18912 58308 18921
rect 34704 18708 34756 18760
rect 34796 18708 34848 18760
rect 37096 18751 37148 18760
rect 37096 18717 37105 18751
rect 37105 18717 37139 18751
rect 37139 18717 37148 18751
rect 37096 18708 37148 18717
rect 39764 18708 39816 18760
rect 40500 18708 40552 18760
rect 41236 18708 41288 18760
rect 45008 18751 45060 18760
rect 45008 18717 45017 18751
rect 45017 18717 45051 18751
rect 45051 18717 45060 18751
rect 45008 18708 45060 18717
rect 48964 18751 49016 18760
rect 48964 18717 48973 18751
rect 48973 18717 49007 18751
rect 49007 18717 49016 18751
rect 48964 18708 49016 18717
rect 49056 18708 49108 18760
rect 30840 18640 30892 18692
rect 31392 18640 31444 18692
rect 32128 18683 32180 18692
rect 32128 18649 32137 18683
rect 32137 18649 32171 18683
rect 32171 18649 32180 18683
rect 32128 18640 32180 18649
rect 38200 18683 38252 18692
rect 38200 18649 38209 18683
rect 38209 18649 38243 18683
rect 38243 18649 38252 18683
rect 38200 18640 38252 18649
rect 38292 18640 38344 18692
rect 39580 18640 39632 18692
rect 44088 18640 44140 18692
rect 47860 18640 47912 18692
rect 48320 18640 48372 18692
rect 49424 18640 49476 18692
rect 49608 18844 49660 18896
rect 50344 18751 50396 18760
rect 50344 18717 50353 18751
rect 50353 18717 50387 18751
rect 50387 18717 50396 18751
rect 50344 18708 50396 18717
rect 53840 18776 53892 18828
rect 51540 18708 51592 18760
rect 51816 18751 51868 18760
rect 51816 18717 51825 18751
rect 51825 18717 51859 18751
rect 51859 18717 51868 18751
rect 51816 18708 51868 18717
rect 52092 18751 52144 18760
rect 52092 18717 52101 18751
rect 52101 18717 52135 18751
rect 52135 18717 52144 18751
rect 52092 18708 52144 18717
rect 56876 18751 56928 18760
rect 56876 18717 56885 18751
rect 56885 18717 56919 18751
rect 56919 18717 56928 18751
rect 56876 18708 56928 18717
rect 57428 18708 57480 18760
rect 51080 18640 51132 18692
rect 31116 18572 31168 18624
rect 36820 18615 36872 18624
rect 36820 18581 36829 18615
rect 36829 18581 36863 18615
rect 36863 18581 36872 18615
rect 36820 18572 36872 18581
rect 37096 18572 37148 18624
rect 40868 18572 40920 18624
rect 48964 18572 49016 18624
rect 4874 18470 4926 18522
rect 4938 18470 4990 18522
rect 5002 18470 5054 18522
rect 5066 18470 5118 18522
rect 5130 18470 5182 18522
rect 35594 18470 35646 18522
rect 35658 18470 35710 18522
rect 35722 18470 35774 18522
rect 35786 18470 35838 18522
rect 35850 18470 35902 18522
rect 19892 18368 19944 18420
rect 21824 18368 21876 18420
rect 16580 18232 16632 18284
rect 18144 18232 18196 18284
rect 19616 18232 19668 18284
rect 17316 18164 17368 18216
rect 20260 18275 20312 18284
rect 20260 18241 20269 18275
rect 20269 18241 20303 18275
rect 20303 18241 20312 18275
rect 20260 18232 20312 18241
rect 20536 18275 20588 18284
rect 20536 18241 20545 18275
rect 20545 18241 20579 18275
rect 20579 18241 20588 18275
rect 20536 18232 20588 18241
rect 23020 18368 23072 18420
rect 23112 18368 23164 18420
rect 24676 18368 24728 18420
rect 24952 18411 25004 18420
rect 24952 18377 24961 18411
rect 24961 18377 24995 18411
rect 24995 18377 25004 18411
rect 24952 18368 25004 18377
rect 24768 18300 24820 18352
rect 28908 18368 28960 18420
rect 26516 18300 26568 18352
rect 20628 18164 20680 18216
rect 22376 18232 22428 18284
rect 22468 18275 22520 18284
rect 22468 18241 22477 18275
rect 22477 18241 22511 18275
rect 22511 18241 22520 18275
rect 22468 18232 22520 18241
rect 23296 18164 23348 18216
rect 23572 18275 23624 18284
rect 23572 18241 23581 18275
rect 23581 18241 23615 18275
rect 23615 18241 23624 18275
rect 23572 18232 23624 18241
rect 23848 18232 23900 18284
rect 25136 18232 25188 18284
rect 27988 18275 28040 18284
rect 27988 18241 27997 18275
rect 27997 18241 28031 18275
rect 28031 18241 28040 18275
rect 27988 18232 28040 18241
rect 28172 18275 28224 18284
rect 28172 18241 28181 18275
rect 28181 18241 28215 18275
rect 28215 18241 28224 18275
rect 28172 18232 28224 18241
rect 28264 18275 28316 18284
rect 28264 18241 28273 18275
rect 28273 18241 28307 18275
rect 28307 18241 28316 18275
rect 28264 18232 28316 18241
rect 29368 18300 29420 18352
rect 30196 18232 30248 18284
rect 25044 18207 25096 18216
rect 25044 18173 25053 18207
rect 25053 18173 25087 18207
rect 25087 18173 25096 18207
rect 25044 18164 25096 18173
rect 26516 18207 26568 18216
rect 26516 18173 26525 18207
rect 26525 18173 26559 18207
rect 26559 18173 26568 18207
rect 26516 18164 26568 18173
rect 26976 18164 27028 18216
rect 30104 18164 30156 18216
rect 30564 18275 30616 18284
rect 30564 18241 30573 18275
rect 30573 18241 30607 18275
rect 30607 18241 30616 18275
rect 30564 18232 30616 18241
rect 16672 18096 16724 18148
rect 22100 18096 22152 18148
rect 24584 18096 24636 18148
rect 29460 18096 29512 18148
rect 22376 18028 22428 18080
rect 23572 18028 23624 18080
rect 26056 18028 26108 18080
rect 30748 18275 30800 18284
rect 30748 18241 30762 18275
rect 30762 18241 30796 18275
rect 30796 18241 30800 18275
rect 32128 18411 32180 18420
rect 32128 18377 32137 18411
rect 32137 18377 32171 18411
rect 32171 18377 32180 18411
rect 32128 18368 32180 18377
rect 37096 18411 37148 18420
rect 37096 18377 37105 18411
rect 37105 18377 37139 18411
rect 37139 18377 37148 18411
rect 37096 18368 37148 18377
rect 37740 18368 37792 18420
rect 38016 18368 38068 18420
rect 40040 18368 40092 18420
rect 40132 18368 40184 18420
rect 37372 18300 37424 18352
rect 30748 18232 30800 18241
rect 32496 18275 32548 18284
rect 32496 18241 32505 18275
rect 32505 18241 32539 18275
rect 32539 18241 32548 18275
rect 32496 18232 32548 18241
rect 34060 18232 34112 18284
rect 37740 18275 37792 18284
rect 37740 18241 37749 18275
rect 37749 18241 37783 18275
rect 37783 18241 37792 18275
rect 37740 18232 37792 18241
rect 31116 18207 31168 18216
rect 31116 18173 31125 18207
rect 31125 18173 31159 18207
rect 31159 18173 31168 18207
rect 31116 18164 31168 18173
rect 33508 18164 33560 18216
rect 35992 18164 36044 18216
rect 31484 18096 31536 18148
rect 32312 18096 32364 18148
rect 38200 18300 38252 18352
rect 40960 18368 41012 18420
rect 43352 18368 43404 18420
rect 45468 18368 45520 18420
rect 56968 18368 57020 18420
rect 38568 18275 38620 18284
rect 38568 18241 38577 18275
rect 38577 18241 38611 18275
rect 38611 18241 38620 18275
rect 38568 18232 38620 18241
rect 38660 18275 38712 18284
rect 38660 18241 38669 18275
rect 38669 18241 38703 18275
rect 38703 18241 38712 18275
rect 38660 18232 38712 18241
rect 38936 18232 38988 18284
rect 39212 18275 39264 18284
rect 39212 18241 39221 18275
rect 39221 18241 39255 18275
rect 39255 18241 39264 18275
rect 39212 18232 39264 18241
rect 38844 18164 38896 18216
rect 39580 18275 39632 18284
rect 39580 18241 39589 18275
rect 39589 18241 39623 18275
rect 39623 18241 39632 18275
rect 39580 18232 39632 18241
rect 39672 18275 39724 18284
rect 39672 18241 39681 18275
rect 39681 18241 39715 18275
rect 39715 18241 39724 18275
rect 39672 18232 39724 18241
rect 39764 18275 39816 18284
rect 39764 18241 39774 18275
rect 39774 18241 39808 18275
rect 39808 18241 39816 18275
rect 39764 18232 39816 18241
rect 38660 18096 38712 18148
rect 39488 18207 39540 18216
rect 39488 18173 39497 18207
rect 39497 18173 39531 18207
rect 39531 18173 39540 18207
rect 39488 18164 39540 18173
rect 40132 18275 40184 18284
rect 40132 18241 40146 18275
rect 40146 18241 40180 18275
rect 40180 18241 40184 18275
rect 40132 18232 40184 18241
rect 40316 18232 40368 18284
rect 40500 18232 40552 18284
rect 40868 18275 40920 18284
rect 40868 18241 40877 18275
rect 40877 18241 40911 18275
rect 40911 18241 40920 18275
rect 40868 18232 40920 18241
rect 40960 18275 41012 18284
rect 40960 18241 40969 18275
rect 40969 18241 41003 18275
rect 41003 18241 41012 18275
rect 40960 18232 41012 18241
rect 50528 18300 50580 18352
rect 51264 18300 51316 18352
rect 40224 18164 40276 18216
rect 41604 18275 41656 18284
rect 41604 18241 41613 18275
rect 41613 18241 41647 18275
rect 41647 18241 41656 18275
rect 41604 18232 41656 18241
rect 46756 18232 46808 18284
rect 49976 18275 50028 18284
rect 49976 18241 49985 18275
rect 49985 18241 50019 18275
rect 50019 18241 50028 18275
rect 49976 18232 50028 18241
rect 50252 18275 50304 18284
rect 50252 18241 50261 18275
rect 50261 18241 50295 18275
rect 50295 18241 50304 18275
rect 50252 18232 50304 18241
rect 40684 18096 40736 18148
rect 31116 18028 31168 18080
rect 32496 18028 32548 18080
rect 37372 18028 37424 18080
rect 38292 18028 38344 18080
rect 38752 18028 38804 18080
rect 42984 18164 43036 18216
rect 49056 18164 49108 18216
rect 50436 18232 50488 18284
rect 50620 18232 50672 18284
rect 40960 18028 41012 18080
rect 41328 18071 41380 18080
rect 41328 18037 41337 18071
rect 41337 18037 41371 18071
rect 41371 18037 41380 18071
rect 41328 18028 41380 18037
rect 41512 18028 41564 18080
rect 50896 18028 50948 18080
rect 52736 18071 52788 18080
rect 52736 18037 52745 18071
rect 52745 18037 52779 18071
rect 52779 18037 52788 18071
rect 52736 18028 52788 18037
rect 52828 18028 52880 18080
rect 53012 18275 53064 18284
rect 53012 18241 53021 18275
rect 53021 18241 53055 18275
rect 53055 18241 53064 18275
rect 53012 18232 53064 18241
rect 56784 18275 56836 18284
rect 56784 18241 56793 18275
rect 56793 18241 56827 18275
rect 56827 18241 56836 18275
rect 56784 18232 56836 18241
rect 56968 18275 57020 18284
rect 56968 18241 56977 18275
rect 56977 18241 57011 18275
rect 57011 18241 57020 18275
rect 56968 18232 57020 18241
rect 58164 18232 58216 18284
rect 54208 18164 54260 18216
rect 53840 18096 53892 18148
rect 54760 18096 54812 18148
rect 54484 18028 54536 18080
rect 56048 18071 56100 18080
rect 56048 18037 56057 18071
rect 56057 18037 56091 18071
rect 56091 18037 56100 18071
rect 56048 18028 56100 18037
rect 56416 18028 56468 18080
rect 57428 18071 57480 18080
rect 57428 18037 57437 18071
rect 57437 18037 57471 18071
rect 57471 18037 57480 18071
rect 57428 18028 57480 18037
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 22100 17824 22152 17876
rect 23112 17824 23164 17876
rect 24584 17824 24636 17876
rect 25780 17867 25832 17876
rect 25780 17833 25789 17867
rect 25789 17833 25823 17867
rect 25823 17833 25832 17867
rect 25780 17824 25832 17833
rect 26516 17824 26568 17876
rect 34704 17824 34756 17876
rect 26148 17756 26200 17808
rect 35992 17867 36044 17876
rect 35992 17833 36001 17867
rect 36001 17833 36035 17867
rect 36035 17833 36044 17867
rect 35992 17824 36044 17833
rect 38016 17824 38068 17876
rect 38476 17824 38528 17876
rect 38660 17867 38712 17876
rect 38660 17833 38669 17867
rect 38669 17833 38703 17867
rect 38703 17833 38712 17867
rect 38660 17824 38712 17833
rect 39948 17867 40000 17876
rect 39948 17833 39957 17867
rect 39957 17833 39991 17867
rect 39991 17833 40000 17867
rect 39948 17824 40000 17833
rect 40684 17867 40736 17876
rect 40684 17833 40693 17867
rect 40693 17833 40727 17867
rect 40727 17833 40736 17867
rect 40684 17824 40736 17833
rect 36176 17756 36228 17808
rect 16672 17663 16724 17672
rect 16672 17629 16681 17663
rect 16681 17629 16715 17663
rect 16715 17629 16724 17663
rect 16672 17620 16724 17629
rect 26608 17688 26660 17740
rect 30380 17688 30432 17740
rect 31576 17688 31628 17740
rect 26332 17663 26384 17672
rect 26332 17629 26341 17663
rect 26341 17629 26375 17663
rect 26375 17629 26384 17663
rect 26332 17620 26384 17629
rect 26424 17663 26476 17672
rect 26424 17629 26433 17663
rect 26433 17629 26467 17663
rect 26467 17629 26476 17663
rect 26424 17620 26476 17629
rect 30288 17663 30340 17672
rect 30288 17629 30297 17663
rect 30297 17629 30331 17663
rect 30331 17629 30340 17663
rect 30288 17620 30340 17629
rect 34520 17620 34572 17672
rect 34888 17663 34940 17672
rect 34888 17629 34897 17663
rect 34897 17629 34931 17663
rect 34931 17629 34940 17663
rect 34888 17620 34940 17629
rect 35072 17620 35124 17672
rect 35256 17663 35308 17672
rect 35256 17629 35281 17663
rect 35281 17629 35308 17663
rect 35256 17620 35308 17629
rect 36176 17663 36228 17672
rect 36176 17629 36185 17663
rect 36185 17629 36219 17663
rect 36219 17629 36228 17663
rect 36176 17620 36228 17629
rect 36544 17663 36596 17672
rect 36544 17629 36553 17663
rect 36553 17629 36587 17663
rect 36587 17629 36596 17663
rect 37096 17756 37148 17808
rect 38108 17756 38160 17808
rect 39212 17756 39264 17808
rect 36544 17620 36596 17629
rect 36820 17663 36872 17672
rect 36820 17629 36829 17663
rect 36829 17629 36863 17663
rect 36863 17629 36872 17663
rect 36820 17620 36872 17629
rect 37740 17688 37792 17740
rect 40040 17731 40092 17740
rect 40040 17697 40049 17731
rect 40049 17697 40083 17731
rect 40083 17697 40092 17731
rect 40040 17688 40092 17697
rect 25044 17552 25096 17604
rect 31024 17595 31076 17604
rect 31024 17561 31033 17595
rect 31033 17561 31067 17595
rect 31067 17561 31076 17595
rect 31024 17552 31076 17561
rect 31484 17552 31536 17604
rect 30472 17527 30524 17536
rect 30472 17493 30481 17527
rect 30481 17493 30515 17527
rect 30515 17493 30524 17527
rect 30472 17484 30524 17493
rect 30748 17484 30800 17536
rect 31668 17484 31720 17536
rect 32312 17484 32364 17536
rect 33784 17484 33836 17536
rect 35256 17484 35308 17536
rect 35992 17552 36044 17604
rect 38752 17620 38804 17672
rect 37004 17595 37056 17604
rect 37004 17561 37013 17595
rect 37013 17561 37047 17595
rect 37047 17561 37056 17595
rect 37004 17552 37056 17561
rect 37096 17552 37148 17604
rect 37556 17552 37608 17604
rect 40592 17620 40644 17672
rect 43812 17867 43864 17876
rect 43812 17833 43821 17867
rect 43821 17833 43855 17867
rect 43855 17833 43864 17867
rect 43812 17824 43864 17833
rect 42616 17756 42668 17808
rect 47492 17824 47544 17876
rect 48596 17824 48648 17876
rect 49332 17824 49384 17876
rect 49516 17867 49568 17876
rect 49516 17833 49525 17867
rect 49525 17833 49559 17867
rect 49559 17833 49568 17867
rect 49516 17824 49568 17833
rect 56600 17824 56652 17876
rect 58164 17824 58216 17876
rect 47952 17756 48004 17808
rect 49700 17756 49752 17808
rect 41512 17731 41564 17740
rect 41512 17697 41521 17731
rect 41521 17697 41555 17731
rect 41555 17697 41564 17731
rect 41512 17688 41564 17697
rect 42984 17731 43036 17740
rect 42984 17697 42993 17731
rect 42993 17697 43027 17731
rect 43027 17697 43036 17731
rect 42984 17688 43036 17697
rect 41236 17663 41288 17672
rect 41236 17629 41245 17663
rect 41245 17629 41279 17663
rect 41279 17629 41288 17663
rect 41236 17620 41288 17629
rect 43076 17663 43128 17672
rect 43076 17629 43085 17663
rect 43085 17629 43119 17663
rect 43119 17629 43128 17663
rect 43076 17620 43128 17629
rect 45008 17688 45060 17740
rect 43352 17663 43404 17672
rect 43352 17629 43361 17663
rect 43361 17629 43395 17663
rect 43395 17629 43404 17663
rect 43352 17620 43404 17629
rect 43444 17663 43496 17672
rect 43444 17629 43453 17663
rect 43453 17629 43487 17663
rect 43487 17629 43496 17663
rect 43444 17620 43496 17629
rect 43812 17620 43864 17672
rect 47860 17620 47912 17672
rect 48964 17688 49016 17740
rect 49056 17620 49108 17672
rect 49976 17688 50028 17740
rect 54484 17756 54536 17808
rect 55956 17756 56008 17808
rect 53932 17688 53984 17740
rect 54760 17731 54812 17740
rect 54760 17697 54769 17731
rect 54769 17697 54803 17731
rect 54803 17697 54812 17731
rect 54760 17688 54812 17697
rect 55220 17688 55272 17740
rect 49700 17663 49752 17672
rect 49700 17629 49709 17663
rect 49709 17629 49743 17663
rect 49743 17629 49752 17663
rect 49700 17620 49752 17629
rect 53840 17620 53892 17672
rect 54484 17663 54536 17672
rect 54484 17629 54493 17663
rect 54493 17629 54527 17663
rect 54527 17629 54536 17663
rect 54484 17620 54536 17629
rect 54576 17663 54628 17672
rect 54576 17629 54585 17663
rect 54585 17629 54619 17663
rect 54619 17629 54628 17663
rect 54576 17620 54628 17629
rect 39856 17595 39908 17604
rect 39856 17561 39865 17595
rect 39865 17561 39899 17595
rect 39899 17561 39908 17595
rect 39856 17552 39908 17561
rect 36452 17484 36504 17536
rect 40132 17484 40184 17536
rect 44088 17552 44140 17604
rect 46756 17595 46808 17604
rect 46756 17561 46765 17595
rect 46765 17561 46799 17595
rect 46799 17561 46808 17595
rect 46756 17552 46808 17561
rect 48412 17552 48464 17604
rect 50620 17552 50672 17604
rect 51356 17552 51408 17604
rect 52736 17595 52788 17604
rect 52736 17561 52745 17595
rect 52745 17561 52779 17595
rect 52779 17561 52788 17595
rect 52736 17552 52788 17561
rect 41144 17527 41196 17536
rect 41144 17493 41153 17527
rect 41153 17493 41187 17527
rect 41187 17493 41196 17527
rect 41144 17484 41196 17493
rect 41328 17484 41380 17536
rect 47584 17484 47636 17536
rect 48228 17484 48280 17536
rect 48320 17527 48372 17536
rect 48320 17493 48329 17527
rect 48329 17493 48363 17527
rect 48363 17493 48372 17527
rect 48320 17484 48372 17493
rect 52368 17527 52420 17536
rect 52368 17493 52377 17527
rect 52377 17493 52411 17527
rect 52411 17493 52420 17527
rect 52368 17484 52420 17493
rect 53104 17484 53156 17536
rect 55772 17552 55824 17604
rect 54208 17527 54260 17536
rect 54208 17493 54217 17527
rect 54217 17493 54251 17527
rect 54251 17493 54260 17527
rect 54208 17484 54260 17493
rect 54392 17484 54444 17536
rect 55680 17527 55732 17536
rect 55680 17493 55689 17527
rect 55689 17493 55723 17527
rect 55723 17493 55732 17527
rect 56416 17663 56468 17672
rect 56416 17629 56425 17663
rect 56425 17629 56459 17663
rect 56459 17629 56468 17663
rect 56416 17620 56468 17629
rect 56600 17620 56652 17672
rect 56876 17663 56928 17672
rect 56876 17629 56885 17663
rect 56885 17629 56919 17663
rect 56919 17629 56928 17663
rect 56876 17620 56928 17629
rect 57428 17620 57480 17672
rect 56692 17552 56744 17604
rect 55680 17484 55732 17493
rect 56232 17527 56284 17536
rect 56232 17493 56241 17527
rect 56241 17493 56275 17527
rect 56275 17493 56284 17527
rect 56232 17484 56284 17493
rect 4874 17382 4926 17434
rect 4938 17382 4990 17434
rect 5002 17382 5054 17434
rect 5066 17382 5118 17434
rect 5130 17382 5182 17434
rect 35594 17382 35646 17434
rect 35658 17382 35710 17434
rect 35722 17382 35774 17434
rect 35786 17382 35838 17434
rect 35850 17382 35902 17434
rect 16764 17280 16816 17332
rect 17960 17212 18012 17264
rect 21640 17212 21692 17264
rect 22284 17212 22336 17264
rect 24676 17255 24728 17264
rect 24676 17221 24685 17255
rect 24685 17221 24719 17255
rect 24719 17221 24728 17255
rect 24676 17212 24728 17221
rect 16672 17076 16724 17128
rect 19340 17119 19392 17128
rect 19340 17085 19349 17119
rect 19349 17085 19383 17119
rect 19383 17085 19392 17119
rect 19340 17076 19392 17085
rect 19800 17187 19852 17196
rect 19800 17153 19809 17187
rect 19809 17153 19843 17187
rect 19843 17153 19852 17187
rect 19800 17144 19852 17153
rect 19708 17076 19760 17128
rect 20352 17144 20404 17196
rect 23204 17144 23256 17196
rect 24032 17187 24084 17196
rect 24032 17153 24041 17187
rect 24041 17153 24075 17187
rect 24075 17153 24084 17187
rect 24032 17144 24084 17153
rect 20168 17076 20220 17128
rect 23020 17076 23072 17128
rect 24584 17144 24636 17196
rect 24952 17144 25004 17196
rect 26792 17280 26844 17332
rect 29000 17280 29052 17332
rect 32220 17323 32272 17332
rect 26240 17212 26292 17264
rect 32220 17289 32229 17323
rect 32229 17289 32263 17323
rect 32263 17289 32272 17323
rect 32220 17280 32272 17289
rect 32404 17323 32456 17332
rect 32404 17289 32413 17323
rect 32413 17289 32447 17323
rect 32447 17289 32456 17323
rect 32404 17280 32456 17289
rect 32496 17323 32548 17332
rect 32496 17289 32505 17323
rect 32505 17289 32539 17323
rect 32539 17289 32548 17323
rect 32496 17280 32548 17289
rect 25228 17119 25280 17128
rect 25228 17085 25237 17119
rect 25237 17085 25271 17119
rect 25271 17085 25280 17119
rect 25228 17076 25280 17085
rect 19248 16983 19300 16992
rect 19248 16949 19257 16983
rect 19257 16949 19291 16983
rect 19291 16949 19300 16983
rect 19248 16940 19300 16949
rect 22744 16940 22796 16992
rect 23112 16940 23164 16992
rect 23664 17008 23716 17060
rect 27896 17144 27948 17196
rect 29828 17144 29880 17196
rect 29920 17187 29972 17196
rect 29920 17153 29929 17187
rect 29929 17153 29963 17187
rect 29963 17153 29972 17187
rect 29920 17144 29972 17153
rect 26332 17119 26384 17128
rect 26332 17085 26341 17119
rect 26341 17085 26375 17119
rect 26375 17085 26384 17119
rect 26332 17076 26384 17085
rect 26424 17076 26476 17128
rect 27804 17119 27856 17128
rect 27804 17085 27813 17119
rect 27813 17085 27847 17119
rect 27847 17085 27856 17119
rect 27804 17076 27856 17085
rect 29368 17119 29420 17128
rect 29368 17085 29377 17119
rect 29377 17085 29411 17119
rect 29411 17085 29420 17119
rect 30656 17187 30708 17196
rect 30656 17153 30665 17187
rect 30665 17153 30699 17187
rect 30699 17153 30708 17187
rect 30656 17144 30708 17153
rect 32128 17212 32180 17264
rect 31024 17187 31076 17196
rect 31024 17153 31033 17187
rect 31033 17153 31067 17187
rect 31067 17153 31076 17187
rect 31024 17144 31076 17153
rect 31116 17187 31168 17196
rect 31116 17153 31125 17187
rect 31125 17153 31159 17187
rect 31159 17153 31168 17187
rect 31116 17144 31168 17153
rect 31208 17187 31260 17196
rect 31208 17153 31218 17187
rect 31218 17153 31252 17187
rect 31252 17153 31260 17187
rect 31208 17144 31260 17153
rect 31392 17187 31444 17196
rect 31392 17153 31401 17187
rect 31401 17153 31435 17187
rect 31435 17153 31444 17187
rect 31392 17144 31444 17153
rect 31668 17144 31720 17196
rect 33784 17255 33836 17264
rect 33784 17221 33793 17255
rect 33793 17221 33827 17255
rect 33827 17221 33836 17255
rect 33784 17212 33836 17221
rect 34244 17212 34296 17264
rect 35164 17280 35216 17332
rect 36084 17280 36136 17332
rect 36820 17280 36872 17332
rect 37188 17280 37240 17332
rect 38108 17323 38160 17332
rect 38108 17289 38117 17323
rect 38117 17289 38151 17323
rect 38151 17289 38160 17323
rect 38108 17280 38160 17289
rect 38936 17280 38988 17332
rect 39304 17280 39356 17332
rect 39764 17323 39816 17332
rect 39764 17289 39773 17323
rect 39773 17289 39807 17323
rect 39807 17289 39816 17323
rect 39764 17280 39816 17289
rect 40408 17280 40460 17332
rect 40592 17323 40644 17332
rect 40592 17289 40601 17323
rect 40601 17289 40635 17323
rect 40635 17289 40644 17323
rect 40592 17280 40644 17289
rect 40684 17280 40736 17332
rect 41972 17280 42024 17332
rect 43076 17280 43128 17332
rect 41144 17255 41196 17264
rect 41144 17221 41153 17255
rect 41153 17221 41187 17255
rect 41187 17221 41196 17255
rect 41144 17212 41196 17221
rect 42616 17255 42668 17264
rect 42616 17221 42625 17255
rect 42625 17221 42659 17255
rect 42659 17221 42668 17255
rect 42616 17212 42668 17221
rect 42708 17255 42760 17264
rect 42708 17221 42717 17255
rect 42717 17221 42751 17255
rect 42751 17221 42760 17255
rect 42708 17212 42760 17221
rect 33508 17187 33560 17196
rect 33508 17153 33517 17187
rect 33517 17153 33551 17187
rect 33551 17153 33560 17187
rect 33508 17144 33560 17153
rect 29368 17076 29420 17085
rect 30748 17076 30800 17128
rect 34520 17076 34572 17128
rect 35716 17144 35768 17196
rect 35900 17187 35952 17196
rect 35900 17153 35909 17187
rect 35909 17153 35943 17187
rect 35943 17153 35952 17187
rect 35900 17144 35952 17153
rect 35256 17119 35308 17128
rect 35256 17085 35265 17119
rect 35265 17085 35299 17119
rect 35299 17085 35308 17119
rect 35256 17076 35308 17085
rect 35532 17076 35584 17128
rect 36084 17187 36136 17196
rect 36084 17153 36093 17187
rect 36093 17153 36127 17187
rect 36127 17153 36136 17187
rect 36084 17144 36136 17153
rect 36544 17144 36596 17196
rect 37280 17076 37332 17128
rect 31208 17008 31260 17060
rect 24216 16940 24268 16992
rect 24400 16940 24452 16992
rect 25412 16940 25464 16992
rect 25872 16983 25924 16992
rect 25872 16949 25881 16983
rect 25881 16949 25915 16983
rect 25915 16949 25924 16983
rect 25872 16940 25924 16949
rect 27252 16940 27304 16992
rect 29460 16983 29512 16992
rect 29460 16949 29469 16983
rect 29469 16949 29503 16983
rect 29503 16949 29512 16983
rect 29460 16940 29512 16949
rect 29644 16940 29696 16992
rect 30288 16940 30340 16992
rect 31760 16983 31812 16992
rect 31760 16949 31769 16983
rect 31769 16949 31803 16983
rect 31803 16949 31812 16983
rect 31760 16940 31812 16949
rect 31852 16983 31904 16992
rect 31852 16949 31861 16983
rect 31861 16949 31895 16983
rect 31895 16949 31904 16983
rect 31852 16940 31904 16949
rect 34888 17008 34940 17060
rect 36176 17008 36228 17060
rect 36544 17008 36596 17060
rect 38752 17187 38804 17196
rect 38752 17153 38761 17187
rect 38761 17153 38795 17187
rect 38795 17153 38804 17187
rect 38752 17144 38804 17153
rect 39764 17144 39816 17196
rect 39948 17187 40000 17196
rect 39948 17153 39957 17187
rect 39957 17153 39991 17187
rect 39991 17153 40000 17187
rect 39948 17144 40000 17153
rect 40316 17187 40368 17196
rect 40316 17153 40325 17187
rect 40325 17153 40359 17187
rect 40359 17153 40368 17187
rect 40316 17144 40368 17153
rect 40868 17187 40920 17196
rect 40868 17153 40877 17187
rect 40877 17153 40911 17187
rect 40911 17153 40920 17187
rect 40868 17144 40920 17153
rect 41052 17144 41104 17196
rect 40592 17076 40644 17128
rect 42340 17144 42392 17196
rect 43904 17280 43956 17332
rect 44088 17280 44140 17332
rect 44548 17280 44600 17332
rect 46756 17280 46808 17332
rect 49056 17280 49108 17332
rect 46572 17212 46624 17264
rect 46020 17187 46072 17196
rect 46020 17153 46029 17187
rect 46029 17153 46063 17187
rect 46063 17153 46072 17187
rect 46020 17144 46072 17153
rect 46204 17187 46256 17196
rect 46204 17153 46211 17187
rect 46211 17153 46256 17187
rect 46204 17144 46256 17153
rect 46296 17187 46348 17196
rect 46296 17153 46305 17187
rect 46305 17153 46339 17187
rect 46339 17153 46348 17187
rect 46296 17144 46348 17153
rect 39396 17008 39448 17060
rect 35900 16940 35952 16992
rect 36636 16983 36688 16992
rect 36636 16949 36645 16983
rect 36645 16949 36679 16983
rect 36679 16949 36688 16983
rect 36636 16940 36688 16949
rect 38476 16983 38528 16992
rect 38476 16949 38485 16983
rect 38485 16949 38519 16983
rect 38519 16949 38528 16983
rect 38476 16940 38528 16949
rect 38660 16940 38712 16992
rect 42984 17076 43036 17128
rect 43444 17119 43496 17128
rect 43444 17085 43453 17119
rect 43453 17085 43487 17119
rect 43487 17085 43496 17119
rect 43444 17076 43496 17085
rect 43812 17076 43864 17128
rect 40868 17008 40920 17060
rect 41604 17008 41656 17060
rect 41788 17008 41840 17060
rect 42616 17008 42668 17060
rect 43536 16940 43588 16992
rect 46480 17187 46532 17196
rect 48504 17212 48556 17264
rect 49516 17323 49568 17332
rect 49516 17289 49525 17323
rect 49525 17289 49559 17323
rect 49559 17289 49568 17323
rect 49516 17280 49568 17289
rect 49700 17323 49752 17332
rect 49700 17289 49709 17323
rect 49709 17289 49743 17323
rect 49743 17289 49752 17323
rect 49700 17280 49752 17289
rect 49792 17280 49844 17332
rect 50620 17323 50672 17332
rect 50620 17289 50629 17323
rect 50629 17289 50663 17323
rect 50663 17289 50672 17323
rect 50620 17280 50672 17289
rect 53012 17280 53064 17332
rect 53472 17280 53524 17332
rect 46480 17153 46494 17187
rect 46494 17153 46528 17187
rect 46528 17153 46532 17187
rect 46480 17144 46532 17153
rect 48320 17144 48372 17196
rect 48872 17187 48924 17196
rect 48872 17153 48881 17187
rect 48881 17153 48915 17187
rect 48915 17153 48924 17187
rect 48872 17144 48924 17153
rect 49056 17187 49108 17196
rect 49056 17153 49063 17187
rect 49063 17153 49108 17187
rect 49056 17144 49108 17153
rect 48780 17076 48832 17128
rect 49332 17187 49384 17196
rect 49332 17153 49346 17187
rect 49346 17153 49380 17187
rect 49380 17153 49384 17187
rect 50068 17255 50120 17264
rect 50068 17221 50077 17255
rect 50077 17221 50111 17255
rect 50111 17221 50120 17255
rect 50068 17212 50120 17221
rect 53380 17212 53432 17264
rect 54576 17280 54628 17332
rect 55772 17280 55824 17332
rect 49332 17144 49384 17153
rect 50252 17187 50304 17196
rect 49792 17076 49844 17128
rect 50252 17153 50260 17187
rect 50260 17153 50294 17187
rect 50294 17153 50304 17187
rect 50252 17144 50304 17153
rect 50344 17187 50396 17196
rect 50344 17153 50353 17187
rect 50353 17153 50387 17187
rect 50387 17153 50396 17187
rect 50344 17144 50396 17153
rect 50804 17187 50856 17196
rect 50804 17153 50813 17187
rect 50813 17153 50847 17187
rect 50847 17153 50856 17187
rect 50804 17144 50856 17153
rect 50896 17187 50948 17196
rect 50896 17153 50905 17187
rect 50905 17153 50939 17187
rect 50939 17153 50948 17187
rect 50896 17144 50948 17153
rect 51632 17144 51684 17196
rect 52368 17144 52420 17196
rect 52920 17187 52972 17196
rect 52920 17153 52929 17187
rect 52929 17153 52963 17187
rect 52963 17153 52972 17187
rect 52920 17144 52972 17153
rect 53012 17187 53064 17196
rect 53012 17153 53021 17187
rect 53021 17153 53055 17187
rect 53055 17153 53064 17187
rect 53012 17144 53064 17153
rect 53196 17144 53248 17196
rect 54392 17255 54444 17264
rect 54392 17221 54401 17255
rect 54401 17221 54435 17255
rect 54435 17221 54444 17255
rect 54392 17212 54444 17221
rect 54852 17212 54904 17264
rect 53748 17187 53800 17196
rect 53748 17153 53749 17187
rect 53749 17153 53783 17187
rect 53783 17153 53800 17187
rect 53748 17144 53800 17153
rect 51540 17008 51592 17060
rect 51816 17008 51868 17060
rect 53196 17008 53248 17060
rect 53564 17008 53616 17060
rect 53932 17076 53984 17128
rect 56876 17280 56928 17332
rect 56232 17255 56284 17264
rect 56232 17221 56241 17255
rect 56241 17221 56275 17255
rect 56275 17221 56284 17255
rect 56232 17212 56284 17221
rect 56784 17212 56836 17264
rect 56692 17076 56744 17128
rect 57520 17076 57572 17128
rect 45284 16983 45336 16992
rect 45284 16949 45293 16983
rect 45293 16949 45327 16983
rect 45327 16949 45336 16983
rect 45284 16940 45336 16949
rect 47492 16940 47544 16992
rect 48320 16983 48372 16992
rect 48320 16949 48329 16983
rect 48329 16949 48363 16983
rect 48363 16949 48372 16983
rect 48320 16940 48372 16949
rect 48504 16983 48556 16992
rect 48504 16949 48513 16983
rect 48513 16949 48547 16983
rect 48547 16949 48556 16983
rect 48504 16940 48556 16949
rect 51080 16983 51132 16992
rect 51080 16949 51089 16983
rect 51089 16949 51123 16983
rect 51123 16949 51132 16983
rect 51080 16940 51132 16949
rect 51264 16940 51316 16992
rect 52920 16940 52972 16992
rect 53472 16940 53524 16992
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 22744 16736 22796 16788
rect 23020 16736 23072 16788
rect 25044 16736 25096 16788
rect 16672 16643 16724 16652
rect 16672 16609 16681 16643
rect 16681 16609 16715 16643
rect 16715 16609 16724 16643
rect 16672 16600 16724 16609
rect 19524 16600 19576 16652
rect 18880 16575 18932 16584
rect 18880 16541 18889 16575
rect 18889 16541 18923 16575
rect 18923 16541 18932 16575
rect 18880 16532 18932 16541
rect 18972 16575 19024 16584
rect 18972 16541 18981 16575
rect 18981 16541 19015 16575
rect 19015 16541 19024 16575
rect 18972 16532 19024 16541
rect 19708 16532 19760 16584
rect 22192 16600 22244 16652
rect 24124 16600 24176 16652
rect 25320 16736 25372 16788
rect 25872 16779 25924 16788
rect 25872 16745 25881 16779
rect 25881 16745 25915 16779
rect 25915 16745 25924 16779
rect 25872 16736 25924 16745
rect 25964 16736 26016 16788
rect 26884 16736 26936 16788
rect 27804 16736 27856 16788
rect 25228 16668 25280 16720
rect 17960 16464 18012 16516
rect 19340 16464 19392 16516
rect 18972 16396 19024 16448
rect 19616 16507 19668 16516
rect 19616 16473 19625 16507
rect 19625 16473 19659 16507
rect 19659 16473 19668 16507
rect 19616 16464 19668 16473
rect 20352 16532 20404 16584
rect 21916 16532 21968 16584
rect 19984 16464 20036 16516
rect 20812 16507 20864 16516
rect 20812 16473 20821 16507
rect 20821 16473 20855 16507
rect 20855 16473 20864 16507
rect 20812 16464 20864 16473
rect 24400 16575 24452 16584
rect 24400 16541 24409 16575
rect 24409 16541 24443 16575
rect 24443 16541 24452 16575
rect 24400 16532 24452 16541
rect 24492 16575 24544 16584
rect 24492 16541 24502 16575
rect 24502 16541 24536 16575
rect 24536 16541 24544 16575
rect 24492 16532 24544 16541
rect 26424 16600 26476 16652
rect 25044 16532 25096 16584
rect 25320 16575 25372 16584
rect 25320 16541 25329 16575
rect 25329 16541 25363 16575
rect 25363 16541 25372 16575
rect 25320 16532 25372 16541
rect 24584 16464 24636 16516
rect 25688 16575 25740 16584
rect 25688 16541 25697 16575
rect 25697 16541 25731 16575
rect 25731 16541 25740 16575
rect 25688 16532 25740 16541
rect 25872 16532 25924 16584
rect 26240 16532 26292 16584
rect 26976 16643 27028 16652
rect 26976 16609 26985 16643
rect 26985 16609 27019 16643
rect 27019 16609 27028 16643
rect 26976 16600 27028 16609
rect 27252 16643 27304 16652
rect 27252 16609 27261 16643
rect 27261 16609 27295 16643
rect 27295 16609 27304 16643
rect 27252 16600 27304 16609
rect 29828 16736 29880 16788
rect 30656 16736 30708 16788
rect 30932 16736 30984 16788
rect 31024 16736 31076 16788
rect 34244 16736 34296 16788
rect 35808 16736 35860 16788
rect 22192 16396 22244 16448
rect 22376 16396 22428 16448
rect 23664 16396 23716 16448
rect 24400 16396 24452 16448
rect 25504 16507 25556 16516
rect 25504 16473 25513 16507
rect 25513 16473 25547 16507
rect 25547 16473 25556 16507
rect 25504 16464 25556 16473
rect 25412 16396 25464 16448
rect 25872 16396 25924 16448
rect 26792 16575 26844 16584
rect 26792 16541 26801 16575
rect 26801 16541 26835 16575
rect 26835 16541 26844 16575
rect 26792 16532 26844 16541
rect 26884 16396 26936 16448
rect 28356 16532 28408 16584
rect 28908 16532 28960 16584
rect 29000 16575 29052 16584
rect 29000 16541 29009 16575
rect 29009 16541 29043 16575
rect 29043 16541 29052 16575
rect 29000 16532 29052 16541
rect 29184 16575 29236 16584
rect 29184 16541 29193 16575
rect 29193 16541 29227 16575
rect 29227 16541 29236 16575
rect 29184 16532 29236 16541
rect 29368 16575 29420 16584
rect 29368 16541 29377 16575
rect 29377 16541 29411 16575
rect 29411 16541 29420 16575
rect 29368 16532 29420 16541
rect 29552 16575 29604 16584
rect 29552 16541 29561 16575
rect 29561 16541 29595 16575
rect 29595 16541 29604 16575
rect 29552 16532 29604 16541
rect 30564 16668 30616 16720
rect 31392 16668 31444 16720
rect 34060 16668 34112 16720
rect 29828 16575 29880 16584
rect 29828 16541 29837 16575
rect 29837 16541 29871 16575
rect 29871 16541 29880 16575
rect 29828 16532 29880 16541
rect 30472 16532 30524 16584
rect 30196 16464 30248 16516
rect 33508 16600 33560 16652
rect 34796 16600 34848 16652
rect 35256 16600 35308 16652
rect 35164 16575 35216 16584
rect 35164 16541 35173 16575
rect 35173 16541 35207 16575
rect 35207 16541 35216 16575
rect 35164 16532 35216 16541
rect 35440 16575 35492 16584
rect 35440 16541 35449 16575
rect 35449 16541 35483 16575
rect 35483 16541 35492 16575
rect 35440 16532 35492 16541
rect 35716 16575 35768 16584
rect 35716 16541 35725 16575
rect 35725 16541 35759 16575
rect 35759 16541 35768 16575
rect 35716 16532 35768 16541
rect 37096 16736 37148 16788
rect 37188 16779 37240 16788
rect 37188 16745 37197 16779
rect 37197 16745 37231 16779
rect 37231 16745 37240 16779
rect 37188 16736 37240 16745
rect 35992 16600 36044 16652
rect 29552 16396 29604 16448
rect 30104 16396 30156 16448
rect 30656 16396 30708 16448
rect 31484 16464 31536 16516
rect 31208 16439 31260 16448
rect 31208 16405 31217 16439
rect 31217 16405 31251 16439
rect 31251 16405 31260 16439
rect 31208 16396 31260 16405
rect 32772 16507 32824 16516
rect 32772 16473 32781 16507
rect 32781 16473 32815 16507
rect 32815 16473 32824 16507
rect 32772 16464 32824 16473
rect 35348 16464 35400 16516
rect 34888 16439 34940 16448
rect 34888 16405 34897 16439
rect 34897 16405 34931 16439
rect 34931 16405 34940 16439
rect 34888 16396 34940 16405
rect 35164 16396 35216 16448
rect 35992 16464 36044 16516
rect 36728 16668 36780 16720
rect 36820 16668 36872 16720
rect 36636 16532 36688 16584
rect 38660 16736 38712 16788
rect 39948 16736 40000 16788
rect 38476 16711 38528 16720
rect 38476 16677 38485 16711
rect 38485 16677 38519 16711
rect 38519 16677 38528 16711
rect 38476 16668 38528 16677
rect 41328 16736 41380 16788
rect 45376 16736 45428 16788
rect 46480 16736 46532 16788
rect 47860 16736 47912 16788
rect 48044 16736 48096 16788
rect 48320 16779 48372 16788
rect 48320 16745 48329 16779
rect 48329 16745 48363 16779
rect 48363 16745 48372 16779
rect 48320 16736 48372 16745
rect 48872 16736 48924 16788
rect 40132 16668 40184 16720
rect 40684 16668 40736 16720
rect 40776 16668 40828 16720
rect 41052 16668 41104 16720
rect 41144 16668 41196 16720
rect 37832 16532 37884 16584
rect 36544 16507 36596 16516
rect 36544 16473 36553 16507
rect 36553 16473 36587 16507
rect 36587 16473 36596 16507
rect 36544 16464 36596 16473
rect 36084 16396 36136 16448
rect 36728 16396 36780 16448
rect 37280 16507 37332 16516
rect 37280 16473 37289 16507
rect 37289 16473 37323 16507
rect 37323 16473 37332 16507
rect 37280 16464 37332 16473
rect 37464 16396 37516 16448
rect 38292 16507 38344 16516
rect 38292 16473 38301 16507
rect 38301 16473 38335 16507
rect 38335 16473 38344 16507
rect 38292 16464 38344 16473
rect 38384 16464 38436 16516
rect 38936 16575 38988 16584
rect 38936 16541 38945 16575
rect 38945 16541 38979 16575
rect 38979 16541 38988 16575
rect 38936 16532 38988 16541
rect 38752 16507 38804 16516
rect 38752 16473 38761 16507
rect 38761 16473 38795 16507
rect 38795 16473 38804 16507
rect 38752 16464 38804 16473
rect 38844 16507 38896 16516
rect 38844 16473 38853 16507
rect 38853 16473 38887 16507
rect 38887 16473 38896 16507
rect 38844 16464 38896 16473
rect 40040 16575 40092 16584
rect 40040 16541 40049 16575
rect 40049 16541 40083 16575
rect 40083 16541 40092 16575
rect 40040 16532 40092 16541
rect 40868 16600 40920 16652
rect 40960 16643 41012 16652
rect 40960 16609 40969 16643
rect 40969 16609 41003 16643
rect 41003 16609 41012 16643
rect 40960 16600 41012 16609
rect 41328 16600 41380 16652
rect 41512 16668 41564 16720
rect 43996 16668 44048 16720
rect 46848 16668 46900 16720
rect 48504 16668 48556 16720
rect 50068 16668 50120 16720
rect 40776 16575 40828 16584
rect 40776 16541 40785 16575
rect 40785 16541 40819 16575
rect 40819 16541 40828 16575
rect 40776 16532 40828 16541
rect 41788 16532 41840 16584
rect 42800 16575 42852 16584
rect 42800 16541 42809 16575
rect 42809 16541 42843 16575
rect 42843 16541 42852 16575
rect 42800 16532 42852 16541
rect 42984 16575 43036 16584
rect 42984 16541 42993 16575
rect 42993 16541 43027 16575
rect 43027 16541 43036 16575
rect 42984 16532 43036 16541
rect 43076 16575 43128 16584
rect 43076 16541 43085 16575
rect 43085 16541 43119 16575
rect 43119 16541 43128 16575
rect 43076 16532 43128 16541
rect 43168 16532 43220 16584
rect 38476 16396 38528 16448
rect 38660 16396 38712 16448
rect 40132 16507 40184 16516
rect 40132 16473 40141 16507
rect 40141 16473 40175 16507
rect 40175 16473 40184 16507
rect 40132 16464 40184 16473
rect 41880 16464 41932 16516
rect 43904 16532 43956 16584
rect 44180 16532 44232 16584
rect 46296 16600 46348 16652
rect 45284 16532 45336 16584
rect 47952 16600 48004 16652
rect 48044 16600 48096 16652
rect 51356 16668 51408 16720
rect 53840 16736 53892 16788
rect 54852 16736 54904 16788
rect 56600 16736 56652 16788
rect 53564 16668 53616 16720
rect 55312 16600 55364 16652
rect 55772 16600 55824 16652
rect 47492 16532 47544 16584
rect 47768 16575 47820 16584
rect 47768 16541 47778 16575
rect 47778 16541 47812 16575
rect 47812 16541 47820 16575
rect 47768 16532 47820 16541
rect 39396 16439 39448 16448
rect 39396 16405 39405 16439
rect 39405 16405 39439 16439
rect 39439 16405 39448 16439
rect 39396 16396 39448 16405
rect 39672 16396 39724 16448
rect 40316 16396 40368 16448
rect 41144 16439 41196 16448
rect 41144 16405 41153 16439
rect 41153 16405 41187 16439
rect 41187 16405 41196 16439
rect 41144 16396 41196 16405
rect 42064 16396 42116 16448
rect 42616 16439 42668 16448
rect 42616 16405 42625 16439
rect 42625 16405 42659 16439
rect 42659 16405 42668 16439
rect 46848 16464 46900 16516
rect 47584 16464 47636 16516
rect 48044 16507 48096 16516
rect 48044 16473 48053 16507
rect 48053 16473 48087 16507
rect 48087 16473 48096 16507
rect 48044 16464 48096 16473
rect 48596 16575 48648 16584
rect 48596 16541 48605 16575
rect 48605 16541 48639 16575
rect 48639 16541 48648 16575
rect 48596 16532 48648 16541
rect 48872 16532 48924 16584
rect 49332 16532 49384 16584
rect 49424 16575 49476 16584
rect 49424 16541 49433 16575
rect 49433 16541 49467 16575
rect 49467 16541 49476 16575
rect 49424 16532 49476 16541
rect 49608 16575 49660 16584
rect 49608 16541 49617 16575
rect 49617 16541 49651 16575
rect 49651 16541 49660 16575
rect 49608 16532 49660 16541
rect 54116 16532 54168 16584
rect 48320 16464 48372 16516
rect 49056 16507 49108 16516
rect 49056 16473 49065 16507
rect 49065 16473 49099 16507
rect 49099 16473 49108 16507
rect 49056 16464 49108 16473
rect 49148 16464 49200 16516
rect 42616 16396 42668 16405
rect 43812 16439 43864 16448
rect 43812 16405 43821 16439
rect 43821 16405 43855 16439
rect 43855 16405 43864 16439
rect 43812 16396 43864 16405
rect 48228 16396 48280 16448
rect 48596 16396 48648 16448
rect 50344 16464 50396 16516
rect 53932 16464 53984 16516
rect 57520 16575 57572 16584
rect 57520 16541 57529 16575
rect 57529 16541 57563 16575
rect 57563 16541 57572 16575
rect 57520 16532 57572 16541
rect 55312 16507 55364 16516
rect 55312 16473 55321 16507
rect 55321 16473 55355 16507
rect 55355 16473 55364 16507
rect 55312 16464 55364 16473
rect 55956 16464 56008 16516
rect 54116 16396 54168 16448
rect 57244 16507 57296 16516
rect 57244 16473 57253 16507
rect 57253 16473 57287 16507
rect 57287 16473 57296 16507
rect 57244 16464 57296 16473
rect 57336 16507 57388 16516
rect 57336 16473 57345 16507
rect 57345 16473 57379 16507
rect 57379 16473 57388 16507
rect 57336 16464 57388 16473
rect 56968 16439 57020 16448
rect 56968 16405 56977 16439
rect 56977 16405 57011 16439
rect 57011 16405 57020 16439
rect 56968 16396 57020 16405
rect 4874 16294 4926 16346
rect 4938 16294 4990 16346
rect 5002 16294 5054 16346
rect 5066 16294 5118 16346
rect 5130 16294 5182 16346
rect 35594 16294 35646 16346
rect 35658 16294 35710 16346
rect 35722 16294 35774 16346
rect 35786 16294 35838 16346
rect 35850 16294 35902 16346
rect 19524 16192 19576 16244
rect 19800 16192 19852 16244
rect 20260 16192 20312 16244
rect 20812 16192 20864 16244
rect 21640 16192 21692 16244
rect 22376 16192 22428 16244
rect 23204 16192 23256 16244
rect 24952 16235 25004 16244
rect 24952 16201 24961 16235
rect 24961 16201 24995 16235
rect 24995 16201 25004 16235
rect 24952 16192 25004 16201
rect 25136 16192 25188 16244
rect 19524 16099 19576 16108
rect 19524 16065 19533 16099
rect 19533 16065 19567 16099
rect 19567 16065 19576 16099
rect 19524 16056 19576 16065
rect 18972 15988 19024 16040
rect 19708 16056 19760 16108
rect 23020 16124 23072 16176
rect 24676 16167 24728 16176
rect 24676 16133 24685 16167
rect 24685 16133 24719 16167
rect 24719 16133 24728 16167
rect 24676 16124 24728 16133
rect 29184 16235 29236 16244
rect 29184 16201 29193 16235
rect 29193 16201 29227 16235
rect 29227 16201 29236 16235
rect 29184 16192 29236 16201
rect 20168 15988 20220 16040
rect 21640 16031 21692 16040
rect 21640 15997 21649 16031
rect 21649 15997 21683 16031
rect 21683 15997 21692 16031
rect 21640 15988 21692 15997
rect 20076 15920 20128 15972
rect 21548 15963 21600 15972
rect 21548 15929 21557 15963
rect 21557 15929 21591 15963
rect 21591 15929 21600 15963
rect 21548 15920 21600 15929
rect 22192 16099 22244 16108
rect 22192 16065 22201 16099
rect 22201 16065 22235 16099
rect 22235 16065 22244 16099
rect 22192 16056 22244 16065
rect 22284 16099 22336 16108
rect 22284 16065 22329 16099
rect 22329 16065 22336 16099
rect 22284 16056 22336 16065
rect 22468 16099 22520 16108
rect 22468 16065 22477 16099
rect 22477 16065 22511 16099
rect 22511 16065 22520 16099
rect 22468 16056 22520 16065
rect 23296 16099 23348 16108
rect 23296 16065 23300 16099
rect 23300 16065 23334 16099
rect 23334 16065 23348 16099
rect 23296 16056 23348 16065
rect 23480 16099 23532 16108
rect 23480 16065 23489 16099
rect 23489 16065 23523 16099
rect 23523 16065 23532 16099
rect 23480 16056 23532 16065
rect 23664 16099 23716 16108
rect 23664 16065 23672 16099
rect 23672 16065 23706 16099
rect 23706 16065 23716 16099
rect 23664 16056 23716 16065
rect 23848 16056 23900 16108
rect 24768 16099 24820 16108
rect 24768 16065 24777 16099
rect 24777 16065 24811 16099
rect 24811 16065 24820 16099
rect 24768 16056 24820 16065
rect 25044 16056 25096 16108
rect 25136 15988 25188 16040
rect 22468 15920 22520 15972
rect 22836 15920 22888 15972
rect 23756 15920 23808 15972
rect 25872 16056 25924 16108
rect 26424 16099 26476 16108
rect 26424 16065 26433 16099
rect 26433 16065 26467 16099
rect 26467 16065 26476 16099
rect 26424 16056 26476 16065
rect 27344 16167 27396 16176
rect 27344 16133 27353 16167
rect 27353 16133 27387 16167
rect 27387 16133 27396 16167
rect 27344 16124 27396 16133
rect 29276 16124 29328 16176
rect 26700 15988 26752 16040
rect 26884 15988 26936 16040
rect 27528 16099 27580 16108
rect 30380 16192 30432 16244
rect 31116 16235 31168 16244
rect 31116 16201 31125 16235
rect 31125 16201 31159 16235
rect 31159 16201 31168 16235
rect 31116 16192 31168 16201
rect 32772 16192 32824 16244
rect 35256 16192 35308 16244
rect 35808 16192 35860 16244
rect 29644 16167 29696 16176
rect 29644 16133 29653 16167
rect 29653 16133 29687 16167
rect 29687 16133 29696 16167
rect 29644 16124 29696 16133
rect 30656 16124 30708 16176
rect 33508 16124 33560 16176
rect 27528 16065 27542 16099
rect 27542 16065 27576 16099
rect 27576 16065 27580 16099
rect 27528 16056 27580 16065
rect 31208 16099 31260 16108
rect 31208 16065 31217 16099
rect 31217 16065 31251 16099
rect 31251 16065 31260 16099
rect 31208 16056 31260 16065
rect 31760 16056 31812 16108
rect 35348 16124 35400 16176
rect 36176 16192 36228 16244
rect 38660 16192 38712 16244
rect 38936 16192 38988 16244
rect 39028 16124 39080 16176
rect 26516 15920 26568 15972
rect 26792 15963 26844 15972
rect 26792 15929 26801 15963
rect 26801 15929 26835 15963
rect 26835 15929 26844 15963
rect 26792 15920 26844 15929
rect 24584 15852 24636 15904
rect 24768 15852 24820 15904
rect 26056 15852 26108 15904
rect 26148 15852 26200 15904
rect 36084 16056 36136 16108
rect 36544 16056 36596 16108
rect 34888 15988 34940 16040
rect 35440 15988 35492 16040
rect 36820 16099 36872 16108
rect 36820 16065 36829 16099
rect 36829 16065 36863 16099
rect 36863 16065 36872 16099
rect 36820 16056 36872 16065
rect 37004 16099 37056 16108
rect 37004 16065 37013 16099
rect 37013 16065 37047 16099
rect 37047 16065 37056 16099
rect 37004 16056 37056 16065
rect 37832 16056 37884 16108
rect 27896 15852 27948 15904
rect 27988 15852 28040 15904
rect 29736 15852 29788 15904
rect 35992 15920 36044 15972
rect 37464 15988 37516 16040
rect 37004 15920 37056 15972
rect 38200 16056 38252 16108
rect 38568 16056 38620 16108
rect 38660 16099 38712 16108
rect 38660 16065 38669 16099
rect 38669 16065 38703 16099
rect 38703 16065 38712 16099
rect 38660 16056 38712 16065
rect 39488 16167 39540 16176
rect 39488 16133 39497 16167
rect 39497 16133 39531 16167
rect 39531 16133 39540 16167
rect 39488 16124 39540 16133
rect 39856 16235 39908 16244
rect 39856 16201 39865 16235
rect 39865 16201 39899 16235
rect 39899 16201 39908 16235
rect 39856 16192 39908 16201
rect 38844 15988 38896 16040
rect 31024 15852 31076 15904
rect 34060 15852 34112 15904
rect 35716 15895 35768 15904
rect 35716 15861 35725 15895
rect 35725 15861 35759 15895
rect 35759 15861 35768 15895
rect 35716 15852 35768 15861
rect 35808 15852 35860 15904
rect 36820 15852 36872 15904
rect 37832 15895 37884 15904
rect 37832 15861 37841 15895
rect 37841 15861 37875 15895
rect 37875 15861 37884 15895
rect 37832 15852 37884 15861
rect 38108 15895 38160 15904
rect 38108 15861 38117 15895
rect 38117 15861 38151 15895
rect 38151 15861 38160 15895
rect 38108 15852 38160 15861
rect 38568 15852 38620 15904
rect 39948 16056 40000 16108
rect 41236 16192 41288 16244
rect 44180 16192 44232 16244
rect 47584 16192 47636 16244
rect 47676 16192 47728 16244
rect 48412 16192 48464 16244
rect 49608 16192 49660 16244
rect 49700 16235 49752 16244
rect 49700 16201 49709 16235
rect 49709 16201 49743 16235
rect 49743 16201 49752 16235
rect 49700 16192 49752 16201
rect 40316 16167 40368 16176
rect 40316 16133 40325 16167
rect 40325 16133 40359 16167
rect 40359 16133 40368 16167
rect 40316 16124 40368 16133
rect 40868 16124 40920 16176
rect 42800 16124 42852 16176
rect 50252 16192 50304 16244
rect 53288 16235 53340 16244
rect 53288 16201 53297 16235
rect 53297 16201 53331 16235
rect 53331 16201 53340 16235
rect 53288 16192 53340 16201
rect 53380 16192 53432 16244
rect 54760 16192 54812 16244
rect 56048 16192 56100 16244
rect 43996 16056 44048 16108
rect 40408 15988 40460 16040
rect 39396 15920 39448 15972
rect 39672 15920 39724 15972
rect 41788 15895 41840 15904
rect 41788 15861 41797 15895
rect 41797 15861 41831 15895
rect 41831 15861 41840 15895
rect 41788 15852 41840 15861
rect 43260 15988 43312 16040
rect 44548 15988 44600 16040
rect 44732 16099 44784 16108
rect 44732 16065 44741 16099
rect 44741 16065 44775 16099
rect 44775 16065 44784 16099
rect 44732 16056 44784 16065
rect 46572 16099 46624 16108
rect 46572 16065 46581 16099
rect 46581 16065 46615 16099
rect 46615 16065 46624 16099
rect 46572 16056 46624 16065
rect 47400 16056 47452 16108
rect 47768 16056 47820 16108
rect 43444 15852 43496 15904
rect 43628 15852 43680 15904
rect 45376 15988 45428 16040
rect 48228 15988 48280 16040
rect 48596 16099 48648 16108
rect 48596 16065 48605 16099
rect 48605 16065 48639 16099
rect 48639 16065 48648 16099
rect 48596 16056 48648 16065
rect 48688 16099 48740 16108
rect 48688 16065 48697 16099
rect 48697 16065 48731 16099
rect 48731 16065 48740 16099
rect 48688 16056 48740 16065
rect 48044 15920 48096 15972
rect 45652 15852 45704 15904
rect 45928 15852 45980 15904
rect 48412 15920 48464 15972
rect 48964 16056 49016 16108
rect 49424 16099 49476 16108
rect 49424 16065 49433 16099
rect 49433 16065 49467 16099
rect 49467 16065 49476 16099
rect 49424 16056 49476 16065
rect 49700 16056 49752 16108
rect 50068 16099 50120 16108
rect 50068 16065 50077 16099
rect 50077 16065 50111 16099
rect 50111 16065 50120 16099
rect 50068 16056 50120 16065
rect 51356 16056 51408 16108
rect 50160 15988 50212 16040
rect 51080 15988 51132 16040
rect 54760 16099 54812 16108
rect 54760 16065 54769 16099
rect 54769 16065 54803 16099
rect 54803 16065 54812 16099
rect 54760 16056 54812 16065
rect 54944 16056 54996 16108
rect 55312 16167 55364 16176
rect 55312 16133 55321 16167
rect 55321 16133 55355 16167
rect 55355 16133 55364 16167
rect 55312 16124 55364 16133
rect 56692 16124 56744 16176
rect 55680 16056 55732 16108
rect 53932 15988 53984 16040
rect 56600 15988 56652 16040
rect 49056 15920 49108 15972
rect 52920 15920 52972 15972
rect 55404 15920 55456 15972
rect 52828 15852 52880 15904
rect 53748 15852 53800 15904
rect 55956 15852 56008 15904
rect 57244 15852 57296 15904
rect 57704 15895 57756 15904
rect 57704 15861 57713 15895
rect 57713 15861 57747 15895
rect 57747 15861 57756 15895
rect 57704 15852 57756 15861
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 13268 15512 13320 15564
rect 18880 15648 18932 15700
rect 20076 15648 20128 15700
rect 20168 15648 20220 15700
rect 22192 15648 22244 15700
rect 22560 15648 22612 15700
rect 23480 15648 23532 15700
rect 24216 15648 24268 15700
rect 24676 15648 24728 15700
rect 19984 15580 20036 15632
rect 24492 15580 24544 15632
rect 24860 15691 24912 15700
rect 24860 15657 24869 15691
rect 24869 15657 24903 15691
rect 24903 15657 24912 15691
rect 24860 15648 24912 15657
rect 26608 15648 26660 15700
rect 26332 15580 26384 15632
rect 26700 15580 26752 15632
rect 28724 15580 28776 15632
rect 21548 15512 21600 15564
rect 23572 15512 23624 15564
rect 23848 15512 23900 15564
rect 24032 15512 24084 15564
rect 24768 15512 24820 15564
rect 26516 15512 26568 15564
rect 30196 15512 30248 15564
rect 14924 15444 14976 15496
rect 12624 15376 12676 15428
rect 12716 15308 12768 15360
rect 13452 15419 13504 15428
rect 13452 15385 13461 15419
rect 13461 15385 13495 15419
rect 13495 15385 13504 15419
rect 13452 15376 13504 15385
rect 19800 15487 19852 15496
rect 19800 15453 19809 15487
rect 19809 15453 19843 15487
rect 19843 15453 19852 15487
rect 19800 15444 19852 15453
rect 20076 15487 20128 15496
rect 20076 15453 20085 15487
rect 20085 15453 20119 15487
rect 20119 15453 20128 15487
rect 20076 15444 20128 15453
rect 20260 15444 20312 15496
rect 22192 15487 22244 15496
rect 22192 15453 22201 15487
rect 22201 15453 22235 15487
rect 22235 15453 22244 15487
rect 22192 15444 22244 15453
rect 22376 15487 22428 15496
rect 22376 15453 22385 15487
rect 22385 15453 22419 15487
rect 22419 15453 22428 15487
rect 22376 15444 22428 15453
rect 22928 15487 22980 15496
rect 22928 15453 22937 15487
rect 22937 15453 22971 15487
rect 22971 15453 22980 15487
rect 22928 15444 22980 15453
rect 23112 15487 23164 15496
rect 23112 15453 23121 15487
rect 23121 15453 23155 15487
rect 23155 15453 23164 15487
rect 23112 15444 23164 15453
rect 23388 15444 23440 15496
rect 24492 15444 24544 15496
rect 23296 15419 23348 15428
rect 23296 15385 23305 15419
rect 23305 15385 23339 15419
rect 23339 15385 23348 15419
rect 23296 15376 23348 15385
rect 24124 15419 24176 15428
rect 24124 15385 24133 15419
rect 24133 15385 24167 15419
rect 24167 15385 24176 15419
rect 24124 15376 24176 15385
rect 25688 15487 25740 15496
rect 25688 15453 25697 15487
rect 25697 15453 25731 15487
rect 25731 15453 25740 15487
rect 25688 15444 25740 15453
rect 29644 15444 29696 15496
rect 25964 15376 26016 15428
rect 26700 15376 26752 15428
rect 27344 15376 27396 15428
rect 15108 15308 15160 15360
rect 18144 15308 18196 15360
rect 20720 15308 20772 15360
rect 21732 15308 21784 15360
rect 22100 15308 22152 15360
rect 23480 15308 23532 15360
rect 26240 15308 26292 15360
rect 34520 15648 34572 15700
rect 30288 15487 30340 15496
rect 30288 15453 30297 15487
rect 30297 15453 30331 15487
rect 30331 15453 30340 15487
rect 30288 15444 30340 15453
rect 30472 15444 30524 15496
rect 31024 15623 31076 15632
rect 31024 15589 31033 15623
rect 31033 15589 31067 15623
rect 31067 15589 31076 15623
rect 31024 15580 31076 15589
rect 36544 15648 36596 15700
rect 38292 15648 38344 15700
rect 30748 15512 30800 15564
rect 32128 15555 32180 15564
rect 32128 15521 32137 15555
rect 32137 15521 32171 15555
rect 32171 15521 32180 15555
rect 32128 15512 32180 15521
rect 32588 15444 32640 15496
rect 33508 15512 33560 15564
rect 35716 15512 35768 15564
rect 38200 15512 38252 15564
rect 38660 15580 38712 15632
rect 39028 15691 39080 15700
rect 39028 15657 39037 15691
rect 39037 15657 39071 15691
rect 39071 15657 39080 15691
rect 39028 15648 39080 15657
rect 39120 15580 39172 15632
rect 40316 15648 40368 15700
rect 40684 15648 40736 15700
rect 43076 15648 43128 15700
rect 47676 15648 47728 15700
rect 48780 15648 48832 15700
rect 49240 15648 49292 15700
rect 51356 15648 51408 15700
rect 54760 15648 54812 15700
rect 39488 15580 39540 15632
rect 42616 15580 42668 15632
rect 48044 15623 48096 15632
rect 48044 15589 48053 15623
rect 48053 15589 48087 15623
rect 48087 15589 48096 15623
rect 48044 15580 48096 15589
rect 48596 15580 48648 15632
rect 48688 15580 48740 15632
rect 51908 15623 51960 15632
rect 51908 15589 51917 15623
rect 51917 15589 51951 15623
rect 51951 15589 51960 15623
rect 51908 15580 51960 15589
rect 40040 15512 40092 15564
rect 37280 15487 37332 15496
rect 37280 15453 37289 15487
rect 37289 15453 37323 15487
rect 37323 15453 37332 15487
rect 37280 15444 37332 15453
rect 39028 15444 39080 15496
rect 40224 15487 40276 15496
rect 40224 15453 40233 15487
rect 40233 15453 40267 15487
rect 40267 15453 40276 15487
rect 40224 15444 40276 15453
rect 40316 15487 40368 15496
rect 40316 15453 40325 15487
rect 40325 15453 40359 15487
rect 40359 15453 40368 15487
rect 40316 15444 40368 15453
rect 43444 15512 43496 15564
rect 44916 15512 44968 15564
rect 47952 15512 48004 15564
rect 49884 15512 49936 15564
rect 29828 15376 29880 15428
rect 32772 15376 32824 15428
rect 30472 15308 30524 15360
rect 36728 15376 36780 15428
rect 37556 15419 37608 15428
rect 37556 15385 37565 15419
rect 37565 15385 37599 15419
rect 37599 15385 37608 15419
rect 37556 15376 37608 15385
rect 37372 15308 37424 15360
rect 39212 15376 39264 15428
rect 39304 15376 39356 15428
rect 39856 15376 39908 15428
rect 41788 15444 41840 15496
rect 43352 15444 43404 15496
rect 43536 15487 43588 15496
rect 43536 15453 43545 15487
rect 43545 15453 43579 15487
rect 43579 15453 43588 15487
rect 43536 15444 43588 15453
rect 43628 15444 43680 15496
rect 44088 15444 44140 15496
rect 39580 15308 39632 15360
rect 40500 15376 40552 15428
rect 40868 15376 40920 15428
rect 40960 15376 41012 15428
rect 42524 15376 42576 15428
rect 40684 15351 40736 15360
rect 40684 15317 40693 15351
rect 40693 15317 40727 15351
rect 40727 15317 40736 15351
rect 40684 15308 40736 15317
rect 41512 15308 41564 15360
rect 43996 15376 44048 15428
rect 44548 15308 44600 15360
rect 45928 15419 45980 15428
rect 45928 15385 45937 15419
rect 45937 15385 45971 15419
rect 45971 15385 45980 15419
rect 45928 15376 45980 15385
rect 47308 15376 47360 15428
rect 47860 15376 47912 15428
rect 48780 15487 48832 15496
rect 48780 15453 48789 15487
rect 48789 15453 48823 15487
rect 48823 15453 48832 15487
rect 48780 15444 48832 15453
rect 51356 15487 51408 15496
rect 51356 15453 51365 15487
rect 51365 15453 51399 15487
rect 51399 15453 51408 15487
rect 51356 15444 51408 15453
rect 52092 15512 52144 15564
rect 52460 15623 52512 15632
rect 52460 15589 52469 15623
rect 52469 15589 52503 15623
rect 52503 15589 52512 15623
rect 52460 15580 52512 15589
rect 53288 15580 53340 15632
rect 51724 15487 51776 15496
rect 51724 15453 51733 15487
rect 51733 15453 51767 15487
rect 51767 15453 51776 15487
rect 51724 15444 51776 15453
rect 49332 15376 49384 15428
rect 51908 15376 51960 15428
rect 46664 15308 46716 15360
rect 47400 15351 47452 15360
rect 47400 15317 47409 15351
rect 47409 15317 47443 15351
rect 47443 15317 47452 15351
rect 47400 15308 47452 15317
rect 48688 15308 48740 15360
rect 49056 15308 49108 15360
rect 51724 15308 51776 15360
rect 52552 15487 52604 15496
rect 52552 15453 52561 15487
rect 52561 15453 52595 15487
rect 52595 15453 52604 15487
rect 52552 15444 52604 15453
rect 52828 15487 52880 15496
rect 52828 15453 52837 15487
rect 52837 15453 52871 15487
rect 52871 15453 52880 15487
rect 52828 15444 52880 15453
rect 53196 15487 53248 15496
rect 53196 15453 53205 15487
rect 53205 15453 53239 15487
rect 53239 15453 53248 15487
rect 53196 15444 53248 15453
rect 53564 15444 53616 15496
rect 52920 15376 52972 15428
rect 53288 15376 53340 15428
rect 54116 15512 54168 15564
rect 56232 15648 56284 15700
rect 56600 15691 56652 15700
rect 56600 15657 56609 15691
rect 56609 15657 56643 15691
rect 56643 15657 56652 15691
rect 56600 15648 56652 15657
rect 52736 15351 52788 15360
rect 52736 15317 52745 15351
rect 52745 15317 52779 15351
rect 52779 15317 52788 15351
rect 52736 15308 52788 15317
rect 53840 15308 53892 15360
rect 55220 15308 55272 15360
rect 55680 15487 55732 15496
rect 55680 15453 55689 15487
rect 55689 15453 55723 15487
rect 55723 15453 55732 15487
rect 55680 15444 55732 15453
rect 55404 15376 55456 15428
rect 57336 15580 57388 15632
rect 56048 15555 56100 15564
rect 56048 15521 56057 15555
rect 56057 15521 56091 15555
rect 56091 15521 56100 15555
rect 56048 15512 56100 15521
rect 55956 15487 56008 15496
rect 55956 15453 55965 15487
rect 55965 15453 55999 15487
rect 55999 15453 56008 15487
rect 55956 15444 56008 15453
rect 56232 15487 56284 15496
rect 56232 15453 56241 15487
rect 56241 15453 56275 15487
rect 56275 15453 56284 15487
rect 56232 15444 56284 15453
rect 56324 15487 56376 15496
rect 56324 15453 56333 15487
rect 56333 15453 56367 15487
rect 56367 15453 56376 15487
rect 56324 15444 56376 15453
rect 56968 15444 57020 15496
rect 57704 15444 57756 15496
rect 56508 15351 56560 15360
rect 56508 15317 56517 15351
rect 56517 15317 56551 15351
rect 56551 15317 56560 15351
rect 56508 15308 56560 15317
rect 4874 15206 4926 15258
rect 4938 15206 4990 15258
rect 5002 15206 5054 15258
rect 5066 15206 5118 15258
rect 5130 15206 5182 15258
rect 35594 15206 35646 15258
rect 35658 15206 35710 15258
rect 35722 15206 35774 15258
rect 35786 15206 35838 15258
rect 35850 15206 35902 15258
rect 12624 15011 12676 15020
rect 12624 14977 12633 15011
rect 12633 14977 12667 15011
rect 12667 14977 12676 15011
rect 12624 14968 12676 14977
rect 12900 15011 12952 15020
rect 12900 14977 12909 15011
rect 12909 14977 12943 15011
rect 12943 14977 12952 15011
rect 12900 14968 12952 14977
rect 16672 15104 16724 15156
rect 13268 15079 13320 15088
rect 13268 15045 13277 15079
rect 13277 15045 13311 15079
rect 13311 15045 13320 15079
rect 13268 15036 13320 15045
rect 18052 15036 18104 15088
rect 18144 15079 18196 15088
rect 18144 15045 18153 15079
rect 18153 15045 18187 15079
rect 18187 15045 18196 15079
rect 18144 15036 18196 15045
rect 20076 15104 20128 15156
rect 22192 15147 22244 15156
rect 22192 15113 22201 15147
rect 22201 15113 22235 15147
rect 22235 15113 22244 15147
rect 22192 15104 22244 15113
rect 22376 15104 22428 15156
rect 23112 15104 23164 15156
rect 23204 15147 23256 15156
rect 23204 15113 23213 15147
rect 23213 15113 23247 15147
rect 23247 15113 23256 15147
rect 23204 15104 23256 15113
rect 25688 15104 25740 15156
rect 26148 15104 26200 15156
rect 19984 15079 20036 15088
rect 19984 15045 19993 15079
rect 19993 15045 20027 15079
rect 20027 15045 20036 15079
rect 19984 15036 20036 15045
rect 14740 14968 14792 15020
rect 13636 14900 13688 14952
rect 15476 14900 15528 14952
rect 17868 14943 17920 14952
rect 17868 14909 17877 14943
rect 17877 14909 17911 14943
rect 17911 14909 17920 14943
rect 17868 14900 17920 14909
rect 12348 14764 12400 14816
rect 14924 14764 14976 14816
rect 16120 14764 16172 14816
rect 19708 14968 19760 15020
rect 19616 14900 19668 14952
rect 20168 14968 20220 15020
rect 20260 15011 20312 15020
rect 20260 14977 20268 15011
rect 20268 14977 20302 15011
rect 20302 14977 20312 15011
rect 20260 14968 20312 14977
rect 20352 15011 20404 15020
rect 20352 14977 20361 15011
rect 20361 14977 20395 15011
rect 20395 14977 20404 15011
rect 20352 14968 20404 14977
rect 20628 14968 20680 15020
rect 21916 14968 21968 15020
rect 22560 15011 22612 15020
rect 22560 14977 22569 15011
rect 22569 14977 22603 15011
rect 22603 14977 22612 15011
rect 22560 14968 22612 14977
rect 22744 15011 22796 15020
rect 22744 14977 22752 15011
rect 22752 14977 22786 15011
rect 22786 14977 22796 15011
rect 22744 14968 22796 14977
rect 22836 15011 22888 15020
rect 22836 14977 22845 15011
rect 22845 14977 22879 15011
rect 22879 14977 22888 15011
rect 22836 14968 22888 14977
rect 23020 15011 23072 15020
rect 23020 14977 23029 15011
rect 23029 14977 23063 15011
rect 23063 14977 23072 15011
rect 25872 15079 25924 15088
rect 25872 15045 25881 15079
rect 25881 15045 25915 15079
rect 25915 15045 25924 15079
rect 25872 15036 25924 15045
rect 25964 15079 26016 15088
rect 25964 15045 25973 15079
rect 25973 15045 26007 15079
rect 26007 15045 26016 15079
rect 25964 15036 26016 15045
rect 23020 14968 23072 14977
rect 24124 14968 24176 15020
rect 24860 14968 24912 15020
rect 32128 15104 32180 15156
rect 37556 15104 37608 15156
rect 38568 15104 38620 15156
rect 39488 15147 39540 15156
rect 39488 15113 39497 15147
rect 39497 15113 39531 15147
rect 39531 15113 39540 15147
rect 39488 15104 39540 15113
rect 39672 15147 39724 15156
rect 39672 15113 39681 15147
rect 39681 15113 39715 15147
rect 39715 15113 39724 15147
rect 39672 15104 39724 15113
rect 30472 15079 30524 15088
rect 30472 15045 30481 15079
rect 30481 15045 30515 15079
rect 30515 15045 30524 15079
rect 30472 15036 30524 15045
rect 30564 15036 30616 15088
rect 34244 15036 34296 15088
rect 42064 15104 42116 15156
rect 42156 15104 42208 15156
rect 43076 15104 43128 15156
rect 41512 15036 41564 15088
rect 43996 15104 44048 15156
rect 46572 15104 46624 15156
rect 49884 15147 49936 15156
rect 49884 15113 49893 15147
rect 49893 15113 49927 15147
rect 49927 15113 49936 15147
rect 49884 15104 49936 15113
rect 49976 15147 50028 15156
rect 49976 15113 49985 15147
rect 49985 15113 50019 15147
rect 50019 15113 50028 15147
rect 49976 15104 50028 15113
rect 19800 14832 19852 14884
rect 25320 14900 25372 14952
rect 22744 14832 22796 14884
rect 23388 14832 23440 14884
rect 35440 14968 35492 15020
rect 30196 14943 30248 14952
rect 30196 14909 30205 14943
rect 30205 14909 30239 14943
rect 30239 14909 30248 14943
rect 30196 14900 30248 14909
rect 20444 14764 20496 14816
rect 26792 14832 26844 14884
rect 30932 14900 30984 14952
rect 37924 15011 37976 15020
rect 37924 14977 37933 15011
rect 37933 14977 37967 15011
rect 37967 14977 37976 15011
rect 37924 14968 37976 14977
rect 38108 14968 38160 15020
rect 39028 14968 39080 15020
rect 41236 14968 41288 15020
rect 42616 14968 42668 15020
rect 42800 15011 42852 15020
rect 42800 14977 42809 15011
rect 42809 14977 42843 15011
rect 42843 14977 42852 15011
rect 42800 14968 42852 14977
rect 46020 15036 46072 15088
rect 46388 15036 46440 15088
rect 47860 15036 47912 15088
rect 52460 15104 52512 15156
rect 52368 15079 52420 15088
rect 52368 15045 52377 15079
rect 52377 15045 52411 15079
rect 52411 15045 52420 15079
rect 52368 15036 52420 15045
rect 37464 14900 37516 14952
rect 38384 14900 38436 14952
rect 40132 14900 40184 14952
rect 41420 14900 41472 14952
rect 41512 14900 41564 14952
rect 43444 14900 43496 14952
rect 44916 15011 44968 15020
rect 44916 14977 44925 15011
rect 44925 14977 44959 15011
rect 44959 14977 44968 15011
rect 44916 14968 44968 14977
rect 46664 15011 46716 15020
rect 46664 14977 46668 15011
rect 46668 14977 46702 15011
rect 46702 14977 46716 15011
rect 46664 14968 46716 14977
rect 34336 14832 34388 14884
rect 25872 14764 25924 14816
rect 27160 14764 27212 14816
rect 34704 14764 34756 14816
rect 36452 14764 36504 14816
rect 37832 14764 37884 14816
rect 38200 14807 38252 14816
rect 38200 14773 38209 14807
rect 38209 14773 38243 14807
rect 38243 14773 38252 14807
rect 38200 14764 38252 14773
rect 40040 14832 40092 14884
rect 40960 14832 41012 14884
rect 42156 14832 42208 14884
rect 42340 14832 42392 14884
rect 42432 14764 42484 14816
rect 42708 14764 42760 14816
rect 43076 14764 43128 14816
rect 43260 14832 43312 14884
rect 44180 14900 44232 14952
rect 44272 14900 44324 14952
rect 47216 14968 47268 15020
rect 47952 14968 48004 15020
rect 51816 15011 51868 15020
rect 51816 14977 51825 15011
rect 51825 14977 51859 15011
rect 51859 14977 51868 15011
rect 51816 14968 51868 14977
rect 53932 15104 53984 15156
rect 55128 15104 55180 15156
rect 53288 15079 53340 15088
rect 53288 15045 53297 15079
rect 53297 15045 53331 15079
rect 53331 15045 53340 15079
rect 53288 15036 53340 15045
rect 53748 15036 53800 15088
rect 56508 15036 56560 15088
rect 49700 14900 49752 14952
rect 50068 14900 50120 14952
rect 52552 14900 52604 14952
rect 53012 14943 53064 14952
rect 53012 14909 53021 14943
rect 53021 14909 53055 14943
rect 53055 14909 53064 14943
rect 53012 14900 53064 14909
rect 53748 14900 53800 14952
rect 44088 14764 44140 14816
rect 44640 14764 44692 14816
rect 45100 14764 45152 14816
rect 47124 14764 47176 14816
rect 47216 14807 47268 14816
rect 47216 14773 47225 14807
rect 47225 14773 47259 14807
rect 47259 14773 47268 14807
rect 47216 14764 47268 14773
rect 48228 14764 48280 14816
rect 48413 14807 48465 14816
rect 48413 14773 48442 14807
rect 48442 14773 48465 14807
rect 48413 14764 48465 14773
rect 54760 14943 54812 14952
rect 54760 14909 54769 14943
rect 54769 14909 54803 14943
rect 54803 14909 54812 14943
rect 54760 14900 54812 14909
rect 55036 14900 55088 14952
rect 55956 14900 56008 14952
rect 56692 14764 56744 14816
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 12900 14560 12952 14612
rect 19708 14560 19760 14612
rect 20260 14560 20312 14612
rect 22928 14560 22980 14612
rect 12716 14467 12768 14476
rect 1216 14356 1268 14408
rect 12716 14433 12725 14467
rect 12725 14433 12759 14467
rect 12759 14433 12768 14467
rect 12716 14424 12768 14433
rect 13176 14424 13228 14476
rect 13452 14424 13504 14476
rect 14740 14467 14792 14476
rect 14740 14433 14749 14467
rect 14749 14433 14783 14467
rect 14783 14433 14792 14467
rect 14740 14424 14792 14433
rect 15200 14424 15252 14476
rect 17316 14424 17368 14476
rect 17868 14424 17920 14476
rect 18052 14424 18104 14476
rect 20628 14424 20680 14476
rect 20720 14467 20772 14476
rect 20720 14433 20729 14467
rect 20729 14433 20763 14467
rect 20763 14433 20772 14467
rect 20720 14424 20772 14433
rect 21732 14467 21784 14476
rect 21732 14433 21741 14467
rect 21741 14433 21775 14467
rect 21775 14433 21784 14467
rect 21732 14424 21784 14433
rect 12348 14399 12400 14408
rect 12348 14365 12357 14399
rect 12357 14365 12391 14399
rect 12391 14365 12400 14399
rect 12348 14356 12400 14365
rect 11704 14288 11756 14340
rect 15292 14356 15344 14408
rect 21456 14399 21508 14408
rect 21456 14365 21465 14399
rect 21465 14365 21499 14399
rect 21499 14365 21508 14399
rect 21456 14356 21508 14365
rect 17960 14288 18012 14340
rect 19432 14288 19484 14340
rect 20444 14288 20496 14340
rect 22008 14288 22060 14340
rect 22192 14288 22244 14340
rect 23112 14492 23164 14544
rect 24768 14603 24820 14612
rect 24768 14569 24777 14603
rect 24777 14569 24811 14603
rect 24811 14569 24820 14603
rect 24768 14560 24820 14569
rect 23204 14356 23256 14408
rect 23572 14399 23624 14408
rect 23572 14365 23581 14399
rect 23581 14365 23615 14399
rect 23615 14365 23624 14399
rect 23572 14356 23624 14365
rect 12256 14263 12308 14272
rect 12256 14229 12265 14263
rect 12265 14229 12299 14263
rect 12299 14229 12308 14263
rect 12256 14220 12308 14229
rect 15476 14263 15528 14272
rect 15476 14229 15485 14263
rect 15485 14229 15519 14263
rect 15519 14229 15528 14263
rect 15476 14220 15528 14229
rect 16764 14220 16816 14272
rect 18144 14220 18196 14272
rect 19156 14220 19208 14272
rect 19892 14220 19944 14272
rect 23480 14220 23532 14272
rect 23756 14288 23808 14340
rect 24216 14356 24268 14408
rect 24676 14399 24728 14408
rect 24676 14365 24685 14399
rect 24685 14365 24719 14399
rect 24719 14365 24728 14399
rect 24676 14356 24728 14365
rect 26700 14603 26752 14612
rect 26700 14569 26709 14603
rect 26709 14569 26743 14603
rect 26743 14569 26752 14603
rect 26700 14560 26752 14569
rect 28356 14560 28408 14612
rect 30288 14560 30340 14612
rect 34336 14603 34388 14612
rect 34336 14569 34345 14603
rect 34345 14569 34379 14603
rect 34379 14569 34388 14603
rect 34336 14560 34388 14569
rect 35992 14560 36044 14612
rect 36268 14560 36320 14612
rect 36912 14560 36964 14612
rect 38200 14560 38252 14612
rect 41328 14560 41380 14612
rect 30012 14492 30064 14544
rect 30748 14492 30800 14544
rect 30932 14492 30984 14544
rect 31668 14492 31720 14544
rect 26240 14467 26292 14476
rect 26240 14433 26249 14467
rect 26249 14433 26283 14467
rect 26283 14433 26292 14467
rect 26240 14424 26292 14433
rect 26976 14424 27028 14476
rect 27068 14424 27120 14476
rect 28632 14424 28684 14476
rect 30196 14424 30248 14476
rect 32588 14467 32640 14476
rect 32588 14433 32597 14467
rect 32597 14433 32631 14467
rect 32631 14433 32640 14467
rect 32588 14424 32640 14433
rect 36820 14535 36872 14544
rect 36820 14501 36829 14535
rect 36829 14501 36863 14535
rect 36863 14501 36872 14535
rect 36820 14492 36872 14501
rect 34704 14424 34756 14476
rect 35256 14424 35308 14476
rect 37280 14424 37332 14476
rect 40408 14424 40460 14476
rect 27160 14399 27212 14408
rect 27160 14365 27169 14399
rect 27169 14365 27203 14399
rect 27203 14365 27212 14399
rect 27160 14356 27212 14365
rect 25964 14288 26016 14340
rect 26332 14288 26384 14340
rect 28356 14288 28408 14340
rect 29828 14399 29880 14408
rect 29828 14365 29837 14399
rect 29837 14365 29871 14399
rect 29871 14365 29880 14399
rect 29828 14356 29880 14365
rect 29920 14399 29972 14408
rect 29920 14365 29929 14399
rect 29929 14365 29963 14399
rect 29963 14365 29972 14399
rect 29920 14356 29972 14365
rect 30932 14399 30984 14408
rect 30932 14365 30941 14399
rect 30941 14365 30975 14399
rect 30975 14365 30984 14399
rect 30932 14356 30984 14365
rect 24308 14220 24360 14272
rect 26148 14220 26200 14272
rect 26516 14220 26568 14272
rect 30288 14331 30340 14340
rect 30288 14297 30297 14331
rect 30297 14297 30331 14331
rect 30331 14297 30340 14331
rect 30288 14288 30340 14297
rect 30472 14288 30524 14340
rect 36176 14399 36228 14408
rect 36176 14365 36185 14399
rect 36185 14365 36219 14399
rect 36219 14365 36228 14399
rect 36176 14356 36228 14365
rect 36452 14356 36504 14408
rect 36820 14356 36872 14408
rect 32864 14331 32916 14340
rect 32864 14297 32873 14331
rect 32873 14297 32907 14331
rect 32907 14297 32916 14331
rect 32864 14288 32916 14297
rect 35348 14288 35400 14340
rect 36912 14288 36964 14340
rect 40132 14356 40184 14408
rect 40960 14399 41012 14408
rect 40960 14365 40969 14399
rect 40969 14365 41003 14399
rect 41003 14365 41012 14399
rect 40960 14356 41012 14365
rect 41144 14399 41196 14408
rect 41144 14365 41153 14399
rect 41153 14365 41187 14399
rect 41187 14365 41196 14399
rect 41144 14356 41196 14365
rect 41328 14424 41380 14476
rect 42524 14560 42576 14612
rect 42800 14560 42852 14612
rect 43812 14560 43864 14612
rect 47032 14560 47084 14612
rect 48780 14560 48832 14612
rect 49240 14560 49292 14612
rect 51264 14560 51316 14612
rect 51816 14560 51868 14612
rect 43076 14424 43128 14476
rect 30012 14220 30064 14272
rect 30380 14263 30432 14272
rect 30380 14229 30389 14263
rect 30389 14229 30423 14263
rect 30423 14229 30432 14263
rect 30380 14220 30432 14229
rect 30564 14220 30616 14272
rect 35256 14220 35308 14272
rect 38476 14220 38528 14272
rect 40132 14220 40184 14272
rect 42064 14263 42116 14272
rect 42064 14229 42073 14263
rect 42073 14229 42107 14263
rect 42107 14229 42116 14263
rect 42064 14220 42116 14229
rect 42432 14356 42484 14408
rect 43352 14399 43404 14408
rect 43352 14365 43361 14399
rect 43361 14365 43395 14399
rect 43395 14365 43404 14399
rect 43352 14356 43404 14365
rect 44456 14492 44508 14544
rect 48964 14492 49016 14544
rect 44088 14424 44140 14476
rect 46020 14424 46072 14476
rect 48228 14424 48280 14476
rect 46572 14399 46624 14408
rect 46572 14365 46581 14399
rect 46581 14365 46615 14399
rect 46615 14365 46624 14399
rect 46572 14356 46624 14365
rect 46756 14399 46808 14408
rect 46756 14365 46765 14399
rect 46765 14365 46799 14399
rect 46799 14365 46808 14399
rect 46756 14356 46808 14365
rect 47584 14356 47636 14408
rect 48780 14399 48832 14408
rect 48780 14365 48789 14399
rect 48789 14365 48823 14399
rect 48823 14365 48832 14399
rect 48780 14356 48832 14365
rect 48964 14399 49016 14408
rect 48964 14365 48973 14399
rect 48973 14365 49007 14399
rect 49007 14365 49016 14399
rect 48964 14356 49016 14365
rect 49792 14424 49844 14476
rect 53012 14424 53064 14476
rect 44180 14288 44232 14340
rect 45652 14288 45704 14340
rect 46664 14288 46716 14340
rect 47032 14331 47084 14340
rect 47032 14297 47041 14331
rect 47041 14297 47075 14331
rect 47075 14297 47084 14331
rect 47032 14288 47084 14297
rect 47216 14331 47268 14340
rect 47216 14297 47225 14331
rect 47225 14297 47259 14331
rect 47259 14297 47268 14331
rect 47216 14288 47268 14297
rect 47400 14288 47452 14340
rect 42616 14220 42668 14272
rect 43904 14220 43956 14272
rect 46020 14220 46072 14272
rect 46296 14220 46348 14272
rect 48596 14220 48648 14272
rect 49148 14220 49200 14272
rect 49608 14399 49660 14408
rect 49608 14365 49617 14399
rect 49617 14365 49651 14399
rect 49651 14365 49660 14399
rect 49608 14356 49660 14365
rect 49976 14399 50028 14408
rect 49976 14365 49985 14399
rect 49985 14365 50019 14399
rect 50019 14365 50028 14399
rect 49976 14356 50028 14365
rect 50068 14356 50120 14408
rect 50528 14399 50580 14408
rect 50528 14365 50537 14399
rect 50537 14365 50571 14399
rect 50571 14365 50580 14399
rect 50528 14356 50580 14365
rect 50620 14399 50672 14408
rect 50620 14365 50629 14399
rect 50629 14365 50663 14399
rect 50663 14365 50672 14399
rect 50620 14356 50672 14365
rect 50436 14331 50488 14340
rect 50436 14297 50445 14331
rect 50445 14297 50479 14331
rect 50479 14297 50488 14331
rect 50436 14288 50488 14297
rect 49700 14220 49752 14272
rect 49792 14263 49844 14272
rect 49792 14229 49801 14263
rect 49801 14229 49835 14263
rect 49835 14229 49844 14263
rect 51724 14331 51776 14340
rect 51724 14297 51733 14331
rect 51733 14297 51767 14331
rect 51767 14297 51776 14331
rect 51724 14288 51776 14297
rect 53748 14288 53800 14340
rect 49792 14220 49844 14229
rect 50804 14263 50856 14272
rect 50804 14229 50813 14263
rect 50813 14229 50847 14263
rect 50847 14229 50856 14263
rect 50804 14220 50856 14229
rect 52552 14220 52604 14272
rect 4874 14118 4926 14170
rect 4938 14118 4990 14170
rect 5002 14118 5054 14170
rect 5066 14118 5118 14170
rect 5130 14118 5182 14170
rect 35594 14118 35646 14170
rect 35658 14118 35710 14170
rect 35722 14118 35774 14170
rect 35786 14118 35838 14170
rect 35850 14118 35902 14170
rect 11704 14016 11756 14068
rect 13176 13991 13228 14000
rect 13176 13957 13185 13991
rect 13185 13957 13219 13991
rect 13219 13957 13228 13991
rect 13176 13948 13228 13957
rect 15292 14059 15344 14068
rect 15292 14025 15301 14059
rect 15301 14025 15335 14059
rect 15335 14025 15344 14059
rect 15292 14016 15344 14025
rect 18052 14016 18104 14068
rect 19432 14016 19484 14068
rect 12164 13812 12216 13864
rect 13636 13812 13688 13864
rect 14740 13812 14792 13864
rect 15476 13880 15528 13932
rect 18144 13923 18196 13932
rect 18144 13889 18153 13923
rect 18153 13889 18187 13923
rect 18187 13889 18196 13923
rect 18144 13880 18196 13889
rect 16764 13812 16816 13864
rect 19156 13923 19208 13932
rect 19156 13889 19165 13923
rect 19165 13889 19199 13923
rect 19199 13889 19208 13923
rect 19156 13880 19208 13889
rect 19340 13812 19392 13864
rect 20260 13923 20312 13932
rect 20260 13889 20269 13923
rect 20269 13889 20303 13923
rect 20303 13889 20312 13923
rect 20260 13880 20312 13889
rect 21456 13880 21508 13932
rect 24584 14016 24636 14068
rect 22100 13991 22152 14000
rect 22100 13957 22109 13991
rect 22109 13957 22143 13991
rect 22143 13957 22152 13991
rect 22100 13948 22152 13957
rect 22192 13948 22244 14000
rect 24124 13948 24176 14000
rect 26976 14016 27028 14068
rect 29920 14016 29972 14068
rect 23848 13923 23900 13932
rect 23848 13889 23857 13923
rect 23857 13889 23891 13923
rect 23891 13889 23900 13923
rect 23848 13880 23900 13889
rect 24216 13923 24268 13932
rect 24216 13889 24225 13923
rect 24225 13889 24259 13923
rect 24259 13889 24268 13923
rect 24216 13880 24268 13889
rect 24308 13923 24360 13932
rect 24308 13889 24317 13923
rect 24317 13889 24351 13923
rect 24351 13889 24360 13923
rect 24308 13880 24360 13889
rect 24400 13923 24452 13932
rect 24400 13889 24410 13923
rect 24410 13889 24444 13923
rect 24444 13889 24452 13923
rect 24400 13880 24452 13889
rect 24492 13812 24544 13864
rect 24676 13923 24728 13932
rect 24676 13889 24685 13923
rect 24685 13889 24719 13923
rect 24719 13889 24728 13923
rect 24676 13880 24728 13889
rect 24860 13880 24912 13932
rect 25596 13948 25648 14000
rect 28356 13948 28408 14000
rect 30380 13948 30432 14000
rect 28632 13923 28684 13932
rect 28632 13889 28641 13923
rect 28641 13889 28675 13923
rect 28675 13889 28684 13923
rect 28632 13880 28684 13889
rect 31024 13948 31076 14000
rect 26792 13855 26844 13864
rect 26792 13821 26801 13855
rect 26801 13821 26835 13855
rect 26835 13821 26844 13855
rect 26792 13812 26844 13821
rect 28908 13855 28960 13864
rect 28908 13821 28917 13855
rect 28917 13821 28951 13855
rect 28951 13821 28960 13855
rect 28908 13812 28960 13821
rect 23388 13744 23440 13796
rect 31024 13855 31076 13864
rect 31024 13821 31033 13855
rect 31033 13821 31067 13855
rect 31067 13821 31076 13855
rect 31024 13812 31076 13821
rect 32864 14016 32916 14068
rect 34336 14016 34388 14068
rect 36176 14016 36228 14068
rect 32772 13991 32824 14000
rect 32772 13957 32781 13991
rect 32781 13957 32815 13991
rect 32815 13957 32824 13991
rect 32772 13948 32824 13957
rect 34244 13991 34296 14000
rect 31668 13880 31720 13932
rect 32588 13923 32640 13932
rect 32588 13889 32597 13923
rect 32597 13889 32631 13923
rect 32631 13889 32640 13923
rect 32588 13880 32640 13889
rect 33508 13855 33560 13864
rect 33508 13821 33517 13855
rect 33517 13821 33551 13855
rect 33551 13821 33560 13855
rect 33508 13812 33560 13821
rect 33692 13855 33744 13864
rect 33692 13821 33701 13855
rect 33701 13821 33735 13855
rect 33735 13821 33744 13855
rect 33692 13812 33744 13821
rect 34244 13957 34253 13991
rect 34253 13957 34287 13991
rect 34287 13957 34296 13991
rect 34244 13948 34296 13957
rect 35992 13991 36044 14000
rect 35992 13957 36001 13991
rect 36001 13957 36035 13991
rect 36035 13957 36044 13991
rect 35992 13948 36044 13957
rect 38568 13948 38620 14000
rect 34520 13880 34572 13932
rect 35256 13880 35308 13932
rect 36268 13923 36320 13932
rect 36268 13889 36277 13923
rect 36277 13889 36311 13923
rect 36311 13889 36320 13923
rect 36268 13880 36320 13889
rect 36544 13880 36596 13932
rect 36360 13812 36412 13864
rect 37004 13923 37056 13932
rect 37004 13889 37013 13923
rect 37013 13889 37047 13923
rect 37047 13889 37056 13923
rect 37004 13880 37056 13889
rect 37280 13880 37332 13932
rect 40684 14016 40736 14068
rect 41328 14016 41380 14068
rect 40500 13948 40552 14000
rect 41512 13948 41564 14000
rect 42064 13948 42116 14000
rect 44088 14016 44140 14068
rect 44272 14059 44324 14068
rect 44272 14025 44281 14059
rect 44281 14025 44315 14059
rect 44315 14025 44324 14059
rect 44272 14016 44324 14025
rect 46020 14016 46072 14068
rect 46572 14016 46624 14068
rect 47584 14059 47636 14068
rect 47584 14025 47593 14059
rect 47593 14025 47627 14059
rect 47627 14025 47636 14059
rect 47584 14016 47636 14025
rect 42708 13991 42760 14000
rect 42708 13957 42717 13991
rect 42717 13957 42751 13991
rect 42751 13957 42760 13991
rect 42708 13948 42760 13957
rect 43444 13948 43496 14000
rect 46204 13948 46256 14000
rect 46664 13991 46716 14000
rect 46664 13957 46673 13991
rect 46673 13957 46707 13991
rect 46707 13957 46716 13991
rect 46664 13948 46716 13957
rect 43996 13880 44048 13932
rect 44456 13923 44508 13932
rect 44456 13889 44465 13923
rect 44465 13889 44499 13923
rect 44499 13889 44508 13923
rect 44456 13880 44508 13889
rect 44548 13923 44600 13932
rect 44548 13889 44557 13923
rect 44557 13889 44591 13923
rect 44591 13889 44600 13923
rect 44548 13880 44600 13889
rect 44640 13880 44692 13932
rect 45652 13880 45704 13932
rect 46480 13923 46532 13932
rect 46480 13889 46484 13923
rect 46484 13889 46518 13923
rect 46518 13889 46532 13923
rect 46480 13880 46532 13889
rect 46572 13923 46624 13932
rect 46572 13889 46581 13923
rect 46581 13889 46615 13923
rect 46615 13889 46624 13923
rect 46572 13880 46624 13889
rect 47400 13948 47452 14000
rect 37740 13812 37792 13864
rect 38936 13855 38988 13864
rect 38936 13821 38945 13855
rect 38945 13821 38979 13855
rect 38979 13821 38988 13855
rect 38936 13812 38988 13821
rect 40408 13855 40460 13864
rect 40408 13821 40417 13855
rect 40417 13821 40451 13855
rect 40451 13821 40460 13855
rect 40408 13812 40460 13821
rect 40592 13812 40644 13864
rect 42340 13812 42392 13864
rect 43076 13812 43128 13864
rect 46756 13812 46808 13864
rect 47124 13880 47176 13932
rect 47216 13812 47268 13864
rect 48320 13880 48372 13932
rect 51080 14016 51132 14068
rect 51172 14016 51224 14068
rect 52000 14016 52052 14068
rect 48780 13880 48832 13932
rect 49056 13923 49108 13932
rect 49056 13889 49065 13923
rect 49065 13889 49099 13923
rect 49099 13889 49108 13923
rect 49056 13880 49108 13889
rect 49148 13923 49200 13932
rect 49148 13889 49157 13923
rect 49157 13889 49191 13923
rect 49191 13889 49200 13923
rect 49148 13880 49200 13889
rect 50804 13948 50856 14000
rect 49792 13923 49844 13932
rect 49792 13889 49801 13923
rect 49801 13889 49835 13923
rect 49835 13889 49844 13923
rect 49792 13880 49844 13889
rect 50528 13880 50580 13932
rect 51632 13923 51684 13932
rect 51632 13889 51641 13923
rect 51641 13889 51675 13923
rect 51675 13889 51684 13923
rect 51632 13880 51684 13889
rect 51908 13880 51960 13932
rect 48596 13812 48648 13864
rect 50988 13812 51040 13864
rect 51816 13812 51868 13864
rect 53748 14016 53800 14068
rect 52368 13948 52420 14000
rect 57612 13880 57664 13932
rect 32772 13744 32824 13796
rect 36084 13744 36136 13796
rect 36544 13744 36596 13796
rect 37096 13744 37148 13796
rect 37648 13744 37700 13796
rect 19984 13676 20036 13728
rect 25780 13676 25832 13728
rect 30472 13719 30524 13728
rect 30472 13685 30481 13719
rect 30481 13685 30515 13719
rect 30515 13685 30524 13719
rect 30472 13676 30524 13685
rect 36452 13719 36504 13728
rect 36452 13685 36461 13719
rect 36461 13685 36495 13719
rect 36495 13685 36504 13719
rect 36452 13676 36504 13685
rect 36820 13676 36872 13728
rect 51724 13744 51776 13796
rect 48688 13719 48740 13728
rect 48688 13685 48697 13719
rect 48697 13685 48731 13719
rect 48731 13685 48740 13719
rect 48688 13676 48740 13685
rect 49056 13676 49108 13728
rect 49240 13676 49292 13728
rect 51448 13719 51500 13728
rect 51448 13685 51457 13719
rect 51457 13685 51491 13719
rect 51491 13685 51500 13719
rect 51448 13676 51500 13685
rect 52276 13719 52328 13728
rect 52276 13685 52285 13719
rect 52285 13685 52319 13719
rect 52319 13685 52328 13719
rect 52276 13676 52328 13685
rect 52736 13676 52788 13728
rect 58440 13719 58492 13728
rect 58440 13685 58449 13719
rect 58449 13685 58483 13719
rect 58483 13685 58492 13719
rect 58440 13676 58492 13685
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 13452 13472 13504 13524
rect 12256 13379 12308 13388
rect 12256 13345 12265 13379
rect 12265 13345 12299 13379
rect 12299 13345 12308 13379
rect 12256 13336 12308 13345
rect 12164 13200 12216 13252
rect 13636 13200 13688 13252
rect 15200 13472 15252 13524
rect 24308 13472 24360 13524
rect 28908 13472 28960 13524
rect 32772 13472 32824 13524
rect 35440 13472 35492 13524
rect 36268 13515 36320 13524
rect 36268 13481 36277 13515
rect 36277 13481 36311 13515
rect 36311 13481 36320 13515
rect 36268 13472 36320 13481
rect 36452 13515 36504 13524
rect 36452 13481 36461 13515
rect 36461 13481 36495 13515
rect 36495 13481 36504 13515
rect 36452 13472 36504 13481
rect 36544 13472 36596 13524
rect 27988 13404 28040 13456
rect 29736 13404 29788 13456
rect 29828 13404 29880 13456
rect 14740 13336 14792 13388
rect 14924 13311 14976 13320
rect 14924 13277 14933 13311
rect 14933 13277 14967 13311
rect 14967 13277 14976 13311
rect 14924 13268 14976 13277
rect 15660 13336 15712 13388
rect 16672 13379 16724 13388
rect 16672 13345 16681 13379
rect 16681 13345 16715 13379
rect 16715 13345 16724 13379
rect 16672 13336 16724 13345
rect 17316 13379 17368 13388
rect 17316 13345 17325 13379
rect 17325 13345 17359 13379
rect 17359 13345 17368 13379
rect 17316 13336 17368 13345
rect 17960 13336 18012 13388
rect 16580 13268 16632 13320
rect 16856 13268 16908 13320
rect 17040 13311 17092 13320
rect 17040 13277 17049 13311
rect 17049 13277 17083 13311
rect 17083 13277 17092 13311
rect 17040 13268 17092 13277
rect 17224 13311 17276 13320
rect 17224 13277 17233 13311
rect 17233 13277 17267 13311
rect 17267 13277 17276 13311
rect 17224 13268 17276 13277
rect 23848 13336 23900 13388
rect 26424 13336 26476 13388
rect 27160 13336 27212 13388
rect 29092 13336 29144 13388
rect 30012 13379 30064 13388
rect 30012 13345 30021 13379
rect 30021 13345 30055 13379
rect 30055 13345 30064 13379
rect 30012 13336 30064 13345
rect 17316 13200 17368 13252
rect 15108 13175 15160 13184
rect 15108 13141 15117 13175
rect 15117 13141 15151 13175
rect 15151 13141 15160 13175
rect 15108 13132 15160 13141
rect 17040 13132 17092 13184
rect 17960 13132 18012 13184
rect 20628 13268 20680 13320
rect 23940 13268 23992 13320
rect 24400 13268 24452 13320
rect 27988 13268 28040 13320
rect 29736 13311 29788 13320
rect 29736 13277 29745 13311
rect 29745 13277 29779 13311
rect 29779 13277 29788 13311
rect 29736 13268 29788 13277
rect 29644 13200 29696 13252
rect 30472 13268 30524 13320
rect 30932 13268 30984 13320
rect 31116 13311 31168 13320
rect 31116 13277 31125 13311
rect 31125 13277 31159 13311
rect 31159 13277 31168 13311
rect 31116 13268 31168 13277
rect 32312 13311 32364 13320
rect 32312 13277 32321 13311
rect 32321 13277 32355 13311
rect 32355 13277 32364 13311
rect 32312 13268 32364 13277
rect 37188 13404 37240 13456
rect 37648 13515 37700 13524
rect 37648 13481 37657 13515
rect 37657 13481 37691 13515
rect 37691 13481 37700 13515
rect 37648 13472 37700 13481
rect 37740 13515 37792 13524
rect 37740 13481 37749 13515
rect 37749 13481 37783 13515
rect 37783 13481 37792 13515
rect 37740 13472 37792 13481
rect 38936 13472 38988 13524
rect 41052 13515 41104 13524
rect 41052 13481 41061 13515
rect 41061 13481 41095 13515
rect 41095 13481 41104 13515
rect 41052 13472 41104 13481
rect 41512 13472 41564 13524
rect 42432 13472 42484 13524
rect 45376 13472 45428 13524
rect 48504 13515 48556 13524
rect 48504 13481 48513 13515
rect 48513 13481 48547 13515
rect 48547 13481 48556 13515
rect 48504 13472 48556 13481
rect 48780 13515 48832 13524
rect 48780 13481 48789 13515
rect 48789 13481 48823 13515
rect 48823 13481 48832 13515
rect 48780 13472 48832 13481
rect 51908 13515 51960 13524
rect 51908 13481 51917 13515
rect 51917 13481 51951 13515
rect 51951 13481 51960 13515
rect 51908 13472 51960 13481
rect 52000 13515 52052 13524
rect 52000 13481 52009 13515
rect 52009 13481 52043 13515
rect 52043 13481 52052 13515
rect 52000 13472 52052 13481
rect 54944 13515 54996 13524
rect 54944 13481 54953 13515
rect 54953 13481 54987 13515
rect 54987 13481 54996 13515
rect 54944 13472 54996 13481
rect 33324 13268 33376 13320
rect 36084 13311 36136 13320
rect 36084 13277 36093 13311
rect 36093 13277 36127 13311
rect 36127 13277 36136 13311
rect 36084 13268 36136 13277
rect 36636 13336 36688 13388
rect 36452 13311 36504 13320
rect 36452 13277 36461 13311
rect 36461 13277 36495 13311
rect 36495 13277 36504 13311
rect 36452 13268 36504 13277
rect 36544 13311 36596 13320
rect 36544 13277 36553 13311
rect 36553 13277 36587 13311
rect 36587 13277 36596 13311
rect 36544 13268 36596 13277
rect 32588 13200 32640 13252
rect 33968 13200 34020 13252
rect 36912 13243 36964 13252
rect 36912 13209 36921 13243
rect 36921 13209 36955 13243
rect 36955 13209 36964 13243
rect 36912 13200 36964 13209
rect 37096 13379 37148 13388
rect 37096 13345 37105 13379
rect 37105 13345 37139 13379
rect 37139 13345 37148 13379
rect 37096 13336 37148 13345
rect 37832 13404 37884 13456
rect 38476 13404 38528 13456
rect 40040 13404 40092 13456
rect 51724 13404 51776 13456
rect 40132 13336 40184 13388
rect 40684 13336 40736 13388
rect 44916 13336 44968 13388
rect 46296 13379 46348 13388
rect 46296 13345 46305 13379
rect 46305 13345 46339 13379
rect 46339 13345 46348 13379
rect 46296 13336 46348 13345
rect 46848 13336 46900 13388
rect 37648 13268 37700 13320
rect 37464 13243 37516 13252
rect 37464 13209 37473 13243
rect 37473 13209 37507 13243
rect 37507 13209 37516 13243
rect 37464 13200 37516 13209
rect 37924 13243 37976 13252
rect 37924 13209 37933 13243
rect 37933 13209 37967 13243
rect 37967 13209 37976 13243
rect 37924 13200 37976 13209
rect 38568 13268 38620 13320
rect 39764 13268 39816 13320
rect 41052 13268 41104 13320
rect 44456 13268 44508 13320
rect 40316 13200 40368 13252
rect 41512 13200 41564 13252
rect 19248 13175 19300 13184
rect 19248 13141 19257 13175
rect 19257 13141 19291 13175
rect 19291 13141 19300 13175
rect 19248 13132 19300 13141
rect 26516 13132 26568 13184
rect 30380 13132 30432 13184
rect 31668 13132 31720 13184
rect 36544 13132 36596 13184
rect 37556 13132 37608 13184
rect 39212 13175 39264 13184
rect 39212 13141 39221 13175
rect 39221 13141 39255 13175
rect 39255 13141 39264 13175
rect 39212 13132 39264 13141
rect 45468 13132 45520 13184
rect 45928 13311 45980 13320
rect 45928 13277 45937 13311
rect 45937 13277 45971 13311
rect 45971 13277 45980 13311
rect 45928 13268 45980 13277
rect 48320 13336 48372 13388
rect 49792 13379 49844 13388
rect 49792 13345 49801 13379
rect 49801 13345 49835 13379
rect 49835 13345 49844 13379
rect 49792 13336 49844 13345
rect 51448 13336 51500 13388
rect 48136 13311 48188 13320
rect 48136 13277 48145 13311
rect 48145 13277 48179 13311
rect 48179 13277 48188 13311
rect 48136 13268 48188 13277
rect 48228 13311 48280 13320
rect 48228 13277 48237 13311
rect 48237 13277 48271 13311
rect 48271 13277 48280 13311
rect 48228 13268 48280 13277
rect 48688 13268 48740 13320
rect 55128 13336 55180 13388
rect 47308 13200 47360 13252
rect 48504 13200 48556 13252
rect 50160 13200 50212 13252
rect 55680 13200 55732 13252
rect 56784 13200 56836 13252
rect 52276 13132 52328 13184
rect 57428 13132 57480 13184
rect 4874 13030 4926 13082
rect 4938 13030 4990 13082
rect 5002 13030 5054 13082
rect 5066 13030 5118 13082
rect 5130 13030 5182 13082
rect 35594 13030 35646 13082
rect 35658 13030 35710 13082
rect 35722 13030 35774 13082
rect 35786 13030 35838 13082
rect 35850 13030 35902 13082
rect 16580 12928 16632 12980
rect 16856 12971 16908 12980
rect 16856 12937 16865 12971
rect 16865 12937 16899 12971
rect 16899 12937 16908 12971
rect 16856 12928 16908 12937
rect 17224 12928 17276 12980
rect 24400 12928 24452 12980
rect 24584 12928 24636 12980
rect 18420 12903 18472 12912
rect 15384 12792 15436 12844
rect 17316 12792 17368 12844
rect 18420 12869 18429 12903
rect 18429 12869 18463 12903
rect 18463 12869 18472 12903
rect 18420 12860 18472 12869
rect 19248 12860 19300 12912
rect 24216 12860 24268 12912
rect 16672 12724 16724 12776
rect 19800 12835 19852 12844
rect 19800 12801 19809 12835
rect 19809 12801 19843 12835
rect 19843 12801 19852 12835
rect 19800 12792 19852 12801
rect 21088 12767 21140 12776
rect 21088 12733 21097 12767
rect 21097 12733 21131 12767
rect 21131 12733 21140 12767
rect 21088 12724 21140 12733
rect 25596 12971 25648 12980
rect 25596 12937 25605 12971
rect 25605 12937 25639 12971
rect 25639 12937 25648 12971
rect 25596 12928 25648 12937
rect 26516 12971 26568 12980
rect 26516 12937 26525 12971
rect 26525 12937 26559 12971
rect 26559 12937 26568 12971
rect 26516 12928 26568 12937
rect 27620 12971 27672 12980
rect 27620 12937 27629 12971
rect 27629 12937 27663 12971
rect 27663 12937 27672 12971
rect 27620 12928 27672 12937
rect 26148 12860 26200 12912
rect 25780 12835 25832 12844
rect 25780 12801 25789 12835
rect 25789 12801 25823 12835
rect 25823 12801 25832 12835
rect 25780 12792 25832 12801
rect 25964 12835 26016 12844
rect 25964 12801 25973 12835
rect 25973 12801 26007 12835
rect 26007 12801 26016 12835
rect 25964 12792 26016 12801
rect 26332 12835 26384 12844
rect 26332 12801 26341 12835
rect 26341 12801 26375 12835
rect 26375 12801 26384 12835
rect 26332 12792 26384 12801
rect 24768 12724 24820 12776
rect 26792 12724 26844 12776
rect 30012 12928 30064 12980
rect 31116 12928 31168 12980
rect 32220 12928 32272 12980
rect 33048 12928 33100 12980
rect 33508 12971 33560 12980
rect 33508 12937 33517 12971
rect 33517 12937 33551 12971
rect 33551 12937 33560 12971
rect 33508 12928 33560 12937
rect 36636 12971 36688 12980
rect 36636 12937 36645 12971
rect 36645 12937 36679 12971
rect 36679 12937 36688 12971
rect 36636 12928 36688 12937
rect 37740 12928 37792 12980
rect 38568 12971 38620 12980
rect 38568 12937 38577 12971
rect 38577 12937 38611 12971
rect 38611 12937 38620 12971
rect 38568 12928 38620 12937
rect 39212 12928 39264 12980
rect 29000 12835 29052 12844
rect 29000 12801 29009 12835
rect 29009 12801 29043 12835
rect 29043 12801 29052 12835
rect 29000 12792 29052 12801
rect 29368 12792 29420 12844
rect 29644 12835 29696 12844
rect 29644 12801 29653 12835
rect 29653 12801 29687 12835
rect 29687 12801 29696 12835
rect 29644 12792 29696 12801
rect 29184 12724 29236 12776
rect 30288 12724 30340 12776
rect 32588 12835 32640 12844
rect 32588 12801 32597 12835
rect 32597 12801 32631 12835
rect 32631 12801 32640 12835
rect 32588 12792 32640 12801
rect 33416 12860 33468 12912
rect 33508 12792 33560 12844
rect 36268 12792 36320 12844
rect 36820 12835 36872 12844
rect 36820 12801 36829 12835
rect 36829 12801 36863 12835
rect 36863 12801 36872 12835
rect 36820 12792 36872 12801
rect 37004 12835 37056 12844
rect 37004 12801 37013 12835
rect 37013 12801 37047 12835
rect 37047 12801 37056 12835
rect 37004 12792 37056 12801
rect 26608 12656 26660 12708
rect 29552 12656 29604 12708
rect 33140 12724 33192 12776
rect 37096 12724 37148 12776
rect 37648 12835 37700 12844
rect 37648 12801 37657 12835
rect 37657 12801 37691 12835
rect 37691 12801 37700 12835
rect 37648 12792 37700 12801
rect 38476 12835 38528 12844
rect 38476 12801 38485 12835
rect 38485 12801 38519 12835
rect 38519 12801 38528 12835
rect 38476 12792 38528 12801
rect 38752 12835 38804 12844
rect 38752 12801 38761 12835
rect 38761 12801 38795 12835
rect 38795 12801 38804 12835
rect 38752 12792 38804 12801
rect 38844 12835 38896 12844
rect 38844 12801 38853 12835
rect 38853 12801 38887 12835
rect 38887 12801 38896 12835
rect 38844 12792 38896 12801
rect 40592 12860 40644 12912
rect 45468 12903 45520 12912
rect 45468 12869 45477 12903
rect 45477 12869 45511 12903
rect 45511 12869 45520 12903
rect 45468 12860 45520 12869
rect 46756 12860 46808 12912
rect 47308 12860 47360 12912
rect 37740 12724 37792 12776
rect 38660 12767 38712 12776
rect 38660 12733 38669 12767
rect 38669 12733 38703 12767
rect 38703 12733 38712 12767
rect 38660 12724 38712 12733
rect 39120 12724 39172 12776
rect 39304 12792 39356 12844
rect 39580 12792 39632 12844
rect 44916 12792 44968 12844
rect 49792 12928 49844 12980
rect 50528 12971 50580 12980
rect 50528 12937 50537 12971
rect 50537 12937 50571 12971
rect 50571 12937 50580 12971
rect 50528 12928 50580 12937
rect 57612 12971 57664 12980
rect 57612 12937 57621 12971
rect 57621 12937 57655 12971
rect 57655 12937 57664 12971
rect 57612 12928 57664 12937
rect 49056 12903 49108 12912
rect 49056 12869 49065 12903
rect 49065 12869 49099 12903
rect 49099 12869 49108 12903
rect 49056 12860 49108 12869
rect 33048 12656 33100 12708
rect 33692 12656 33744 12708
rect 19616 12631 19668 12640
rect 19616 12597 19625 12631
rect 19625 12597 19659 12631
rect 19659 12597 19668 12631
rect 19616 12588 19668 12597
rect 19708 12588 19760 12640
rect 27252 12631 27304 12640
rect 27252 12597 27261 12631
rect 27261 12597 27295 12631
rect 27295 12597 27304 12631
rect 27252 12588 27304 12597
rect 30472 12588 30524 12640
rect 33232 12588 33284 12640
rect 37924 12656 37976 12708
rect 39948 12724 40000 12776
rect 42892 12767 42944 12776
rect 42892 12733 42901 12767
rect 42901 12733 42935 12767
rect 42935 12733 42944 12767
rect 42892 12724 42944 12733
rect 39764 12656 39816 12708
rect 44272 12767 44324 12776
rect 44272 12733 44281 12767
rect 44281 12733 44315 12767
rect 44315 12733 44324 12767
rect 44272 12724 44324 12733
rect 48136 12724 48188 12776
rect 50160 12792 50212 12844
rect 57428 12835 57480 12844
rect 57428 12801 57437 12835
rect 57437 12801 57471 12835
rect 57471 12801 57480 12835
rect 57428 12792 57480 12801
rect 42800 12588 42852 12640
rect 45928 12588 45980 12640
rect 46572 12588 46624 12640
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 12164 12291 12216 12300
rect 12164 12257 12173 12291
rect 12173 12257 12207 12291
rect 12207 12257 12216 12291
rect 15384 12384 15436 12436
rect 17040 12384 17092 12436
rect 12164 12248 12216 12257
rect 14740 12291 14792 12300
rect 14740 12257 14749 12291
rect 14749 12257 14783 12291
rect 14783 12257 14792 12291
rect 14740 12248 14792 12257
rect 15660 12291 15712 12300
rect 15660 12257 15669 12291
rect 15669 12257 15703 12291
rect 15703 12257 15712 12291
rect 15660 12248 15712 12257
rect 17960 12316 18012 12368
rect 14832 12223 14884 12232
rect 14832 12189 14841 12223
rect 14841 12189 14875 12223
rect 14875 12189 14884 12223
rect 14832 12180 14884 12189
rect 15292 12180 15344 12232
rect 16764 12180 16816 12232
rect 13452 12112 13504 12164
rect 16948 12112 17000 12164
rect 19800 12384 19852 12436
rect 24860 12384 24912 12436
rect 19248 12316 19300 12368
rect 26332 12316 26384 12368
rect 26792 12384 26844 12436
rect 27988 12427 28040 12436
rect 27988 12393 27997 12427
rect 27997 12393 28031 12427
rect 28031 12393 28040 12427
rect 27988 12384 28040 12393
rect 29000 12384 29052 12436
rect 29736 12384 29788 12436
rect 26884 12316 26936 12368
rect 31668 12427 31720 12436
rect 31668 12393 31677 12427
rect 31677 12393 31711 12427
rect 31711 12393 31720 12427
rect 31668 12384 31720 12393
rect 32588 12384 32640 12436
rect 33140 12384 33192 12436
rect 33784 12384 33836 12436
rect 35716 12384 35768 12436
rect 37648 12384 37700 12436
rect 37740 12384 37792 12436
rect 39672 12384 39724 12436
rect 40868 12384 40920 12436
rect 43720 12384 43772 12436
rect 46204 12427 46256 12436
rect 46204 12393 46213 12427
rect 46213 12393 46247 12427
rect 46247 12393 46256 12427
rect 46204 12384 46256 12393
rect 46756 12384 46808 12436
rect 18420 12180 18472 12232
rect 19248 12223 19300 12232
rect 19248 12189 19257 12223
rect 19257 12189 19291 12223
rect 19291 12189 19300 12223
rect 19248 12180 19300 12189
rect 24584 12291 24636 12300
rect 24584 12257 24593 12291
rect 24593 12257 24627 12291
rect 24627 12257 24636 12291
rect 24584 12248 24636 12257
rect 26700 12248 26752 12300
rect 27344 12248 27396 12300
rect 19708 12180 19760 12232
rect 26608 12180 26660 12232
rect 14096 12087 14148 12096
rect 14096 12053 14105 12087
rect 14105 12053 14139 12087
rect 14139 12053 14148 12087
rect 14096 12044 14148 12053
rect 15292 12044 15344 12096
rect 17500 12087 17552 12096
rect 17500 12053 17509 12087
rect 17509 12053 17543 12087
rect 17543 12053 17552 12087
rect 17500 12044 17552 12053
rect 17868 12087 17920 12096
rect 17868 12053 17877 12087
rect 17877 12053 17911 12087
rect 17911 12053 17920 12087
rect 17868 12044 17920 12053
rect 20904 12044 20956 12096
rect 22192 12112 22244 12164
rect 27160 12223 27212 12232
rect 27160 12189 27169 12223
rect 27169 12189 27203 12223
rect 27203 12189 27212 12223
rect 27160 12180 27212 12189
rect 28724 12180 28776 12232
rect 28908 12223 28960 12232
rect 28908 12189 28917 12223
rect 28917 12189 28951 12223
rect 28951 12189 28960 12223
rect 28908 12180 28960 12189
rect 32680 12316 32732 12368
rect 24768 12044 24820 12096
rect 30380 12180 30432 12232
rect 30472 12223 30524 12232
rect 30472 12189 30481 12223
rect 30481 12189 30515 12223
rect 30515 12189 30524 12223
rect 30472 12180 30524 12189
rect 30564 12223 30616 12232
rect 30564 12189 30573 12223
rect 30573 12189 30607 12223
rect 30607 12189 30616 12223
rect 30564 12180 30616 12189
rect 29920 12112 29972 12164
rect 31484 12223 31536 12232
rect 31484 12189 31493 12223
rect 31493 12189 31527 12223
rect 31527 12189 31536 12223
rect 31484 12180 31536 12189
rect 31760 12223 31812 12232
rect 31760 12189 31769 12223
rect 31769 12189 31803 12223
rect 31803 12189 31812 12223
rect 31760 12180 31812 12189
rect 33048 12223 33100 12232
rect 33048 12189 33057 12223
rect 33057 12189 33091 12223
rect 33091 12189 33100 12223
rect 33048 12180 33100 12189
rect 38660 12316 38712 12368
rect 34244 12291 34296 12300
rect 34244 12257 34253 12291
rect 34253 12257 34287 12291
rect 34287 12257 34296 12291
rect 34244 12248 34296 12257
rect 33324 12180 33376 12232
rect 33692 12223 33744 12232
rect 33692 12189 33701 12223
rect 33701 12189 33735 12223
rect 33735 12189 33744 12223
rect 33692 12180 33744 12189
rect 33784 12223 33836 12232
rect 33784 12189 33793 12223
rect 33793 12189 33827 12223
rect 33827 12189 33836 12223
rect 33784 12180 33836 12189
rect 26240 12044 26292 12096
rect 26884 12044 26936 12096
rect 26976 12044 27028 12096
rect 27620 12044 27672 12096
rect 29460 12044 29512 12096
rect 30288 12044 30340 12096
rect 31024 12112 31076 12164
rect 33968 12223 34020 12232
rect 33968 12189 33977 12223
rect 33977 12189 34011 12223
rect 34011 12189 34020 12223
rect 33968 12180 34020 12189
rect 34428 12180 34480 12232
rect 34888 12223 34940 12232
rect 34888 12189 34897 12223
rect 34897 12189 34931 12223
rect 34931 12189 34940 12223
rect 34888 12180 34940 12189
rect 35164 12223 35216 12232
rect 35164 12189 35173 12223
rect 35173 12189 35207 12223
rect 35207 12189 35216 12223
rect 35164 12180 35216 12189
rect 35440 12180 35492 12232
rect 35716 12223 35768 12232
rect 35716 12189 35720 12223
rect 35720 12189 35754 12223
rect 35754 12189 35768 12223
rect 35716 12180 35768 12189
rect 35992 12180 36044 12232
rect 32588 12044 32640 12096
rect 35348 12044 35400 12096
rect 36268 12112 36320 12164
rect 37832 12180 37884 12232
rect 38752 12180 38804 12232
rect 39212 12223 39264 12232
rect 39212 12189 39221 12223
rect 39221 12189 39255 12223
rect 39255 12189 39264 12223
rect 39212 12180 39264 12189
rect 39488 12180 39540 12232
rect 39948 12223 40000 12232
rect 39948 12189 39958 12223
rect 39958 12189 39992 12223
rect 39992 12189 40000 12223
rect 39948 12180 40000 12189
rect 40316 12223 40368 12232
rect 40316 12189 40330 12223
rect 40330 12189 40364 12223
rect 40364 12189 40368 12223
rect 40316 12180 40368 12189
rect 40592 12223 40644 12232
rect 40592 12189 40601 12223
rect 40601 12189 40635 12223
rect 40635 12189 40644 12223
rect 40592 12180 40644 12189
rect 40868 12223 40920 12232
rect 40868 12189 40877 12223
rect 40877 12189 40911 12223
rect 40911 12189 40920 12223
rect 40868 12180 40920 12189
rect 40960 12223 41012 12232
rect 40960 12189 40969 12223
rect 40969 12189 41003 12223
rect 41003 12189 41012 12223
rect 40960 12180 41012 12189
rect 35992 12044 36044 12096
rect 36452 12044 36504 12096
rect 37740 12044 37792 12096
rect 38660 12044 38712 12096
rect 38844 12087 38896 12096
rect 38844 12053 38853 12087
rect 38853 12053 38887 12087
rect 38887 12053 38896 12087
rect 38844 12044 38896 12053
rect 39396 12044 39448 12096
rect 39672 12112 39724 12164
rect 40776 12155 40828 12164
rect 40776 12121 40785 12155
rect 40785 12121 40819 12155
rect 40819 12121 40828 12155
rect 40776 12112 40828 12121
rect 40684 12044 40736 12096
rect 41328 12248 41380 12300
rect 45928 12248 45980 12300
rect 46204 12180 46256 12232
rect 42432 12112 42484 12164
rect 4874 11942 4926 11994
rect 4938 11942 4990 11994
rect 5002 11942 5054 11994
rect 5066 11942 5118 11994
rect 5130 11942 5182 11994
rect 35594 11942 35646 11994
rect 35658 11942 35710 11994
rect 35722 11942 35774 11994
rect 35786 11942 35838 11994
rect 35850 11942 35902 11994
rect 17500 11840 17552 11892
rect 19248 11840 19300 11892
rect 26700 11840 26752 11892
rect 27252 11840 27304 11892
rect 29552 11883 29604 11892
rect 29552 11849 29561 11883
rect 29561 11849 29595 11883
rect 29595 11849 29604 11883
rect 29552 11840 29604 11849
rect 13452 11772 13504 11824
rect 19616 11772 19668 11824
rect 22192 11772 22244 11824
rect 12164 11747 12216 11756
rect 12164 11713 12173 11747
rect 12173 11713 12207 11747
rect 12207 11713 12216 11747
rect 12164 11704 12216 11713
rect 14740 11747 14792 11756
rect 14740 11713 14749 11747
rect 14749 11713 14783 11747
rect 14783 11713 14792 11747
rect 14740 11704 14792 11713
rect 12440 11679 12492 11688
rect 12440 11645 12449 11679
rect 12449 11645 12483 11679
rect 12483 11645 12492 11679
rect 12440 11636 12492 11645
rect 14280 11636 14332 11688
rect 17316 11704 17368 11756
rect 26700 11704 26752 11756
rect 21088 11636 21140 11688
rect 22468 11636 22520 11688
rect 28356 11704 28408 11756
rect 28816 11747 28868 11756
rect 28816 11713 28825 11747
rect 28825 11713 28859 11747
rect 28859 11713 28868 11747
rect 28816 11704 28868 11713
rect 29276 11636 29328 11688
rect 29552 11704 29604 11756
rect 29736 11747 29788 11756
rect 29736 11713 29740 11747
rect 29740 11713 29774 11747
rect 29774 11713 29788 11747
rect 29736 11704 29788 11713
rect 30380 11772 30432 11824
rect 29644 11568 29696 11620
rect 30196 11747 30248 11756
rect 30196 11713 30205 11747
rect 30205 11713 30239 11747
rect 30239 11713 30248 11747
rect 30196 11704 30248 11713
rect 31024 11815 31076 11824
rect 31024 11781 31033 11815
rect 31033 11781 31067 11815
rect 31067 11781 31076 11815
rect 31024 11772 31076 11781
rect 31116 11815 31168 11824
rect 31116 11781 31151 11815
rect 31151 11781 31168 11815
rect 32496 11840 32548 11892
rect 33232 11883 33284 11892
rect 33232 11849 33241 11883
rect 33241 11849 33275 11883
rect 33275 11849 33284 11883
rect 33232 11840 33284 11849
rect 33324 11883 33376 11892
rect 33324 11849 33333 11883
rect 33333 11849 33367 11883
rect 33367 11849 33376 11883
rect 33324 11840 33376 11849
rect 34888 11840 34940 11892
rect 35072 11840 35124 11892
rect 35256 11840 35308 11892
rect 37556 11840 37608 11892
rect 38384 11840 38436 11892
rect 39396 11883 39448 11892
rect 39396 11849 39405 11883
rect 39405 11849 39439 11883
rect 39439 11849 39448 11883
rect 39396 11840 39448 11849
rect 40776 11840 40828 11892
rect 42432 11840 42484 11892
rect 31116 11772 31168 11781
rect 35992 11815 36044 11824
rect 35992 11781 36001 11815
rect 36001 11781 36035 11815
rect 36035 11781 36044 11815
rect 35992 11772 36044 11781
rect 36084 11772 36136 11824
rect 30748 11636 30800 11688
rect 32312 11704 32364 11756
rect 32588 11747 32640 11756
rect 32588 11713 32597 11747
rect 32597 11713 32631 11747
rect 32631 11713 32640 11747
rect 32588 11704 32640 11713
rect 32772 11747 32824 11756
rect 32772 11713 32779 11747
rect 32779 11713 32824 11747
rect 32772 11704 32824 11713
rect 32864 11747 32916 11756
rect 32864 11713 32873 11747
rect 32873 11713 32907 11747
rect 32907 11713 32916 11747
rect 32864 11704 32916 11713
rect 33048 11747 33100 11756
rect 33048 11713 33062 11747
rect 33062 11713 33096 11747
rect 33096 11713 33100 11747
rect 33048 11704 33100 11713
rect 33324 11747 33376 11756
rect 33324 11713 33333 11747
rect 33333 11713 33367 11747
rect 33367 11713 33376 11747
rect 33324 11704 33376 11713
rect 33600 11747 33652 11756
rect 33600 11713 33609 11747
rect 33609 11713 33643 11747
rect 33643 11713 33652 11747
rect 33600 11704 33652 11713
rect 33784 11747 33836 11756
rect 33784 11713 33793 11747
rect 33793 11713 33827 11747
rect 33827 11713 33836 11747
rect 33784 11704 33836 11713
rect 34612 11704 34664 11756
rect 35256 11704 35308 11756
rect 31484 11568 31536 11620
rect 32680 11568 32732 11620
rect 35348 11636 35400 11688
rect 36268 11747 36320 11756
rect 36268 11713 36277 11747
rect 36277 11713 36311 11747
rect 36311 11713 36320 11747
rect 36268 11704 36320 11713
rect 36544 11704 36596 11756
rect 36636 11704 36688 11756
rect 37740 11704 37792 11756
rect 37924 11704 37976 11756
rect 38292 11747 38344 11756
rect 38292 11713 38298 11747
rect 38298 11713 38332 11747
rect 38332 11713 38344 11747
rect 38292 11704 38344 11713
rect 40040 11772 40092 11824
rect 40960 11772 41012 11824
rect 42800 11815 42852 11824
rect 42800 11781 42809 11815
rect 42809 11781 42843 11815
rect 42843 11781 42852 11815
rect 42800 11772 42852 11781
rect 44272 11883 44324 11892
rect 44272 11849 44281 11883
rect 44281 11849 44315 11883
rect 44315 11849 44324 11883
rect 44272 11840 44324 11849
rect 38476 11704 38528 11756
rect 38752 11704 38804 11756
rect 38936 11747 38988 11756
rect 38936 11713 38946 11747
rect 38946 11713 38980 11747
rect 38980 11713 38988 11747
rect 38936 11704 38988 11713
rect 14004 11543 14056 11552
rect 14004 11509 14013 11543
rect 14013 11509 14047 11543
rect 14047 11509 14056 11543
rect 14004 11500 14056 11509
rect 15476 11500 15528 11552
rect 16396 11500 16448 11552
rect 20168 11500 20220 11552
rect 22008 11500 22060 11552
rect 27620 11500 27672 11552
rect 27988 11500 28040 11552
rect 28724 11500 28776 11552
rect 29184 11543 29236 11552
rect 29184 11509 29193 11543
rect 29193 11509 29227 11543
rect 29227 11509 29236 11543
rect 29184 11500 29236 11509
rect 30472 11500 30524 11552
rect 30932 11500 30984 11552
rect 33416 11500 33468 11552
rect 34336 11500 34388 11552
rect 35348 11500 35400 11552
rect 36268 11568 36320 11620
rect 39028 11679 39080 11688
rect 39028 11645 39037 11679
rect 39037 11645 39071 11679
rect 39071 11645 39080 11679
rect 39028 11636 39080 11645
rect 39120 11679 39172 11688
rect 39120 11645 39129 11679
rect 39129 11645 39163 11679
rect 39163 11645 39172 11679
rect 39120 11636 39172 11645
rect 39672 11636 39724 11688
rect 39856 11747 39908 11756
rect 39856 11713 39865 11747
rect 39865 11713 39899 11747
rect 39899 11713 39908 11747
rect 39856 11704 39908 11713
rect 39948 11747 40000 11756
rect 39948 11713 39957 11747
rect 39957 11713 39991 11747
rect 39991 11713 40000 11747
rect 39948 11704 40000 11713
rect 41328 11704 41380 11756
rect 36636 11500 36688 11552
rect 37832 11500 37884 11552
rect 40592 11568 40644 11620
rect 39028 11500 39080 11552
rect 39212 11500 39264 11552
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 12440 11296 12492 11348
rect 14832 11296 14884 11348
rect 15660 11296 15712 11348
rect 16396 11339 16448 11348
rect 16396 11305 16405 11339
rect 16405 11305 16439 11339
rect 16439 11305 16448 11339
rect 16396 11296 16448 11305
rect 16672 11296 16724 11348
rect 22468 11339 22520 11348
rect 22468 11305 22477 11339
rect 22477 11305 22511 11339
rect 22511 11305 22520 11339
rect 22468 11296 22520 11305
rect 13544 11160 13596 11212
rect 14004 11092 14056 11144
rect 14096 11135 14148 11144
rect 14096 11101 14105 11135
rect 14105 11101 14139 11135
rect 14139 11101 14148 11135
rect 14096 11092 14148 11101
rect 14280 11135 14332 11144
rect 14280 11101 14289 11135
rect 14289 11101 14323 11135
rect 14323 11101 14332 11135
rect 14280 11092 14332 11101
rect 14740 11160 14792 11212
rect 15292 11271 15344 11280
rect 15292 11237 15301 11271
rect 15301 11237 15335 11271
rect 15335 11237 15344 11271
rect 15292 11228 15344 11237
rect 17224 11228 17276 11280
rect 18236 11228 18288 11280
rect 15476 11135 15528 11144
rect 15476 11101 15485 11135
rect 15485 11101 15519 11135
rect 15519 11101 15528 11135
rect 15476 11092 15528 11101
rect 15844 11067 15896 11076
rect 15844 11033 15853 11067
rect 15853 11033 15887 11067
rect 15887 11033 15896 11067
rect 15844 11024 15896 11033
rect 16028 11092 16080 11144
rect 17868 11160 17920 11212
rect 16948 11135 17000 11144
rect 16948 11101 16957 11135
rect 16957 11101 16991 11135
rect 16991 11101 17000 11135
rect 16948 11092 17000 11101
rect 17316 11135 17368 11144
rect 17316 11101 17325 11135
rect 17325 11101 17359 11135
rect 17359 11101 17368 11135
rect 17316 11092 17368 11101
rect 22560 11228 22612 11280
rect 28540 11228 28592 11280
rect 28908 11339 28960 11348
rect 28908 11305 28917 11339
rect 28917 11305 28951 11339
rect 28951 11305 28960 11339
rect 28908 11296 28960 11305
rect 29828 11296 29880 11348
rect 30564 11296 30616 11348
rect 33324 11296 33376 11348
rect 36452 11296 36504 11348
rect 37924 11296 37976 11348
rect 38660 11296 38712 11348
rect 39120 11339 39172 11348
rect 39120 11305 39129 11339
rect 39129 11305 39163 11339
rect 39163 11305 39172 11339
rect 39120 11296 39172 11305
rect 39212 11296 39264 11348
rect 29920 11228 29972 11280
rect 30380 11228 30432 11280
rect 32864 11228 32916 11280
rect 35440 11271 35492 11280
rect 35440 11237 35449 11271
rect 35449 11237 35483 11271
rect 35483 11237 35492 11271
rect 35440 11228 35492 11237
rect 37832 11228 37884 11280
rect 39856 11296 39908 11348
rect 21364 11160 21416 11212
rect 29276 11160 29328 11212
rect 19892 11135 19944 11144
rect 19892 11101 19901 11135
rect 19901 11101 19935 11135
rect 19935 11101 19944 11135
rect 19892 11092 19944 11101
rect 15568 10999 15620 11008
rect 15568 10965 15577 10999
rect 15577 10965 15611 10999
rect 15611 10965 15620 10999
rect 15568 10956 15620 10965
rect 15660 10999 15712 11008
rect 15660 10965 15669 10999
rect 15669 10965 15703 10999
rect 15703 10965 15712 10999
rect 15660 10956 15712 10965
rect 17132 10999 17184 11008
rect 17132 10965 17141 10999
rect 17141 10965 17175 10999
rect 17175 10965 17184 10999
rect 17132 10956 17184 10965
rect 17960 10956 18012 11008
rect 19248 10956 19300 11008
rect 20720 11092 20772 11144
rect 22008 11135 22060 11144
rect 22008 11101 22017 11135
rect 22017 11101 22051 11135
rect 22051 11101 22060 11135
rect 22008 11092 22060 11101
rect 24952 11092 25004 11144
rect 22928 11024 22980 11076
rect 27620 11024 27672 11076
rect 27896 11067 27948 11076
rect 27896 11033 27905 11067
rect 27905 11033 27939 11067
rect 27939 11033 27948 11067
rect 27896 11024 27948 11033
rect 28356 11092 28408 11144
rect 29000 11092 29052 11144
rect 29092 11135 29144 11144
rect 29092 11101 29101 11135
rect 29101 11101 29135 11135
rect 29135 11101 29144 11135
rect 29092 11092 29144 11101
rect 30472 11135 30524 11144
rect 30472 11101 30481 11135
rect 30481 11101 30515 11135
rect 30515 11101 30524 11135
rect 30472 11092 30524 11101
rect 31116 11160 31168 11212
rect 32312 11203 32364 11212
rect 32312 11169 32321 11203
rect 32321 11169 32355 11203
rect 32355 11169 32364 11203
rect 32312 11160 32364 11169
rect 29552 11024 29604 11076
rect 33508 11160 33560 11212
rect 32496 11135 32548 11144
rect 32496 11101 32505 11135
rect 32505 11101 32539 11135
rect 32539 11101 32548 11135
rect 32496 11092 32548 11101
rect 33324 11092 33376 11144
rect 34796 11135 34848 11144
rect 34796 11101 34805 11135
rect 34805 11101 34839 11135
rect 34839 11101 34848 11135
rect 34796 11092 34848 11101
rect 34888 11135 34940 11144
rect 34888 11101 34897 11135
rect 34897 11101 34931 11135
rect 34931 11101 34940 11135
rect 34888 11092 34940 11101
rect 20076 10999 20128 11008
rect 20076 10965 20085 10999
rect 20085 10965 20119 10999
rect 20119 10965 20128 10999
rect 20076 10956 20128 10965
rect 34336 11024 34388 11076
rect 35440 11092 35492 11144
rect 36544 11160 36596 11212
rect 40316 11203 40368 11212
rect 40316 11169 40325 11203
rect 40325 11169 40359 11203
rect 40359 11169 40368 11203
rect 40316 11160 40368 11169
rect 38292 11135 38344 11144
rect 38292 11101 38301 11135
rect 38301 11101 38335 11135
rect 38335 11101 38344 11135
rect 38292 11092 38344 11101
rect 35348 11024 35400 11076
rect 38108 11024 38160 11076
rect 38568 11135 38620 11144
rect 38568 11101 38577 11135
rect 38577 11101 38611 11135
rect 38611 11101 38620 11135
rect 38568 11092 38620 11101
rect 39212 11092 39264 11144
rect 39580 11067 39632 11076
rect 39580 11033 39589 11067
rect 39589 11033 39623 11067
rect 39623 11033 39632 11067
rect 39580 11024 39632 11033
rect 41696 11024 41748 11076
rect 34428 10956 34480 11008
rect 34520 10956 34572 11008
rect 37372 10956 37424 11008
rect 39212 10956 39264 11008
rect 39488 10956 39540 11008
rect 4874 10854 4926 10906
rect 4938 10854 4990 10906
rect 5002 10854 5054 10906
rect 5066 10854 5118 10906
rect 5130 10854 5182 10906
rect 35594 10854 35646 10906
rect 35658 10854 35710 10906
rect 35722 10854 35774 10906
rect 35786 10854 35838 10906
rect 35850 10854 35902 10906
rect 13544 10795 13596 10804
rect 13544 10761 13553 10795
rect 13553 10761 13587 10795
rect 13587 10761 13596 10795
rect 13544 10752 13596 10761
rect 17132 10752 17184 10804
rect 20168 10795 20220 10804
rect 20168 10761 20177 10795
rect 20177 10761 20211 10795
rect 20211 10761 20220 10795
rect 20168 10752 20220 10761
rect 22468 10752 22520 10804
rect 26700 10795 26752 10804
rect 26700 10761 26709 10795
rect 26709 10761 26743 10795
rect 26743 10761 26752 10795
rect 26700 10752 26752 10761
rect 13912 10727 13964 10736
rect 13912 10693 13921 10727
rect 13921 10693 13955 10727
rect 13955 10693 13964 10727
rect 13912 10684 13964 10693
rect 15844 10684 15896 10736
rect 14832 10616 14884 10668
rect 15660 10616 15712 10668
rect 17960 10684 18012 10736
rect 19984 10684 20036 10736
rect 18052 10659 18104 10668
rect 16120 10548 16172 10600
rect 14096 10480 14148 10532
rect 15568 10480 15620 10532
rect 18052 10625 18061 10659
rect 18061 10625 18095 10659
rect 18095 10625 18104 10659
rect 18052 10616 18104 10625
rect 18236 10659 18288 10668
rect 18236 10625 18245 10659
rect 18245 10625 18279 10659
rect 18279 10625 18288 10659
rect 18236 10616 18288 10625
rect 22100 10684 22152 10736
rect 22928 10684 22980 10736
rect 26608 10684 26660 10736
rect 27896 10795 27948 10804
rect 27896 10761 27905 10795
rect 27905 10761 27939 10795
rect 27939 10761 27948 10795
rect 27896 10752 27948 10761
rect 28448 10752 28500 10804
rect 20720 10659 20772 10668
rect 20720 10625 20729 10659
rect 20729 10625 20763 10659
rect 20763 10625 20772 10659
rect 20720 10616 20772 10625
rect 18328 10591 18380 10600
rect 18328 10557 18337 10591
rect 18337 10557 18371 10591
rect 18371 10557 18380 10591
rect 18328 10548 18380 10557
rect 19248 10548 19300 10600
rect 21364 10659 21416 10668
rect 21364 10625 21373 10659
rect 21373 10625 21407 10659
rect 21407 10625 21416 10659
rect 21364 10616 21416 10625
rect 26516 10616 26568 10668
rect 27252 10616 27304 10668
rect 13452 10455 13504 10464
rect 13452 10421 13461 10455
rect 13461 10421 13495 10455
rect 13495 10421 13504 10455
rect 13452 10412 13504 10421
rect 14832 10412 14884 10464
rect 19892 10412 19944 10464
rect 20260 10480 20312 10532
rect 22836 10548 22888 10600
rect 23940 10548 23992 10600
rect 24952 10591 25004 10600
rect 24952 10557 24961 10591
rect 24961 10557 24995 10591
rect 24995 10557 25004 10591
rect 24952 10548 25004 10557
rect 25872 10548 25924 10600
rect 27988 10659 28040 10668
rect 27988 10625 27997 10659
rect 27997 10625 28031 10659
rect 28031 10625 28040 10659
rect 27988 10616 28040 10625
rect 29552 10752 29604 10804
rect 30196 10752 30248 10804
rect 31760 10752 31812 10804
rect 32680 10795 32732 10804
rect 32680 10761 32689 10795
rect 32689 10761 32723 10795
rect 32723 10761 32732 10795
rect 32680 10752 32732 10761
rect 32772 10752 32824 10804
rect 34796 10752 34848 10804
rect 36176 10752 36228 10804
rect 37096 10795 37148 10804
rect 37096 10761 37105 10795
rect 37105 10761 37139 10795
rect 37139 10761 37148 10795
rect 37096 10752 37148 10761
rect 37372 10795 37424 10804
rect 37372 10761 37381 10795
rect 37381 10761 37415 10795
rect 37415 10761 37424 10795
rect 37372 10752 37424 10761
rect 28356 10659 28408 10668
rect 28356 10625 28366 10659
rect 28366 10625 28400 10659
rect 28400 10625 28408 10659
rect 28356 10616 28408 10625
rect 28540 10659 28592 10668
rect 28540 10625 28549 10659
rect 28549 10625 28583 10659
rect 28583 10625 28592 10659
rect 28540 10616 28592 10625
rect 28908 10616 28960 10668
rect 29184 10659 29236 10668
rect 29184 10625 29193 10659
rect 29193 10625 29227 10659
rect 29227 10625 29236 10659
rect 29184 10616 29236 10625
rect 30748 10727 30800 10736
rect 30748 10693 30757 10727
rect 30757 10693 30791 10727
rect 30791 10693 30800 10727
rect 30748 10684 30800 10693
rect 31024 10684 31076 10736
rect 29460 10659 29512 10668
rect 29460 10625 29469 10659
rect 29469 10625 29503 10659
rect 29503 10625 29512 10659
rect 29460 10616 29512 10625
rect 30380 10616 30432 10668
rect 29092 10548 29144 10600
rect 31024 10548 31076 10600
rect 31208 10591 31260 10600
rect 31208 10557 31217 10591
rect 31217 10557 31251 10591
rect 31251 10557 31260 10591
rect 31208 10548 31260 10557
rect 32588 10659 32640 10668
rect 32588 10625 32597 10659
rect 32597 10625 32631 10659
rect 32631 10625 32640 10659
rect 32588 10616 32640 10625
rect 32772 10659 32824 10668
rect 32772 10625 32781 10659
rect 32781 10625 32815 10659
rect 32815 10625 32824 10659
rect 32772 10616 32824 10625
rect 34888 10684 34940 10736
rect 35072 10727 35124 10736
rect 35072 10693 35081 10727
rect 35081 10693 35115 10727
rect 35115 10693 35124 10727
rect 35072 10684 35124 10693
rect 33048 10659 33100 10668
rect 33048 10625 33057 10659
rect 33057 10625 33091 10659
rect 33091 10625 33100 10659
rect 33048 10616 33100 10625
rect 34428 10659 34480 10668
rect 34428 10625 34437 10659
rect 34437 10625 34471 10659
rect 34471 10625 34480 10659
rect 34428 10616 34480 10625
rect 35348 10616 35400 10668
rect 36084 10684 36136 10736
rect 35624 10659 35676 10668
rect 35624 10625 35633 10659
rect 35633 10625 35667 10659
rect 35667 10625 35676 10659
rect 35624 10616 35676 10625
rect 35900 10659 35952 10668
rect 35900 10625 35909 10659
rect 35909 10625 35943 10659
rect 35943 10625 35952 10659
rect 35900 10616 35952 10625
rect 36452 10659 36504 10668
rect 36452 10625 36461 10659
rect 36461 10625 36495 10659
rect 36495 10625 36504 10659
rect 36452 10616 36504 10625
rect 36636 10616 36688 10668
rect 37188 10684 37240 10736
rect 39580 10752 39632 10804
rect 38200 10727 38252 10736
rect 38200 10693 38209 10727
rect 38209 10693 38243 10727
rect 38243 10693 38252 10727
rect 38200 10684 38252 10693
rect 38384 10684 38436 10736
rect 38476 10616 38528 10668
rect 22008 10523 22060 10532
rect 22008 10489 22017 10523
rect 22017 10489 22051 10523
rect 22051 10489 22060 10523
rect 22008 10480 22060 10489
rect 21640 10455 21692 10464
rect 21640 10421 21649 10455
rect 21649 10421 21683 10455
rect 21683 10421 21692 10455
rect 21640 10412 21692 10421
rect 28724 10480 28776 10532
rect 27252 10412 27304 10464
rect 31760 10480 31812 10532
rect 34704 10523 34756 10532
rect 34704 10489 34713 10523
rect 34713 10489 34747 10523
rect 34747 10489 34756 10523
rect 34704 10480 34756 10489
rect 35624 10480 35676 10532
rect 38292 10548 38344 10600
rect 39304 10659 39356 10668
rect 39304 10625 39313 10659
rect 39313 10625 39347 10659
rect 39347 10625 39356 10659
rect 39304 10616 39356 10625
rect 40592 10616 40644 10668
rect 29460 10455 29512 10464
rect 29460 10421 29469 10455
rect 29469 10421 29503 10455
rect 29503 10421 29512 10455
rect 29460 10412 29512 10421
rect 30472 10412 30524 10464
rect 32312 10412 32364 10464
rect 34612 10412 34664 10464
rect 35808 10455 35860 10464
rect 35808 10421 35817 10455
rect 35817 10421 35851 10455
rect 35851 10421 35860 10455
rect 35808 10412 35860 10421
rect 35900 10412 35952 10464
rect 36084 10412 36136 10464
rect 37464 10412 37516 10464
rect 37556 10455 37608 10464
rect 37556 10421 37565 10455
rect 37565 10421 37599 10455
rect 37599 10421 37608 10455
rect 37556 10412 37608 10421
rect 37832 10455 37884 10464
rect 37832 10421 37841 10455
rect 37841 10421 37875 10455
rect 37875 10421 37884 10455
rect 37832 10412 37884 10421
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 13544 10140 13596 10192
rect 13912 10183 13964 10192
rect 13912 10149 13921 10183
rect 13921 10149 13955 10183
rect 13955 10149 13964 10183
rect 13912 10140 13964 10149
rect 14096 10047 14148 10056
rect 14096 10013 14105 10047
rect 14105 10013 14139 10047
rect 14139 10013 14148 10047
rect 14096 10004 14148 10013
rect 17316 10208 17368 10260
rect 17960 10208 18012 10260
rect 22008 10208 22060 10260
rect 22560 10251 22612 10260
rect 22560 10217 22569 10251
rect 22569 10217 22603 10251
rect 22603 10217 22612 10251
rect 22560 10208 22612 10217
rect 22836 10251 22888 10260
rect 22836 10217 22845 10251
rect 22845 10217 22879 10251
rect 22879 10217 22888 10251
rect 22836 10208 22888 10217
rect 25872 10251 25924 10260
rect 25872 10217 25881 10251
rect 25881 10217 25915 10251
rect 25915 10217 25924 10251
rect 25872 10208 25924 10217
rect 27712 10251 27764 10260
rect 27712 10217 27721 10251
rect 27721 10217 27755 10251
rect 27755 10217 27764 10251
rect 27712 10208 27764 10217
rect 29368 10208 29420 10260
rect 29460 10208 29512 10260
rect 18052 10140 18104 10192
rect 21640 10140 21692 10192
rect 18328 10072 18380 10124
rect 23112 10072 23164 10124
rect 16120 10047 16172 10056
rect 16120 10013 16129 10047
rect 16129 10013 16163 10047
rect 16163 10013 16172 10047
rect 16120 10004 16172 10013
rect 19984 10004 20036 10056
rect 20076 10004 20128 10056
rect 20260 10047 20312 10056
rect 20260 10013 20269 10047
rect 20269 10013 20303 10047
rect 20303 10013 20312 10047
rect 20260 10004 20312 10013
rect 22560 10004 22612 10056
rect 23020 10047 23072 10056
rect 23020 10013 23029 10047
rect 23029 10013 23063 10047
rect 23063 10013 23072 10047
rect 23020 10004 23072 10013
rect 27620 10140 27672 10192
rect 30472 10208 30524 10260
rect 30932 10208 30984 10260
rect 31208 10208 31260 10260
rect 32220 10208 32272 10260
rect 32956 10208 33008 10260
rect 30380 10115 30432 10124
rect 30380 10081 30389 10115
rect 30389 10081 30423 10115
rect 30423 10081 30432 10115
rect 30380 10072 30432 10081
rect 30472 10072 30524 10124
rect 12348 9936 12400 9988
rect 13728 9936 13780 9988
rect 13912 9936 13964 9988
rect 16856 9979 16908 9988
rect 16856 9945 16865 9979
rect 16865 9945 16899 9979
rect 16899 9945 16908 9979
rect 16856 9936 16908 9945
rect 14832 9868 14884 9920
rect 16764 9868 16816 9920
rect 17684 9868 17736 9920
rect 22100 9936 22152 9988
rect 21364 9868 21416 9920
rect 22376 9911 22428 9920
rect 22376 9877 22401 9911
rect 22401 9877 22428 9911
rect 22376 9868 22428 9877
rect 23664 9868 23716 9920
rect 27344 10047 27396 10056
rect 27344 10013 27353 10047
rect 27353 10013 27387 10047
rect 27387 10013 27396 10047
rect 27344 10004 27396 10013
rect 27712 10004 27764 10056
rect 28724 9936 28776 9988
rect 29000 9936 29052 9988
rect 29092 9979 29144 9988
rect 29092 9945 29101 9979
rect 29101 9945 29135 9979
rect 29135 9945 29144 9979
rect 29092 9936 29144 9945
rect 31300 10140 31352 10192
rect 32128 10140 32180 10192
rect 31208 10004 31260 10056
rect 31484 10072 31536 10124
rect 32312 10072 32364 10124
rect 32680 10115 32732 10124
rect 32680 10081 32689 10115
rect 32689 10081 32723 10115
rect 32723 10081 32732 10115
rect 32680 10072 32732 10081
rect 31944 10004 31996 10056
rect 32036 9868 32088 9920
rect 32312 9936 32364 9988
rect 32588 10047 32640 10056
rect 32588 10013 32597 10047
rect 32597 10013 32631 10047
rect 32631 10013 32640 10047
rect 35348 10208 35400 10260
rect 35808 10208 35860 10260
rect 38108 10208 38160 10260
rect 38568 10208 38620 10260
rect 34796 10140 34848 10192
rect 36176 10183 36228 10192
rect 36176 10149 36185 10183
rect 36185 10149 36219 10183
rect 36219 10149 36228 10183
rect 36176 10140 36228 10149
rect 36268 10140 36320 10192
rect 35900 10115 35952 10124
rect 35900 10081 35909 10115
rect 35909 10081 35943 10115
rect 35943 10081 35952 10115
rect 35900 10072 35952 10081
rect 32588 10004 32640 10013
rect 33784 10004 33836 10056
rect 33692 9936 33744 9988
rect 36176 9936 36228 9988
rect 36360 10047 36412 10056
rect 36360 10013 36372 10047
rect 36372 10013 36406 10047
rect 36406 10013 36412 10047
rect 36360 10004 36412 10013
rect 36452 9936 36504 9988
rect 37004 10004 37056 10056
rect 37188 10047 37240 10056
rect 37188 10013 37197 10047
rect 37197 10013 37231 10047
rect 37231 10013 37240 10047
rect 37188 10004 37240 10013
rect 39212 10115 39264 10124
rect 39212 10081 39221 10115
rect 39221 10081 39255 10115
rect 39255 10081 39264 10115
rect 39212 10072 39264 10081
rect 40132 10072 40184 10124
rect 40592 10072 40644 10124
rect 41236 10072 41288 10124
rect 32772 9868 32824 9920
rect 35808 9868 35860 9920
rect 36084 9868 36136 9920
rect 37280 9936 37332 9988
rect 37556 9936 37608 9988
rect 40040 10004 40092 10056
rect 37096 9868 37148 9920
rect 41512 9936 41564 9988
rect 4874 9766 4926 9818
rect 4938 9766 4990 9818
rect 5002 9766 5054 9818
rect 5066 9766 5118 9818
rect 5130 9766 5182 9818
rect 35594 9766 35646 9818
rect 35658 9766 35710 9818
rect 35722 9766 35774 9818
rect 35786 9766 35838 9818
rect 35850 9766 35902 9818
rect 14832 9707 14884 9716
rect 14832 9673 14841 9707
rect 14841 9673 14875 9707
rect 14875 9673 14884 9707
rect 14832 9664 14884 9673
rect 16856 9707 16908 9716
rect 16856 9673 16865 9707
rect 16865 9673 16899 9707
rect 16899 9673 16908 9707
rect 16856 9664 16908 9673
rect 23296 9664 23348 9716
rect 27712 9664 27764 9716
rect 29276 9707 29328 9716
rect 29276 9673 29285 9707
rect 29285 9673 29319 9707
rect 29319 9673 29328 9707
rect 29276 9664 29328 9673
rect 30380 9664 30432 9716
rect 13452 9596 13504 9648
rect 12348 9460 12400 9512
rect 12440 9460 12492 9512
rect 13728 9460 13780 9512
rect 15476 9596 15528 9648
rect 16764 9571 16816 9580
rect 16764 9537 16773 9571
rect 16773 9537 16807 9571
rect 16807 9537 16816 9571
rect 16764 9528 16816 9537
rect 16948 9571 17000 9580
rect 16948 9537 16957 9571
rect 16957 9537 16991 9571
rect 16991 9537 17000 9571
rect 16948 9528 17000 9537
rect 21824 9571 21876 9580
rect 21824 9537 21833 9571
rect 21833 9537 21867 9571
rect 21867 9537 21876 9571
rect 21824 9528 21876 9537
rect 21916 9571 21968 9580
rect 21916 9537 21925 9571
rect 21925 9537 21959 9571
rect 21959 9537 21968 9571
rect 21916 9528 21968 9537
rect 29000 9596 29052 9648
rect 32588 9664 32640 9716
rect 32956 9664 33008 9716
rect 28724 9571 28776 9580
rect 28724 9537 28733 9571
rect 28733 9537 28767 9571
rect 28767 9537 28776 9571
rect 28724 9528 28776 9537
rect 29092 9571 29144 9580
rect 29092 9537 29101 9571
rect 29101 9537 29135 9571
rect 29135 9537 29144 9571
rect 29092 9528 29144 9537
rect 32036 9596 32088 9648
rect 21732 9460 21784 9512
rect 23480 9503 23532 9512
rect 23480 9469 23489 9503
rect 23489 9469 23523 9503
rect 23523 9469 23532 9503
rect 23480 9460 23532 9469
rect 28816 9460 28868 9512
rect 23020 9392 23072 9444
rect 32128 9528 32180 9580
rect 31484 9460 31536 9512
rect 32588 9571 32640 9580
rect 32588 9537 32597 9571
rect 32597 9537 32631 9571
rect 32631 9537 32640 9571
rect 32588 9528 32640 9537
rect 32956 9571 33008 9580
rect 32956 9537 32965 9571
rect 32965 9537 32999 9571
rect 32999 9537 33008 9571
rect 32956 9528 33008 9537
rect 36912 9596 36964 9648
rect 40132 9664 40184 9716
rect 39212 9596 39264 9648
rect 33232 9571 33284 9580
rect 33232 9537 33241 9571
rect 33241 9537 33275 9571
rect 33275 9537 33284 9571
rect 33232 9528 33284 9537
rect 33784 9571 33836 9580
rect 33784 9537 33793 9571
rect 33793 9537 33827 9571
rect 33827 9537 33836 9571
rect 33784 9528 33836 9537
rect 33416 9460 33468 9512
rect 36636 9528 36688 9580
rect 37096 9571 37148 9580
rect 37096 9537 37105 9571
rect 37105 9537 37139 9571
rect 37139 9537 37148 9571
rect 37096 9528 37148 9537
rect 37280 9528 37332 9580
rect 41236 9571 41288 9580
rect 41236 9537 41245 9571
rect 41245 9537 41279 9571
rect 41279 9537 41288 9571
rect 41236 9528 41288 9537
rect 31852 9392 31904 9444
rect 31944 9392 31996 9444
rect 32588 9392 32640 9444
rect 22468 9324 22520 9376
rect 27988 9324 28040 9376
rect 28816 9324 28868 9376
rect 31208 9324 31260 9376
rect 32312 9367 32364 9376
rect 32312 9333 32321 9367
rect 32321 9333 32355 9367
rect 32355 9333 32364 9367
rect 32312 9324 32364 9333
rect 32404 9324 32456 9376
rect 33416 9367 33468 9376
rect 33416 9333 33425 9367
rect 33425 9333 33459 9367
rect 33459 9333 33468 9367
rect 33416 9324 33468 9333
rect 34704 9392 34756 9444
rect 36820 9324 36872 9376
rect 39396 9324 39448 9376
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 21180 9120 21232 9172
rect 21916 9163 21968 9172
rect 16672 8916 16724 8968
rect 21916 9129 21925 9163
rect 21925 9129 21959 9163
rect 21959 9129 21968 9163
rect 21916 9120 21968 9129
rect 21732 9052 21784 9104
rect 28080 9120 28132 9172
rect 28816 9163 28868 9172
rect 28816 9129 28825 9163
rect 28825 9129 28859 9163
rect 28859 9129 28868 9163
rect 28816 9120 28868 9129
rect 29092 9120 29144 9172
rect 31944 9120 31996 9172
rect 32220 9163 32272 9172
rect 32220 9129 32229 9163
rect 32229 9129 32263 9163
rect 32263 9129 32272 9163
rect 32220 9120 32272 9129
rect 33232 9120 33284 9172
rect 36636 9120 36688 9172
rect 36728 9120 36780 9172
rect 38016 9120 38068 9172
rect 22376 9052 22428 9104
rect 27804 9052 27856 9104
rect 32128 9052 32180 9104
rect 33048 9052 33100 9104
rect 23664 9027 23716 9036
rect 23664 8993 23673 9027
rect 23673 8993 23707 9027
rect 23707 8993 23716 9027
rect 23664 8984 23716 8993
rect 28540 9027 28592 9036
rect 28540 8993 28549 9027
rect 28549 8993 28583 9027
rect 28583 8993 28592 9027
rect 28540 8984 28592 8993
rect 19984 8848 20036 8900
rect 23940 8959 23992 8968
rect 23940 8925 23949 8959
rect 23949 8925 23983 8959
rect 23983 8925 23992 8959
rect 23940 8916 23992 8925
rect 21548 8891 21600 8900
rect 21548 8857 21557 8891
rect 21557 8857 21591 8891
rect 21591 8857 21600 8891
rect 21548 8848 21600 8857
rect 21732 8891 21784 8900
rect 21732 8857 21741 8891
rect 21741 8857 21775 8891
rect 21775 8857 21784 8891
rect 21732 8848 21784 8857
rect 21824 8848 21876 8900
rect 27620 8959 27672 8968
rect 27620 8925 27629 8959
rect 27629 8925 27663 8959
rect 27663 8925 27672 8959
rect 27620 8916 27672 8925
rect 28632 8916 28684 8968
rect 31760 8916 31812 8968
rect 32312 8959 32364 8968
rect 32312 8925 32321 8959
rect 32321 8925 32355 8959
rect 32355 8925 32364 8959
rect 32312 8916 32364 8925
rect 32496 8916 32548 8968
rect 36728 8984 36780 9036
rect 36820 9027 36872 9036
rect 36820 8993 36829 9027
rect 36829 8993 36863 9027
rect 36863 8993 36872 9027
rect 36820 8984 36872 8993
rect 40040 8984 40092 9036
rect 37096 8959 37148 8968
rect 37096 8925 37105 8959
rect 37105 8925 37139 8959
rect 37139 8925 37148 8959
rect 37096 8916 37148 8925
rect 27804 8848 27856 8900
rect 36544 8848 36596 8900
rect 18144 8780 18196 8832
rect 20720 8823 20772 8832
rect 20720 8789 20729 8823
rect 20729 8789 20763 8823
rect 20763 8789 20772 8823
rect 20720 8780 20772 8789
rect 21088 8780 21140 8832
rect 21364 8823 21416 8832
rect 21364 8789 21373 8823
rect 21373 8789 21407 8823
rect 21407 8789 21416 8823
rect 21364 8780 21416 8789
rect 27344 8780 27396 8832
rect 32956 8780 33008 8832
rect 35992 8780 36044 8832
rect 36728 8780 36780 8832
rect 38016 8848 38068 8900
rect 39396 8891 39448 8900
rect 39396 8857 39405 8891
rect 39405 8857 39439 8891
rect 39439 8857 39448 8891
rect 39396 8848 39448 8857
rect 4874 8678 4926 8730
rect 4938 8678 4990 8730
rect 5002 8678 5054 8730
rect 5066 8678 5118 8730
rect 5130 8678 5182 8730
rect 35594 8678 35646 8730
rect 35658 8678 35710 8730
rect 35722 8678 35774 8730
rect 35786 8678 35838 8730
rect 35850 8678 35902 8730
rect 15292 8440 15344 8492
rect 18328 8576 18380 8628
rect 21180 8619 21232 8628
rect 21180 8585 21189 8619
rect 21189 8585 21223 8619
rect 21223 8585 21232 8619
rect 21180 8576 21232 8585
rect 17684 8508 17736 8560
rect 15844 8483 15896 8492
rect 15844 8449 15853 8483
rect 15853 8449 15887 8483
rect 15887 8449 15896 8483
rect 15844 8440 15896 8449
rect 16028 8483 16080 8492
rect 16028 8449 16037 8483
rect 16037 8449 16071 8483
rect 16071 8449 16080 8483
rect 16028 8440 16080 8449
rect 18420 8483 18472 8492
rect 18420 8449 18429 8483
rect 18429 8449 18463 8483
rect 18463 8449 18472 8483
rect 18420 8440 18472 8449
rect 20720 8440 20772 8492
rect 21732 8508 21784 8560
rect 15936 8372 15988 8424
rect 16672 8415 16724 8424
rect 16672 8381 16681 8415
rect 16681 8381 16715 8415
rect 16715 8381 16724 8415
rect 16672 8372 16724 8381
rect 18052 8372 18104 8424
rect 19432 8415 19484 8424
rect 19432 8381 19441 8415
rect 19441 8381 19475 8415
rect 19475 8381 19484 8415
rect 19432 8372 19484 8381
rect 21548 8440 21600 8492
rect 23480 8576 23532 8628
rect 29000 8619 29052 8628
rect 29000 8585 29009 8619
rect 29009 8585 29043 8619
rect 29043 8585 29052 8619
rect 29000 8576 29052 8585
rect 31484 8619 31536 8628
rect 31484 8585 31493 8619
rect 31493 8585 31527 8619
rect 31527 8585 31536 8619
rect 31484 8576 31536 8585
rect 32588 8576 32640 8628
rect 37280 8576 37332 8628
rect 37832 8576 37884 8628
rect 22928 8508 22980 8560
rect 26608 8508 26660 8560
rect 32312 8508 32364 8560
rect 22468 8483 22520 8492
rect 22468 8449 22477 8483
rect 22477 8449 22511 8483
rect 22511 8449 22520 8483
rect 22468 8440 22520 8449
rect 31300 8483 31352 8492
rect 31300 8449 31309 8483
rect 31309 8449 31343 8483
rect 31343 8449 31352 8483
rect 31300 8440 31352 8449
rect 21824 8372 21876 8424
rect 22928 8304 22980 8356
rect 16120 8236 16172 8288
rect 21364 8279 21416 8288
rect 21364 8245 21373 8279
rect 21373 8245 21407 8279
rect 21407 8245 21416 8279
rect 21364 8236 21416 8245
rect 23940 8236 23992 8288
rect 25320 8415 25372 8424
rect 25320 8381 25329 8415
rect 25329 8381 25363 8415
rect 25363 8381 25372 8415
rect 25320 8372 25372 8381
rect 27068 8372 27120 8424
rect 27620 8372 27672 8424
rect 28540 8372 28592 8424
rect 32496 8440 32548 8492
rect 28080 8304 28132 8356
rect 32220 8372 32272 8424
rect 36084 8551 36136 8560
rect 36084 8517 36093 8551
rect 36093 8517 36127 8551
rect 36127 8517 36136 8551
rect 36084 8508 36136 8517
rect 35808 8483 35860 8492
rect 35808 8449 35817 8483
rect 35817 8449 35851 8483
rect 35851 8449 35860 8483
rect 35808 8440 35860 8449
rect 35992 8483 36044 8492
rect 35992 8449 36001 8483
rect 36001 8449 36035 8483
rect 36035 8449 36044 8483
rect 35992 8440 36044 8449
rect 26976 8279 27028 8288
rect 26976 8245 26985 8279
rect 26985 8245 27019 8279
rect 27019 8245 27028 8279
rect 26976 8236 27028 8245
rect 28448 8236 28500 8288
rect 28632 8279 28684 8288
rect 28632 8245 28641 8279
rect 28641 8245 28675 8279
rect 28675 8245 28684 8279
rect 28632 8236 28684 8245
rect 31760 8279 31812 8288
rect 31760 8245 31769 8279
rect 31769 8245 31803 8279
rect 31803 8245 31812 8279
rect 31760 8236 31812 8245
rect 32496 8279 32548 8288
rect 32496 8245 32505 8279
rect 32505 8245 32539 8279
rect 32539 8245 32548 8279
rect 32496 8236 32548 8245
rect 36636 8483 36688 8492
rect 36636 8449 36645 8483
rect 36645 8449 36679 8483
rect 36679 8449 36688 8483
rect 36636 8440 36688 8449
rect 36728 8483 36780 8492
rect 36728 8449 36737 8483
rect 36737 8449 36771 8483
rect 36771 8449 36780 8483
rect 36728 8440 36780 8449
rect 37372 8483 37424 8492
rect 37372 8449 37381 8483
rect 37381 8449 37415 8483
rect 37415 8449 37424 8483
rect 37372 8440 37424 8449
rect 38016 8508 38068 8560
rect 41512 8576 41564 8628
rect 40040 8508 40092 8560
rect 36912 8372 36964 8424
rect 40316 8415 40368 8424
rect 40316 8381 40325 8415
rect 40325 8381 40359 8415
rect 40359 8381 40368 8415
rect 40316 8372 40368 8381
rect 36360 8304 36412 8356
rect 32680 8236 32732 8288
rect 36268 8236 36320 8288
rect 37556 8236 37608 8288
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 16028 8032 16080 8084
rect 12072 7896 12124 7948
rect 12440 7896 12492 7948
rect 15384 7896 15436 7948
rect 19432 8032 19484 8084
rect 21732 8075 21784 8084
rect 21732 8041 21741 8075
rect 21741 8041 21775 8075
rect 21775 8041 21784 8075
rect 21732 8032 21784 8041
rect 21824 8032 21876 8084
rect 25320 8032 25372 8084
rect 28632 8032 28684 8084
rect 29092 8032 29144 8084
rect 32128 8075 32180 8084
rect 32128 8041 32137 8075
rect 32137 8041 32171 8075
rect 32171 8041 32180 8075
rect 32128 8032 32180 8041
rect 37832 8075 37884 8084
rect 37832 8041 37841 8075
rect 37841 8041 37875 8075
rect 37875 8041 37884 8075
rect 37832 8032 37884 8041
rect 40316 8032 40368 8084
rect 16212 7964 16264 8016
rect 16488 7896 16540 7948
rect 15476 7828 15528 7880
rect 17684 7896 17736 7948
rect 16672 7871 16724 7880
rect 16672 7837 16681 7871
rect 16681 7837 16715 7871
rect 16715 7837 16724 7871
rect 16672 7828 16724 7837
rect 16856 7871 16908 7880
rect 16856 7837 16865 7871
rect 16865 7837 16899 7871
rect 16899 7837 16908 7871
rect 16856 7828 16908 7837
rect 17224 7871 17276 7880
rect 17224 7837 17233 7871
rect 17233 7837 17267 7871
rect 17267 7837 17276 7871
rect 17224 7828 17276 7837
rect 27804 7964 27856 8016
rect 28448 8007 28500 8016
rect 28448 7973 28457 8007
rect 28457 7973 28491 8007
rect 28491 7973 28500 8007
rect 28448 7964 28500 7973
rect 31760 7964 31812 8016
rect 32496 7964 32548 8016
rect 33784 7964 33836 8016
rect 36268 7964 36320 8016
rect 21088 7896 21140 7948
rect 21548 7896 21600 7948
rect 26792 7896 26844 7948
rect 12440 7803 12492 7812
rect 12440 7769 12449 7803
rect 12449 7769 12483 7803
rect 12483 7769 12492 7803
rect 12440 7760 12492 7769
rect 13728 7760 13780 7812
rect 14372 7803 14424 7812
rect 14372 7769 14381 7803
rect 14381 7769 14415 7803
rect 14415 7769 14424 7803
rect 14372 7760 14424 7769
rect 18144 7871 18196 7880
rect 18144 7837 18153 7871
rect 18153 7837 18187 7871
rect 18187 7837 18196 7871
rect 18144 7828 18196 7837
rect 14004 7692 14056 7744
rect 15844 7692 15896 7744
rect 21180 7760 21232 7812
rect 26976 7828 27028 7880
rect 27068 7871 27120 7880
rect 27068 7837 27077 7871
rect 27077 7837 27111 7871
rect 27111 7837 27120 7871
rect 27068 7828 27120 7837
rect 27344 7896 27396 7948
rect 28540 7896 28592 7948
rect 30840 7896 30892 7948
rect 31300 7896 31352 7948
rect 28080 7871 28132 7880
rect 28080 7837 28089 7871
rect 28089 7837 28123 7871
rect 28123 7837 28132 7871
rect 28080 7828 28132 7837
rect 28724 7828 28776 7880
rect 29552 7871 29604 7880
rect 29552 7837 29561 7871
rect 29561 7837 29595 7871
rect 29595 7837 29604 7871
rect 29552 7828 29604 7837
rect 32680 7828 32732 7880
rect 34428 7896 34480 7948
rect 34520 7896 34572 7948
rect 35808 7896 35860 7948
rect 33876 7828 33928 7880
rect 36360 7871 36412 7880
rect 36360 7837 36369 7871
rect 36369 7837 36403 7871
rect 36403 7837 36412 7871
rect 36360 7828 36412 7837
rect 36636 7939 36688 7948
rect 36636 7905 36645 7939
rect 36645 7905 36679 7939
rect 36679 7905 36688 7939
rect 36636 7896 36688 7905
rect 37004 7939 37056 7948
rect 37004 7905 37013 7939
rect 37013 7905 37047 7939
rect 37047 7905 37056 7939
rect 37004 7896 37056 7905
rect 37556 7828 37608 7880
rect 37648 7871 37700 7880
rect 37648 7837 37657 7871
rect 37657 7837 37691 7871
rect 37691 7837 37700 7871
rect 37648 7828 37700 7837
rect 38016 7871 38068 7880
rect 38016 7837 38025 7871
rect 38025 7837 38059 7871
rect 38059 7837 38068 7871
rect 38016 7828 38068 7837
rect 40040 7871 40092 7880
rect 40040 7837 40049 7871
rect 40049 7837 40083 7871
rect 40083 7837 40092 7871
rect 40040 7828 40092 7837
rect 41052 8032 41104 8084
rect 16028 7692 16080 7744
rect 16948 7692 17000 7744
rect 17592 7692 17644 7744
rect 21364 7692 21416 7744
rect 26148 7692 26200 7744
rect 29828 7803 29880 7812
rect 29828 7769 29837 7803
rect 29837 7769 29871 7803
rect 29871 7769 29880 7803
rect 29828 7760 29880 7769
rect 30380 7760 30432 7812
rect 31300 7735 31352 7744
rect 31300 7701 31309 7735
rect 31309 7701 31343 7735
rect 31343 7701 31352 7735
rect 31300 7692 31352 7701
rect 37188 7692 37240 7744
rect 38752 7692 38804 7744
rect 4874 7590 4926 7642
rect 4938 7590 4990 7642
rect 5002 7590 5054 7642
rect 5066 7590 5118 7642
rect 5130 7590 5182 7642
rect 35594 7590 35646 7642
rect 35658 7590 35710 7642
rect 35722 7590 35774 7642
rect 35786 7590 35838 7642
rect 35850 7590 35902 7642
rect 14372 7488 14424 7540
rect 16672 7488 16724 7540
rect 18052 7488 18104 7540
rect 21088 7488 21140 7540
rect 23296 7531 23348 7540
rect 15292 7463 15344 7472
rect 15292 7429 15301 7463
rect 15301 7429 15335 7463
rect 15335 7429 15344 7463
rect 15292 7420 15344 7429
rect 16580 7420 16632 7472
rect 23296 7497 23305 7531
rect 23305 7497 23339 7531
rect 23339 7497 23348 7531
rect 23296 7488 23348 7497
rect 27252 7488 27304 7540
rect 14004 7395 14056 7404
rect 14004 7361 14013 7395
rect 14013 7361 14047 7395
rect 14047 7361 14056 7395
rect 14004 7352 14056 7361
rect 16120 7395 16172 7404
rect 16120 7361 16129 7395
rect 16129 7361 16163 7395
rect 16163 7361 16172 7395
rect 16120 7352 16172 7361
rect 16212 7395 16264 7404
rect 16212 7361 16221 7395
rect 16221 7361 16255 7395
rect 16255 7361 16264 7395
rect 16212 7352 16264 7361
rect 16488 7352 16540 7404
rect 12440 7327 12492 7336
rect 12440 7293 12449 7327
rect 12449 7293 12483 7327
rect 12483 7293 12492 7327
rect 12440 7284 12492 7293
rect 12900 7327 12952 7336
rect 12900 7293 12909 7327
rect 12909 7293 12943 7327
rect 12943 7293 12952 7327
rect 12900 7284 12952 7293
rect 16948 7284 17000 7336
rect 15844 7216 15896 7268
rect 17408 7395 17460 7404
rect 17408 7361 17417 7395
rect 17417 7361 17451 7395
rect 17451 7361 17460 7395
rect 17408 7352 17460 7361
rect 17592 7395 17644 7404
rect 17592 7361 17601 7395
rect 17601 7361 17635 7395
rect 17635 7361 17644 7395
rect 17592 7352 17644 7361
rect 20352 7395 20404 7404
rect 20352 7361 20361 7395
rect 20361 7361 20395 7395
rect 20395 7361 20404 7395
rect 20352 7352 20404 7361
rect 20444 7395 20496 7404
rect 20444 7361 20453 7395
rect 20453 7361 20487 7395
rect 20487 7361 20496 7395
rect 20444 7352 20496 7361
rect 20536 7395 20588 7404
rect 20536 7361 20545 7395
rect 20545 7361 20579 7395
rect 20579 7361 20588 7395
rect 20536 7352 20588 7361
rect 20260 7284 20312 7336
rect 17132 7216 17184 7268
rect 20720 7259 20772 7268
rect 20720 7225 20729 7259
rect 20729 7225 20763 7259
rect 20763 7225 20772 7259
rect 20720 7216 20772 7225
rect 21364 7395 21416 7404
rect 21364 7361 21373 7395
rect 21373 7361 21407 7395
rect 21407 7361 21416 7395
rect 21364 7352 21416 7361
rect 23020 7395 23072 7404
rect 23020 7361 23029 7395
rect 23029 7361 23063 7395
rect 23063 7361 23072 7395
rect 23020 7352 23072 7361
rect 23112 7352 23164 7404
rect 27620 7395 27672 7404
rect 27620 7361 27629 7395
rect 27629 7361 27663 7395
rect 27663 7361 27672 7395
rect 27620 7352 27672 7361
rect 22008 7284 22060 7336
rect 23940 7284 23992 7336
rect 26240 7284 26292 7336
rect 23112 7216 23164 7268
rect 26608 7284 26660 7336
rect 28540 7352 28592 7404
rect 30380 7488 30432 7540
rect 31852 7531 31904 7540
rect 31852 7497 31861 7531
rect 31861 7497 31895 7531
rect 31895 7497 31904 7531
rect 31852 7488 31904 7497
rect 33876 7531 33928 7540
rect 33876 7497 33885 7531
rect 33885 7497 33919 7531
rect 33919 7497 33928 7531
rect 33876 7488 33928 7497
rect 29552 7420 29604 7472
rect 31300 7395 31352 7404
rect 31300 7361 31309 7395
rect 31309 7361 31343 7395
rect 31343 7361 31352 7395
rect 31300 7352 31352 7361
rect 32864 7420 32916 7472
rect 34796 7420 34848 7472
rect 36636 7488 36688 7540
rect 38016 7488 38068 7540
rect 37188 7420 37240 7472
rect 37924 7420 37976 7472
rect 26792 7216 26844 7268
rect 16764 7148 16816 7200
rect 21272 7148 21324 7200
rect 23848 7148 23900 7200
rect 25964 7191 26016 7200
rect 25964 7157 25973 7191
rect 25973 7157 26007 7191
rect 26007 7157 26016 7191
rect 25964 7148 26016 7157
rect 28172 7148 28224 7200
rect 29828 7216 29880 7268
rect 30656 7216 30708 7268
rect 29276 7148 29328 7200
rect 32404 7327 32456 7336
rect 32404 7293 32413 7327
rect 32413 7293 32447 7327
rect 32447 7293 32456 7327
rect 32404 7284 32456 7293
rect 35440 7284 35492 7336
rect 36360 7284 36412 7336
rect 36544 7395 36596 7404
rect 36544 7361 36553 7395
rect 36553 7361 36587 7395
rect 36587 7361 36596 7395
rect 36544 7352 36596 7361
rect 36728 7395 36780 7404
rect 36728 7361 36737 7395
rect 36737 7361 36771 7395
rect 36771 7361 36780 7395
rect 36728 7352 36780 7361
rect 37004 7352 37056 7404
rect 38752 7395 38804 7404
rect 38752 7361 38761 7395
rect 38761 7361 38795 7395
rect 38795 7361 38804 7395
rect 38752 7352 38804 7361
rect 40040 7352 40092 7404
rect 37648 7284 37700 7336
rect 37004 7216 37056 7268
rect 31668 7148 31720 7200
rect 32956 7148 33008 7200
rect 33140 7148 33192 7200
rect 35348 7191 35400 7200
rect 35348 7157 35357 7191
rect 35357 7157 35391 7191
rect 35391 7157 35400 7191
rect 35348 7148 35400 7157
rect 36176 7148 36228 7200
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 23848 6944 23900 6996
rect 25964 6944 26016 6996
rect 26240 6944 26292 6996
rect 15844 6876 15896 6928
rect 14740 6783 14792 6792
rect 14740 6749 14749 6783
rect 14749 6749 14783 6783
rect 14783 6749 14792 6783
rect 14740 6740 14792 6749
rect 16488 6808 16540 6860
rect 16580 6851 16632 6860
rect 16580 6817 16589 6851
rect 16589 6817 16623 6851
rect 16623 6817 16632 6851
rect 16580 6808 16632 6817
rect 16764 6740 16816 6792
rect 17684 6740 17736 6792
rect 20720 6808 20772 6860
rect 21364 6808 21416 6860
rect 20260 6740 20312 6792
rect 20536 6783 20588 6792
rect 20536 6749 20545 6783
rect 20545 6749 20579 6783
rect 20579 6749 20588 6783
rect 20536 6740 20588 6749
rect 20812 6740 20864 6792
rect 21732 6740 21784 6792
rect 22008 6783 22060 6792
rect 22008 6749 22017 6783
rect 22017 6749 22051 6783
rect 22051 6749 22060 6783
rect 22008 6740 22060 6749
rect 17408 6672 17460 6724
rect 20352 6672 20404 6724
rect 14096 6647 14148 6656
rect 14096 6613 14105 6647
rect 14105 6613 14139 6647
rect 14139 6613 14148 6647
rect 14096 6604 14148 6613
rect 14924 6604 14976 6656
rect 16028 6604 16080 6656
rect 18144 6647 18196 6656
rect 18144 6613 18153 6647
rect 18153 6613 18187 6647
rect 18187 6613 18196 6647
rect 18144 6604 18196 6613
rect 20628 6647 20680 6656
rect 20628 6613 20637 6647
rect 20637 6613 20671 6647
rect 20671 6613 20680 6647
rect 20628 6604 20680 6613
rect 21916 6672 21968 6724
rect 22928 6808 22980 6860
rect 23572 6808 23624 6860
rect 27252 6740 27304 6792
rect 27344 6783 27396 6792
rect 27344 6749 27353 6783
rect 27353 6749 27387 6783
rect 27387 6749 27396 6783
rect 27344 6740 27396 6749
rect 27436 6783 27488 6792
rect 27436 6749 27445 6783
rect 27445 6749 27479 6783
rect 27479 6749 27488 6783
rect 27436 6740 27488 6749
rect 22928 6672 22980 6724
rect 26056 6672 26108 6724
rect 28540 6944 28592 6996
rect 32404 6944 32456 6996
rect 32864 6944 32916 6996
rect 34612 6944 34664 6996
rect 36544 6987 36596 6996
rect 36544 6953 36553 6987
rect 36553 6953 36587 6987
rect 36587 6953 36596 6987
rect 36544 6944 36596 6953
rect 36728 6944 36780 6996
rect 33048 6876 33100 6928
rect 34520 6876 34572 6928
rect 30656 6851 30708 6860
rect 30656 6817 30665 6851
rect 30665 6817 30699 6851
rect 30699 6817 30708 6851
rect 30656 6808 30708 6817
rect 32864 6851 32916 6860
rect 32864 6817 32873 6851
rect 32873 6817 32907 6851
rect 32907 6817 32916 6851
rect 32864 6808 32916 6817
rect 35348 6808 35400 6860
rect 31300 6740 31352 6792
rect 33140 6740 33192 6792
rect 33968 6740 34020 6792
rect 34428 6783 34480 6792
rect 34428 6749 34437 6783
rect 34437 6749 34471 6783
rect 34471 6749 34480 6783
rect 34428 6740 34480 6749
rect 35440 6715 35492 6724
rect 20904 6604 20956 6656
rect 23020 6604 23072 6656
rect 35440 6681 35449 6715
rect 35449 6681 35483 6715
rect 35483 6681 35492 6715
rect 35440 6672 35492 6681
rect 36176 6740 36228 6792
rect 36912 6783 36964 6792
rect 36912 6749 36921 6783
rect 36921 6749 36955 6783
rect 36955 6749 36964 6783
rect 36912 6740 36964 6749
rect 30380 6647 30432 6656
rect 30380 6613 30389 6647
rect 30389 6613 30423 6647
rect 30423 6613 30432 6647
rect 30380 6604 30432 6613
rect 32680 6604 32732 6656
rect 35348 6604 35400 6656
rect 35992 6672 36044 6724
rect 36636 6672 36688 6724
rect 36268 6604 36320 6656
rect 4874 6502 4926 6554
rect 4938 6502 4990 6554
rect 5002 6502 5054 6554
rect 5066 6502 5118 6554
rect 5130 6502 5182 6554
rect 35594 6502 35646 6554
rect 35658 6502 35710 6554
rect 35722 6502 35774 6554
rect 35786 6502 35838 6554
rect 35850 6502 35902 6554
rect 12992 6400 13044 6452
rect 13636 6332 13688 6384
rect 14740 6400 14792 6452
rect 14924 6375 14976 6384
rect 14924 6341 14933 6375
rect 14933 6341 14967 6375
rect 14967 6341 14976 6375
rect 14924 6332 14976 6341
rect 14004 6264 14056 6316
rect 14096 6307 14148 6316
rect 14096 6273 14105 6307
rect 14105 6273 14139 6307
rect 14139 6273 14148 6307
rect 14096 6264 14148 6273
rect 14556 6307 14608 6316
rect 14556 6273 14565 6307
rect 14565 6273 14599 6307
rect 14599 6273 14608 6307
rect 14556 6264 14608 6273
rect 12072 6239 12124 6248
rect 12072 6205 12081 6239
rect 12081 6205 12115 6239
rect 12115 6205 12124 6239
rect 12072 6196 12124 6205
rect 12992 6196 13044 6248
rect 14832 6307 14884 6316
rect 14832 6273 14841 6307
rect 14841 6273 14875 6307
rect 14875 6273 14884 6307
rect 14832 6264 14884 6273
rect 15384 6264 15436 6316
rect 20444 6400 20496 6452
rect 20720 6400 20772 6452
rect 21364 6400 21416 6452
rect 19984 6332 20036 6384
rect 20628 6332 20680 6384
rect 16856 6264 16908 6316
rect 17408 6307 17460 6316
rect 17408 6273 17417 6307
rect 17417 6273 17451 6307
rect 17451 6273 17460 6307
rect 17408 6264 17460 6273
rect 14740 6128 14792 6180
rect 15844 6239 15896 6248
rect 15844 6205 15853 6239
rect 15853 6205 15887 6239
rect 15887 6205 15896 6239
rect 15844 6196 15896 6205
rect 17684 6239 17736 6248
rect 17684 6205 17693 6239
rect 17693 6205 17727 6239
rect 17727 6205 17736 6239
rect 17684 6196 17736 6205
rect 19156 6239 19208 6248
rect 19156 6205 19165 6239
rect 19165 6205 19199 6239
rect 19199 6205 19208 6239
rect 19156 6196 19208 6205
rect 20812 6264 20864 6316
rect 20996 6332 21048 6384
rect 21916 6332 21968 6384
rect 30380 6443 30432 6452
rect 30380 6409 30389 6443
rect 30389 6409 30423 6443
rect 30423 6409 30432 6443
rect 30380 6400 30432 6409
rect 36360 6400 36412 6452
rect 34796 6332 34848 6384
rect 35348 6332 35400 6384
rect 20628 6196 20680 6248
rect 19708 6128 19760 6180
rect 20904 6128 20956 6180
rect 21364 6239 21416 6248
rect 21364 6205 21373 6239
rect 21373 6205 21407 6239
rect 21407 6205 21416 6239
rect 21364 6196 21416 6205
rect 27436 6264 27488 6316
rect 29460 6264 29512 6316
rect 31852 6264 31904 6316
rect 34520 6264 34572 6316
rect 36176 6307 36228 6316
rect 36176 6273 36184 6307
rect 36184 6273 36218 6307
rect 36218 6273 36228 6307
rect 36176 6264 36228 6273
rect 36268 6307 36320 6316
rect 36268 6273 36277 6307
rect 36277 6273 36311 6307
rect 36311 6273 36320 6307
rect 36268 6264 36320 6273
rect 23296 6239 23348 6248
rect 23296 6205 23305 6239
rect 23305 6205 23339 6239
rect 23339 6205 23348 6239
rect 23296 6196 23348 6205
rect 23572 6239 23624 6248
rect 23572 6205 23581 6239
rect 23581 6205 23615 6239
rect 23615 6205 23624 6239
rect 23572 6196 23624 6205
rect 27804 6196 27856 6248
rect 28632 6239 28684 6248
rect 28632 6205 28641 6239
rect 28641 6205 28675 6239
rect 28675 6205 28684 6239
rect 28632 6196 28684 6205
rect 31392 6196 31444 6248
rect 31760 6196 31812 6248
rect 33784 6196 33836 6248
rect 33968 6239 34020 6248
rect 33968 6205 33977 6239
rect 33977 6205 34011 6239
rect 34011 6205 34020 6239
rect 33968 6196 34020 6205
rect 36636 6196 36688 6248
rect 12348 6060 12400 6112
rect 13912 6103 13964 6112
rect 13912 6069 13921 6103
rect 13921 6069 13955 6103
rect 13955 6069 13964 6103
rect 13912 6060 13964 6069
rect 14280 6060 14332 6112
rect 15752 6103 15804 6112
rect 15752 6069 15761 6103
rect 15761 6069 15795 6103
rect 15795 6069 15804 6103
rect 15752 6060 15804 6069
rect 17500 6103 17552 6112
rect 17500 6069 17509 6103
rect 17509 6069 17543 6103
rect 17543 6069 17552 6103
rect 17500 6060 17552 6069
rect 21088 6060 21140 6112
rect 21364 6060 21416 6112
rect 27896 6060 27948 6112
rect 29184 6103 29236 6112
rect 29184 6069 29193 6103
rect 29193 6069 29227 6103
rect 29227 6069 29236 6103
rect 29184 6060 29236 6069
rect 37004 6103 37056 6112
rect 37004 6069 37013 6103
rect 37013 6069 37047 6103
rect 37047 6069 37056 6103
rect 37004 6060 37056 6069
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 12992 5899 13044 5908
rect 12992 5865 13001 5899
rect 13001 5865 13035 5899
rect 13035 5865 13044 5899
rect 12992 5856 13044 5865
rect 14556 5899 14608 5908
rect 14556 5865 14565 5899
rect 14565 5865 14599 5899
rect 14599 5865 14608 5899
rect 14556 5856 14608 5865
rect 14832 5899 14884 5908
rect 14832 5865 14841 5899
rect 14841 5865 14875 5899
rect 14875 5865 14884 5899
rect 14832 5856 14884 5865
rect 18144 5899 18196 5908
rect 18144 5865 18153 5899
rect 18153 5865 18187 5899
rect 18187 5865 18196 5899
rect 18144 5856 18196 5865
rect 19156 5856 19208 5908
rect 20536 5856 20588 5908
rect 21364 5856 21416 5908
rect 23296 5856 23348 5908
rect 27436 5899 27488 5908
rect 27436 5865 27445 5899
rect 27445 5865 27479 5899
rect 27479 5865 27488 5899
rect 27436 5856 27488 5865
rect 29276 5899 29328 5908
rect 29276 5865 29285 5899
rect 29285 5865 29319 5899
rect 29319 5865 29328 5899
rect 29276 5856 29328 5865
rect 31852 5899 31904 5908
rect 31852 5865 31861 5899
rect 31861 5865 31895 5899
rect 31895 5865 31904 5899
rect 31852 5856 31904 5865
rect 34520 5899 34572 5908
rect 34520 5865 34529 5899
rect 34529 5865 34563 5899
rect 34563 5865 34572 5899
rect 34520 5856 34572 5865
rect 36176 5856 36228 5908
rect 12900 5652 12952 5704
rect 13912 5652 13964 5704
rect 14004 5652 14056 5704
rect 15384 5788 15436 5840
rect 14280 5695 14332 5704
rect 14280 5661 14289 5695
rect 14289 5661 14323 5695
rect 14323 5661 14332 5695
rect 14280 5652 14332 5661
rect 15752 5720 15804 5772
rect 15844 5763 15896 5772
rect 15844 5729 15853 5763
rect 15853 5729 15887 5763
rect 15887 5729 15896 5763
rect 15844 5720 15896 5729
rect 14556 5627 14608 5636
rect 14556 5593 14583 5627
rect 14583 5593 14608 5627
rect 16580 5652 16632 5704
rect 14556 5584 14608 5593
rect 14740 5627 14792 5636
rect 14740 5593 14749 5627
rect 14749 5593 14783 5627
rect 14783 5593 14792 5627
rect 16488 5627 16540 5636
rect 14740 5584 14792 5593
rect 16488 5593 16497 5627
rect 16497 5593 16531 5627
rect 16531 5593 16540 5627
rect 16488 5584 16540 5593
rect 16948 5652 17000 5704
rect 17776 5695 17828 5704
rect 17776 5661 17785 5695
rect 17785 5661 17819 5695
rect 17819 5661 17828 5695
rect 17776 5652 17828 5661
rect 16856 5584 16908 5636
rect 17500 5584 17552 5636
rect 19616 5720 19668 5772
rect 19984 5720 20036 5772
rect 20720 5720 20772 5772
rect 20996 5720 21048 5772
rect 21088 5763 21140 5772
rect 21088 5729 21097 5763
rect 21097 5729 21131 5763
rect 21131 5729 21140 5763
rect 21088 5720 21140 5729
rect 36636 5899 36688 5908
rect 36636 5865 36645 5899
rect 36645 5865 36679 5899
rect 36679 5865 36688 5899
rect 36636 5856 36688 5865
rect 37372 5856 37424 5908
rect 21272 5695 21324 5704
rect 21272 5661 21281 5695
rect 21281 5661 21315 5695
rect 21315 5661 21324 5695
rect 21272 5652 21324 5661
rect 24768 5652 24820 5704
rect 27896 5695 27948 5704
rect 27896 5661 27905 5695
rect 27905 5661 27939 5695
rect 27939 5661 27948 5695
rect 27896 5652 27948 5661
rect 29184 5652 29236 5704
rect 31852 5652 31904 5704
rect 32772 5695 32824 5704
rect 32772 5661 32781 5695
rect 32781 5661 32815 5695
rect 32815 5661 32824 5695
rect 32772 5652 32824 5661
rect 19432 5584 19484 5636
rect 13820 5516 13872 5568
rect 16212 5559 16264 5568
rect 16212 5525 16221 5559
rect 16221 5525 16255 5559
rect 16255 5525 16264 5559
rect 16212 5516 16264 5525
rect 19984 5584 20036 5636
rect 27620 5584 27672 5636
rect 30380 5627 30432 5636
rect 30380 5593 30389 5627
rect 30389 5593 30423 5627
rect 30423 5593 30432 5627
rect 30380 5584 30432 5593
rect 30472 5584 30524 5636
rect 27896 5516 27948 5568
rect 28080 5516 28132 5568
rect 28724 5516 28776 5568
rect 33324 5584 33376 5636
rect 36268 5652 36320 5704
rect 31944 5559 31996 5568
rect 31944 5525 31953 5559
rect 31953 5525 31987 5559
rect 31987 5525 31996 5559
rect 31944 5516 31996 5525
rect 32864 5516 32916 5568
rect 37832 5584 37884 5636
rect 34704 5559 34756 5568
rect 34704 5525 34713 5559
rect 34713 5525 34747 5559
rect 34747 5525 34756 5559
rect 34704 5516 34756 5525
rect 36176 5559 36228 5568
rect 36176 5525 36185 5559
rect 36185 5525 36219 5559
rect 36219 5525 36228 5559
rect 36176 5516 36228 5525
rect 4874 5414 4926 5466
rect 4938 5414 4990 5466
rect 5002 5414 5054 5466
rect 5066 5414 5118 5466
rect 5130 5414 5182 5466
rect 35594 5414 35646 5466
rect 35658 5414 35710 5466
rect 35722 5414 35774 5466
rect 35786 5414 35838 5466
rect 35850 5414 35902 5466
rect 13544 5244 13596 5296
rect 14556 5355 14608 5364
rect 14556 5321 14565 5355
rect 14565 5321 14599 5355
rect 14599 5321 14608 5355
rect 14556 5312 14608 5321
rect 14740 5355 14792 5364
rect 14740 5321 14749 5355
rect 14749 5321 14783 5355
rect 14783 5321 14792 5355
rect 14740 5312 14792 5321
rect 15292 5312 15344 5364
rect 15568 5312 15620 5364
rect 12348 5176 12400 5228
rect 13820 5108 13872 5160
rect 16212 5287 16264 5296
rect 16212 5253 16221 5287
rect 16221 5253 16255 5287
rect 16255 5253 16264 5287
rect 16212 5244 16264 5253
rect 16580 5312 16632 5364
rect 19432 5312 19484 5364
rect 23572 5244 23624 5296
rect 24768 5312 24820 5364
rect 26240 5312 26292 5364
rect 27620 5312 27672 5364
rect 27804 5312 27856 5364
rect 28172 5312 28224 5364
rect 29460 5355 29512 5364
rect 29460 5321 29469 5355
rect 29469 5321 29503 5355
rect 29503 5321 29512 5355
rect 29460 5312 29512 5321
rect 30380 5312 30432 5364
rect 31944 5312 31996 5364
rect 33324 5355 33376 5364
rect 33324 5321 33333 5355
rect 33333 5321 33367 5355
rect 33367 5321 33376 5355
rect 33324 5312 33376 5321
rect 34704 5312 34756 5364
rect 36268 5312 36320 5364
rect 16580 5176 16632 5228
rect 16856 5219 16908 5228
rect 16856 5185 16865 5219
rect 16865 5185 16899 5219
rect 16899 5185 16908 5219
rect 16856 5176 16908 5185
rect 17316 5176 17368 5228
rect 20536 5219 20588 5228
rect 20536 5185 20545 5219
rect 20545 5185 20579 5219
rect 20579 5185 20588 5219
rect 20536 5176 20588 5185
rect 26056 5244 26108 5296
rect 28080 5244 28132 5296
rect 31668 5244 31720 5296
rect 16120 5108 16172 5160
rect 23940 5151 23992 5160
rect 23940 5117 23949 5151
rect 23949 5117 23983 5151
rect 23983 5117 23992 5151
rect 23940 5108 23992 5117
rect 31392 5151 31444 5160
rect 31392 5117 31401 5151
rect 31401 5117 31435 5151
rect 31435 5117 31444 5151
rect 31392 5108 31444 5117
rect 37372 5312 37424 5364
rect 37004 5244 37056 5296
rect 33784 5151 33836 5160
rect 33784 5117 33793 5151
rect 33793 5117 33827 5151
rect 33827 5117 33836 5151
rect 33784 5108 33836 5117
rect 37096 5176 37148 5228
rect 34152 5151 34204 5160
rect 34152 5117 34161 5151
rect 34161 5117 34195 5151
rect 34195 5117 34204 5151
rect 34152 5108 34204 5117
rect 28080 4972 28132 5024
rect 34796 5015 34848 5024
rect 34796 4981 34805 5015
rect 34805 4981 34839 5015
rect 34839 4981 34848 5015
rect 34796 4972 34848 4981
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 17776 4768 17828 4820
rect 23940 4768 23992 4820
rect 26148 4811 26200 4820
rect 26148 4777 26157 4811
rect 26157 4777 26191 4811
rect 26191 4777 26200 4811
rect 26148 4768 26200 4777
rect 27712 4811 27764 4820
rect 27712 4777 27721 4811
rect 27721 4777 27755 4811
rect 27755 4777 27764 4811
rect 27712 4768 27764 4777
rect 34152 4768 34204 4820
rect 34612 4768 34664 4820
rect 34796 4768 34848 4820
rect 36176 4768 36228 4820
rect 15568 4675 15620 4684
rect 15568 4641 15577 4675
rect 15577 4641 15611 4675
rect 15611 4641 15620 4675
rect 15568 4632 15620 4641
rect 21916 4632 21968 4684
rect 24768 4632 24820 4684
rect 31484 4675 31536 4684
rect 31484 4641 31493 4675
rect 31493 4641 31527 4675
rect 31527 4641 31536 4675
rect 31484 4632 31536 4641
rect 32772 4632 32824 4684
rect 16120 4496 16172 4548
rect 22928 4496 22980 4548
rect 23388 4496 23440 4548
rect 27712 4564 27764 4616
rect 30748 4564 30800 4616
rect 32864 4564 32916 4616
rect 24676 4539 24728 4548
rect 24676 4505 24685 4539
rect 24685 4505 24719 4539
rect 24719 4505 24728 4539
rect 24676 4496 24728 4505
rect 26056 4496 26108 4548
rect 27804 4496 27856 4548
rect 28080 4539 28132 4548
rect 28080 4505 28089 4539
rect 28089 4505 28123 4539
rect 28123 4505 28132 4539
rect 28080 4496 28132 4505
rect 34612 4496 34664 4548
rect 16672 4428 16724 4480
rect 17316 4471 17368 4480
rect 17316 4437 17325 4471
rect 17325 4437 17359 4471
rect 17359 4437 17368 4471
rect 17316 4428 17368 4437
rect 19984 4428 20036 4480
rect 21180 4428 21232 4480
rect 23204 4471 23256 4480
rect 23204 4437 23213 4471
rect 23213 4437 23247 4471
rect 23247 4437 23256 4471
rect 23204 4428 23256 4437
rect 4874 4326 4926 4378
rect 4938 4326 4990 4378
rect 5002 4326 5054 4378
rect 5066 4326 5118 4378
rect 5130 4326 5182 4378
rect 35594 4326 35646 4378
rect 35658 4326 35710 4378
rect 35722 4326 35774 4378
rect 35786 4326 35838 4378
rect 35850 4326 35902 4378
rect 23204 4224 23256 4276
rect 19984 4199 20036 4208
rect 19984 4165 19993 4199
rect 19993 4165 20027 4199
rect 20027 4165 20036 4199
rect 19984 4156 20036 4165
rect 20720 4156 20772 4208
rect 23480 4156 23532 4208
rect 26056 4156 26108 4208
rect 16672 4131 16724 4140
rect 16672 4097 16681 4131
rect 16681 4097 16715 4131
rect 16715 4097 16724 4131
rect 16672 4088 16724 4097
rect 17316 4131 17368 4140
rect 17316 4097 17325 4131
rect 17325 4097 17359 4131
rect 17359 4097 17368 4131
rect 17316 4088 17368 4097
rect 22560 4131 22612 4140
rect 22560 4097 22569 4131
rect 22569 4097 22603 4131
rect 22603 4097 22612 4131
rect 22560 4088 22612 4097
rect 22928 4131 22980 4140
rect 22928 4097 22937 4131
rect 22937 4097 22971 4131
rect 22971 4097 22980 4131
rect 22928 4088 22980 4097
rect 23112 4131 23164 4140
rect 23112 4097 23121 4131
rect 23121 4097 23155 4131
rect 23155 4097 23164 4131
rect 23112 4088 23164 4097
rect 25320 4088 25372 4140
rect 26516 4131 26568 4140
rect 26516 4097 26525 4131
rect 26525 4097 26559 4131
rect 26559 4097 26568 4131
rect 26516 4088 26568 4097
rect 27804 4156 27856 4208
rect 19708 4063 19760 4072
rect 19708 4029 19717 4063
rect 19717 4029 19751 4063
rect 19751 4029 19760 4063
rect 19708 4020 19760 4029
rect 21364 4020 21416 4072
rect 21916 4020 21968 4072
rect 23388 4020 23440 4072
rect 22008 3952 22060 4004
rect 23756 4063 23808 4072
rect 23756 4029 23765 4063
rect 23765 4029 23799 4063
rect 23799 4029 23808 4063
rect 23756 4020 23808 4029
rect 21364 3884 21416 3936
rect 21548 3884 21600 3936
rect 22836 3927 22888 3936
rect 22836 3893 22845 3927
rect 22845 3893 22879 3927
rect 22879 3893 22888 3927
rect 22836 3884 22888 3893
rect 23296 3884 23348 3936
rect 25964 3884 26016 3936
rect 28724 4063 28776 4072
rect 28724 4029 28733 4063
rect 28733 4029 28767 4063
rect 28767 4029 28776 4063
rect 28724 4020 28776 4029
rect 27988 3884 28040 3936
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 24676 3680 24728 3732
rect 25320 3723 25372 3732
rect 25320 3689 25329 3723
rect 25329 3689 25363 3723
rect 25363 3689 25372 3723
rect 25320 3680 25372 3689
rect 25780 3680 25832 3732
rect 26516 3680 26568 3732
rect 23480 3655 23532 3664
rect 23480 3621 23489 3655
rect 23489 3621 23523 3655
rect 23523 3621 23532 3655
rect 23480 3612 23532 3621
rect 27896 3680 27948 3732
rect 30748 3680 30800 3732
rect 31392 3680 31444 3732
rect 19708 3587 19760 3596
rect 19708 3553 19717 3587
rect 19717 3553 19751 3587
rect 19751 3553 19760 3587
rect 19708 3544 19760 3553
rect 19984 3451 20036 3460
rect 19984 3417 19993 3451
rect 19993 3417 20027 3451
rect 20027 3417 20036 3451
rect 19984 3408 20036 3417
rect 20720 3408 20772 3460
rect 21824 3408 21876 3460
rect 23940 3544 23992 3596
rect 24768 3544 24820 3596
rect 28080 3544 28132 3596
rect 30380 3544 30432 3596
rect 31484 3544 31536 3596
rect 23388 3519 23440 3528
rect 23388 3485 23397 3519
rect 23397 3485 23431 3519
rect 23431 3485 23440 3519
rect 23388 3476 23440 3485
rect 22928 3408 22980 3460
rect 21916 3383 21968 3392
rect 21916 3349 21925 3383
rect 21925 3349 21959 3383
rect 21959 3349 21968 3383
rect 21916 3340 21968 3349
rect 22652 3340 22704 3392
rect 23296 3340 23348 3392
rect 23388 3340 23440 3392
rect 25688 3476 25740 3528
rect 25780 3519 25832 3528
rect 25780 3485 25789 3519
rect 25789 3485 25823 3519
rect 25823 3485 25832 3519
rect 25780 3476 25832 3485
rect 25964 3519 26016 3528
rect 25964 3485 25973 3519
rect 25973 3485 26007 3519
rect 26007 3485 26016 3519
rect 25964 3476 26016 3485
rect 29368 3476 29420 3528
rect 30288 3519 30340 3528
rect 30288 3485 30297 3519
rect 30297 3485 30331 3519
rect 30331 3485 30340 3519
rect 30288 3476 30340 3485
rect 27804 3408 27856 3460
rect 28816 3408 28868 3460
rect 30564 3408 30616 3460
rect 32312 3408 32364 3460
rect 32864 3408 32916 3460
rect 28356 3340 28408 3392
rect 32404 3340 32456 3392
rect 4874 3238 4926 3290
rect 4938 3238 4990 3290
rect 5002 3238 5054 3290
rect 5066 3238 5118 3290
rect 5130 3238 5182 3290
rect 35594 3238 35646 3290
rect 35658 3238 35710 3290
rect 35722 3238 35774 3290
rect 35786 3238 35838 3290
rect 35850 3238 35902 3290
rect 19984 3136 20036 3188
rect 22192 3136 22244 3188
rect 22560 3136 22612 3188
rect 23296 3136 23348 3188
rect 23756 3179 23808 3188
rect 23756 3145 23765 3179
rect 23765 3145 23799 3179
rect 23799 3145 23808 3179
rect 23756 3136 23808 3145
rect 25688 3179 25740 3188
rect 25688 3145 25697 3179
rect 25697 3145 25731 3179
rect 25731 3145 25740 3179
rect 25688 3136 25740 3145
rect 28080 3136 28132 3188
rect 22652 3111 22704 3120
rect 22652 3077 22661 3111
rect 22661 3077 22695 3111
rect 22695 3077 22704 3111
rect 22652 3068 22704 3077
rect 22836 3068 22888 3120
rect 26056 3068 26108 3120
rect 21916 3000 21968 3052
rect 23940 3043 23992 3052
rect 23940 3009 23949 3043
rect 23949 3009 23983 3043
rect 23983 3009 23992 3043
rect 23940 3000 23992 3009
rect 28356 3111 28408 3120
rect 28356 3077 28365 3111
rect 28365 3077 28399 3111
rect 28399 3077 28408 3111
rect 28356 3068 28408 3077
rect 28816 3068 28868 3120
rect 32680 3136 32732 3188
rect 33784 3136 33836 3188
rect 30380 3068 30432 3120
rect 32312 3068 32364 3120
rect 32404 3111 32456 3120
rect 32404 3077 32413 3111
rect 32413 3077 32447 3111
rect 32447 3077 32456 3111
rect 32404 3068 32456 3077
rect 32864 3068 32916 3120
rect 21180 2975 21232 2984
rect 21180 2941 21189 2975
rect 21189 2941 21223 2975
rect 21223 2941 21232 2975
rect 21180 2932 21232 2941
rect 21548 2932 21600 2984
rect 21824 2975 21876 2984
rect 21824 2941 21833 2975
rect 21833 2941 21867 2975
rect 21867 2941 21876 2975
rect 21824 2932 21876 2941
rect 22192 2864 22244 2916
rect 22928 2932 22980 2984
rect 23296 2975 23348 2984
rect 23296 2941 23305 2975
rect 23305 2941 23339 2975
rect 23339 2941 23348 2975
rect 23296 2932 23348 2941
rect 29000 2932 29052 2984
rect 31484 2932 31536 2984
rect 35348 3000 35400 3052
rect 37280 3043 37332 3052
rect 37280 3009 37289 3043
rect 37289 3009 37323 3043
rect 37323 3009 37332 3043
rect 37280 3000 37332 3009
rect 42432 3043 42484 3052
rect 42432 3009 42441 3043
rect 42441 3009 42475 3043
rect 42475 3009 42484 3043
rect 42432 3000 42484 3009
rect 43628 3043 43680 3052
rect 43628 3009 43637 3043
rect 43637 3009 43671 3043
rect 43671 3009 43680 3043
rect 43628 3000 43680 3009
rect 23388 2864 23440 2916
rect 30656 2796 30708 2848
rect 34152 2796 34204 2848
rect 34796 2796 34848 2848
rect 35440 2839 35492 2848
rect 35440 2805 35449 2839
rect 35449 2805 35483 2839
rect 35483 2805 35492 2839
rect 35440 2796 35492 2805
rect 36084 2796 36136 2848
rect 36728 2796 36780 2848
rect 37372 2796 37424 2848
rect 38016 2796 38068 2848
rect 38660 2796 38712 2848
rect 39304 2796 39356 2848
rect 39948 2796 40000 2848
rect 40592 2796 40644 2848
rect 41236 2796 41288 2848
rect 41880 2796 41932 2848
rect 42524 2796 42576 2848
rect 43168 2796 43220 2848
rect 43812 2839 43864 2848
rect 43812 2805 43821 2839
rect 43821 2805 43855 2839
rect 43855 2805 43864 2839
rect 43812 2796 43864 2805
rect 44456 2796 44508 2848
rect 45100 2796 45152 2848
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 19340 2592 19392 2644
rect 29000 2592 29052 2644
rect 29368 2635 29420 2644
rect 29368 2601 29377 2635
rect 29377 2601 29411 2635
rect 29411 2601 29420 2635
rect 29368 2592 29420 2601
rect 30104 2592 30156 2644
rect 30288 2592 30340 2644
rect 22560 2524 22612 2576
rect 30380 2524 30432 2576
rect 21824 2456 21876 2508
rect 22192 2431 22244 2440
rect 22192 2397 22201 2431
rect 22201 2397 22235 2431
rect 22235 2397 22244 2431
rect 22192 2388 22244 2397
rect 23296 2456 23348 2508
rect 21364 2320 21416 2372
rect 22652 2320 22704 2372
rect 23388 2388 23440 2440
rect 29000 2456 29052 2508
rect 19340 2295 19392 2304
rect 19340 2261 19349 2295
rect 19349 2261 19383 2295
rect 19383 2261 19392 2295
rect 19340 2252 19392 2261
rect 20628 2252 20680 2304
rect 21272 2252 21324 2304
rect 23204 2252 23256 2304
rect 29644 2320 29696 2372
rect 30104 2431 30156 2440
rect 30104 2397 30113 2431
rect 30113 2397 30147 2431
rect 30147 2397 30156 2431
rect 30104 2388 30156 2397
rect 30288 2431 30340 2440
rect 30288 2397 30297 2431
rect 30297 2397 30331 2431
rect 30331 2397 30340 2431
rect 30288 2388 30340 2397
rect 30748 2388 30800 2440
rect 35348 2499 35400 2508
rect 35348 2465 35357 2499
rect 35357 2465 35391 2499
rect 35391 2465 35400 2499
rect 35348 2456 35400 2465
rect 37280 2499 37332 2508
rect 37280 2465 37289 2499
rect 37289 2465 37323 2499
rect 37323 2465 37332 2499
rect 37280 2456 37332 2465
rect 42432 2499 42484 2508
rect 42432 2465 42441 2499
rect 42441 2465 42475 2499
rect 42475 2465 42484 2499
rect 42432 2456 42484 2465
rect 43628 2499 43680 2508
rect 43628 2465 43637 2499
rect 43637 2465 43671 2499
rect 43671 2465 43680 2499
rect 43628 2456 43680 2465
rect 30288 2252 30340 2304
rect 30932 2252 30984 2304
rect 4874 2150 4926 2202
rect 4938 2150 4990 2202
rect 5002 2150 5054 2202
rect 5066 2150 5118 2202
rect 5130 2150 5182 2202
rect 35594 2150 35646 2202
rect 35658 2150 35710 2202
rect 35722 2150 35774 2202
rect 35786 2150 35838 2202
rect 35850 2150 35902 2202
<< metal2 >>
rect 22558 39200 22614 40000
rect 23202 39200 23258 40000
rect 24490 39200 24546 40000
rect 25134 39200 25190 40000
rect 25778 39200 25834 40000
rect 26422 39200 26478 40000
rect 27066 39200 27122 40000
rect 27710 39200 27766 40000
rect 28354 39200 28410 40000
rect 28998 39200 29054 40000
rect 29642 39200 29698 40000
rect 30286 39200 30342 40000
rect 30930 39200 30986 40000
rect 31574 39200 31630 40000
rect 32218 39200 32274 40000
rect 32862 39200 32918 40000
rect 33506 39200 33562 40000
rect 34150 39200 34206 40000
rect 34794 39200 34850 40000
rect 35438 39200 35494 40000
rect 36082 39200 36138 40000
rect 36726 39200 36782 40000
rect 37370 39200 37426 40000
rect 38014 39200 38070 40000
rect 38658 39200 38714 40000
rect 39302 39200 39358 40000
rect 39946 39200 40002 40000
rect 40590 39200 40646 40000
rect 41234 39200 41290 40000
rect 41878 39200 41934 40000
rect 42522 39200 42578 40000
rect 43166 39200 43222 40000
rect 43810 39200 43866 40000
rect 44454 39200 44510 40000
rect 45098 39200 45154 40000
rect 45742 39200 45798 40000
rect 46386 39200 46442 40000
rect 47030 39200 47086 40000
rect 47674 39200 47730 40000
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37499 4522 37508
rect 22572 37466 22600 39200
rect 23216 37466 23244 39200
rect 22560 37460 22612 37466
rect 22560 37402 22612 37408
rect 23204 37460 23256 37466
rect 23204 37402 23256 37408
rect 23020 37188 23072 37194
rect 23020 37130 23072 37136
rect 24216 37188 24268 37194
rect 24216 37130 24268 37136
rect 4874 37020 5182 37029
rect 4874 37018 4880 37020
rect 4936 37018 4960 37020
rect 5016 37018 5040 37020
rect 5096 37018 5120 37020
rect 5176 37018 5182 37020
rect 4936 36966 4938 37018
rect 5118 36966 5120 37018
rect 4874 36964 4880 36966
rect 4936 36964 4960 36966
rect 5016 36964 5040 36966
rect 5096 36964 5120 36966
rect 5176 36964 5182 36966
rect 4874 36955 5182 36964
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 22100 36168 22152 36174
rect 22100 36110 22152 36116
rect 4874 35932 5182 35941
rect 4874 35930 4880 35932
rect 4936 35930 4960 35932
rect 5016 35930 5040 35932
rect 5096 35930 5120 35932
rect 5176 35930 5182 35932
rect 4936 35878 4938 35930
rect 5118 35878 5120 35930
rect 4874 35876 4880 35878
rect 4936 35876 4960 35878
rect 5016 35876 5040 35878
rect 5096 35876 5120 35878
rect 5176 35876 5182 35878
rect 4874 35867 5182 35876
rect 21916 35692 21968 35698
rect 21916 35634 21968 35640
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 21928 35290 21956 35634
rect 22112 35494 22140 36110
rect 23032 35834 23060 37130
rect 24228 36378 24256 37130
rect 24504 36922 24532 39200
rect 25148 36922 25176 39200
rect 25792 36922 25820 39200
rect 26436 37466 26464 39200
rect 26424 37460 26476 37466
rect 26424 37402 26476 37408
rect 27080 36922 27108 39200
rect 27724 36922 27752 39200
rect 28368 37466 28396 39200
rect 28356 37460 28408 37466
rect 28356 37402 28408 37408
rect 29012 36922 29040 39200
rect 29656 36922 29684 39200
rect 29736 37188 29788 37194
rect 29736 37130 29788 37136
rect 24492 36916 24544 36922
rect 24492 36858 24544 36864
rect 25136 36916 25188 36922
rect 25136 36858 25188 36864
rect 25780 36916 25832 36922
rect 25780 36858 25832 36864
rect 27068 36916 27120 36922
rect 27068 36858 27120 36864
rect 27712 36916 27764 36922
rect 27712 36858 27764 36864
rect 29000 36916 29052 36922
rect 29000 36858 29052 36864
rect 29644 36916 29696 36922
rect 29644 36858 29696 36864
rect 25320 36780 25372 36786
rect 25320 36722 25372 36728
rect 25332 36378 25360 36722
rect 24216 36372 24268 36378
rect 24216 36314 24268 36320
rect 25320 36372 25372 36378
rect 25320 36314 25372 36320
rect 29748 36106 29776 37130
rect 30300 36922 30328 39200
rect 30944 36922 30972 39200
rect 31588 36922 31616 39200
rect 31668 37256 31720 37262
rect 31668 37198 31720 37204
rect 30288 36916 30340 36922
rect 30288 36858 30340 36864
rect 30932 36916 30984 36922
rect 30932 36858 30984 36864
rect 31576 36916 31628 36922
rect 31576 36858 31628 36864
rect 23296 36100 23348 36106
rect 23296 36042 23348 36048
rect 23572 36100 23624 36106
rect 23572 36042 23624 36048
rect 28816 36100 28868 36106
rect 28816 36042 28868 36048
rect 29736 36100 29788 36106
rect 29736 36042 29788 36048
rect 23308 35834 23336 36042
rect 23020 35828 23072 35834
rect 23020 35770 23072 35776
rect 23296 35828 23348 35834
rect 23296 35770 23348 35776
rect 22100 35488 22152 35494
rect 22100 35430 22152 35436
rect 21916 35284 21968 35290
rect 21916 35226 21968 35232
rect 18604 35080 18656 35086
rect 18604 35022 18656 35028
rect 16856 34944 16908 34950
rect 16856 34886 16908 34892
rect 4874 34844 5182 34853
rect 4874 34842 4880 34844
rect 4936 34842 4960 34844
rect 5016 34842 5040 34844
rect 5096 34842 5120 34844
rect 5176 34842 5182 34844
rect 4936 34790 4938 34842
rect 5118 34790 5120 34842
rect 4874 34788 4880 34790
rect 4936 34788 4960 34790
rect 5016 34788 5040 34790
rect 5096 34788 5120 34790
rect 5176 34788 5182 34790
rect 4874 34779 5182 34788
rect 16868 34610 16896 34886
rect 18052 34672 18104 34678
rect 18052 34614 18104 34620
rect 16856 34604 16908 34610
rect 16856 34546 16908 34552
rect 16948 34536 17000 34542
rect 16948 34478 17000 34484
rect 17224 34536 17276 34542
rect 18064 34524 18092 34614
rect 18616 34542 18644 35022
rect 21272 34604 21324 34610
rect 21272 34546 21324 34552
rect 17224 34478 17276 34484
rect 17972 34496 18092 34524
rect 18144 34536 18196 34542
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 16960 33862 16988 34478
rect 17132 33992 17184 33998
rect 17132 33934 17184 33940
rect 16948 33856 17000 33862
rect 16948 33798 17000 33804
rect 4874 33756 5182 33765
rect 4874 33754 4880 33756
rect 4936 33754 4960 33756
rect 5016 33754 5040 33756
rect 5096 33754 5120 33756
rect 5176 33754 5182 33756
rect 4936 33702 4938 33754
rect 5118 33702 5120 33754
rect 4874 33700 4880 33702
rect 4936 33700 4960 33702
rect 5016 33700 5040 33702
rect 5096 33700 5120 33702
rect 5176 33700 5182 33702
rect 4874 33691 5182 33700
rect 15936 33584 15988 33590
rect 15936 33526 15988 33532
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 13912 32904 13964 32910
rect 13912 32846 13964 32852
rect 4874 32668 5182 32677
rect 4874 32666 4880 32668
rect 4936 32666 4960 32668
rect 5016 32666 5040 32668
rect 5096 32666 5120 32668
rect 5176 32666 5182 32668
rect 4936 32614 4938 32666
rect 5118 32614 5120 32666
rect 4874 32612 4880 32614
rect 4936 32612 4960 32614
rect 5016 32612 5040 32614
rect 5096 32612 5120 32614
rect 5176 32612 5182 32614
rect 4874 32603 5182 32612
rect 13924 32502 13952 32846
rect 15948 32842 15976 33526
rect 16960 33522 16988 33798
rect 17144 33522 17172 33934
rect 16948 33516 17000 33522
rect 16948 33458 17000 33464
rect 17132 33516 17184 33522
rect 17132 33458 17184 33464
rect 17236 33454 17264 34478
rect 17868 33992 17920 33998
rect 17868 33934 17920 33940
rect 17776 33856 17828 33862
rect 17776 33798 17828 33804
rect 17224 33448 17276 33454
rect 17224 33390 17276 33396
rect 17040 33312 17092 33318
rect 17040 33254 17092 33260
rect 14648 32836 14700 32842
rect 14648 32778 14700 32784
rect 15936 32836 15988 32842
rect 15936 32778 15988 32784
rect 14660 32570 14688 32778
rect 14648 32564 14700 32570
rect 14648 32506 14700 32512
rect 13912 32496 13964 32502
rect 13912 32438 13964 32444
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 4874 31580 5182 31589
rect 4874 31578 4880 31580
rect 4936 31578 4960 31580
rect 5016 31578 5040 31580
rect 5096 31578 5120 31580
rect 5176 31578 5182 31580
rect 4936 31526 4938 31578
rect 5118 31526 5120 31578
rect 4874 31524 4880 31526
rect 4936 31524 4960 31526
rect 5016 31524 5040 31526
rect 5096 31524 5120 31526
rect 5176 31524 5182 31526
rect 4874 31515 5182 31524
rect 13924 31346 13952 32438
rect 15568 31816 15620 31822
rect 15568 31758 15620 31764
rect 15844 31816 15896 31822
rect 15844 31758 15896 31764
rect 15580 31482 15608 31758
rect 15568 31476 15620 31482
rect 15568 31418 15620 31424
rect 13912 31340 13964 31346
rect 13912 31282 13964 31288
rect 15856 31210 15884 31758
rect 15948 31414 15976 32778
rect 16304 32768 16356 32774
rect 16304 32710 16356 32716
rect 16488 32768 16540 32774
rect 16488 32710 16540 32716
rect 16316 32434 16344 32710
rect 16304 32428 16356 32434
rect 16304 32370 16356 32376
rect 16500 32026 16528 32710
rect 17052 32366 17080 33254
rect 17236 32858 17264 33390
rect 17236 32830 17356 32858
rect 17788 32842 17816 33798
rect 17880 32910 17908 33934
rect 17972 33590 18000 34496
rect 18144 34478 18196 34484
rect 18604 34536 18656 34542
rect 18604 34478 18656 34484
rect 18156 34202 18184 34478
rect 21180 34400 21232 34406
rect 21180 34342 21232 34348
rect 18144 34196 18196 34202
rect 18144 34138 18196 34144
rect 18052 34060 18104 34066
rect 18052 34002 18104 34008
rect 17960 33584 18012 33590
rect 17960 33526 18012 33532
rect 18064 33318 18092 34002
rect 18052 33312 18104 33318
rect 18052 33254 18104 33260
rect 18064 32910 18092 33254
rect 18156 32910 18184 34138
rect 20260 34128 20312 34134
rect 20260 34070 20312 34076
rect 19800 34060 19852 34066
rect 19800 34002 19852 34008
rect 18328 33856 18380 33862
rect 18328 33798 18380 33804
rect 18236 33448 18288 33454
rect 18236 33390 18288 33396
rect 18248 33114 18276 33390
rect 18236 33108 18288 33114
rect 18236 33050 18288 33056
rect 18340 33046 18368 33798
rect 18972 33312 19024 33318
rect 18972 33254 19024 33260
rect 18328 33040 18380 33046
rect 18328 32982 18380 32988
rect 18984 32978 19012 33254
rect 19812 33114 19840 34002
rect 20272 33590 20300 34070
rect 21192 33930 21220 34342
rect 21284 34202 21312 34546
rect 22112 34542 22140 35430
rect 22284 35284 22336 35290
rect 22284 35226 22336 35232
rect 22296 35086 22324 35226
rect 23032 35154 23060 35770
rect 23584 35698 23612 36042
rect 28828 35834 28856 36042
rect 29552 36032 29604 36038
rect 29552 35974 29604 35980
rect 25228 35828 25280 35834
rect 25228 35770 25280 35776
rect 28816 35828 28868 35834
rect 28816 35770 28868 35776
rect 23572 35692 23624 35698
rect 23572 35634 23624 35640
rect 23664 35692 23716 35698
rect 23664 35634 23716 35640
rect 23756 35692 23808 35698
rect 23756 35634 23808 35640
rect 23676 35290 23704 35634
rect 23664 35284 23716 35290
rect 23664 35226 23716 35232
rect 23020 35148 23072 35154
rect 23020 35090 23072 35096
rect 22284 35080 22336 35086
rect 22284 35022 22336 35028
rect 22468 35080 22520 35086
rect 22468 35022 22520 35028
rect 22652 35080 22704 35086
rect 22652 35022 22704 35028
rect 22100 34536 22152 34542
rect 22100 34478 22152 34484
rect 21272 34196 21324 34202
rect 21272 34138 21324 34144
rect 21640 34128 21692 34134
rect 21640 34070 21692 34076
rect 21180 33924 21232 33930
rect 21180 33866 21232 33872
rect 21652 33658 21680 34070
rect 22008 33992 22060 33998
rect 22008 33934 22060 33940
rect 21640 33652 21692 33658
rect 21640 33594 21692 33600
rect 20260 33584 20312 33590
rect 20260 33526 20312 33532
rect 22020 33522 22048 33934
rect 22008 33516 22060 33522
rect 22008 33458 22060 33464
rect 20628 33448 20680 33454
rect 20628 33390 20680 33396
rect 19800 33108 19852 33114
rect 19800 33050 19852 33056
rect 18972 32972 19024 32978
rect 18972 32914 19024 32920
rect 20640 32910 20668 33390
rect 21824 33312 21876 33318
rect 21824 33254 21876 33260
rect 21836 32978 21864 33254
rect 21824 32972 21876 32978
rect 21824 32914 21876 32920
rect 17868 32904 17920 32910
rect 17868 32846 17920 32852
rect 18052 32904 18104 32910
rect 18052 32846 18104 32852
rect 18144 32904 18196 32910
rect 18144 32846 18196 32852
rect 20628 32904 20680 32910
rect 20628 32846 20680 32852
rect 17328 32434 17356 32830
rect 17776 32836 17828 32842
rect 17776 32778 17828 32784
rect 18236 32836 18288 32842
rect 18236 32778 18288 32784
rect 18248 32722 18276 32778
rect 18156 32694 18276 32722
rect 19248 32768 19300 32774
rect 19248 32710 19300 32716
rect 17316 32428 17368 32434
rect 17316 32370 17368 32376
rect 17040 32360 17092 32366
rect 17040 32302 17092 32308
rect 16488 32020 16540 32026
rect 16488 31962 16540 31968
rect 16120 31680 16172 31686
rect 16120 31622 16172 31628
rect 15936 31408 15988 31414
rect 15936 31350 15988 31356
rect 15844 31204 15896 31210
rect 15844 31146 15896 31152
rect 15948 31142 15976 31350
rect 16132 31346 16160 31622
rect 16120 31340 16172 31346
rect 16120 31282 16172 31288
rect 16500 31278 16528 31962
rect 17328 31754 17356 32370
rect 17960 32224 18012 32230
rect 17960 32166 18012 32172
rect 17972 31822 18000 32166
rect 18156 32026 18184 32694
rect 18328 32224 18380 32230
rect 18328 32166 18380 32172
rect 18144 32020 18196 32026
rect 18144 31962 18196 31968
rect 17960 31816 18012 31822
rect 17960 31758 18012 31764
rect 17316 31748 17368 31754
rect 17316 31690 17368 31696
rect 16488 31272 16540 31278
rect 16488 31214 16540 31220
rect 17224 31272 17276 31278
rect 17224 31214 17276 31220
rect 15936 31136 15988 31142
rect 15936 31078 15988 31084
rect 16488 31136 16540 31142
rect 16488 31078 16540 31084
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 16500 30666 16528 31078
rect 17236 30938 17264 31214
rect 17224 30932 17276 30938
rect 17224 30874 17276 30880
rect 17328 30734 17356 31690
rect 18156 31482 18184 31962
rect 18236 31680 18288 31686
rect 18236 31622 18288 31628
rect 18144 31476 18196 31482
rect 18144 31418 18196 31424
rect 17868 31408 17920 31414
rect 17920 31368 18000 31396
rect 17868 31350 17920 31356
rect 17776 31136 17828 31142
rect 17776 31078 17828 31084
rect 17788 30734 17816 31078
rect 17316 30728 17368 30734
rect 17316 30670 17368 30676
rect 17776 30728 17828 30734
rect 17776 30670 17828 30676
rect 16488 30660 16540 30666
rect 16488 30602 16540 30608
rect 4874 30492 5182 30501
rect 4874 30490 4880 30492
rect 4936 30490 4960 30492
rect 5016 30490 5040 30492
rect 5096 30490 5120 30492
rect 5176 30490 5182 30492
rect 4936 30438 4938 30490
rect 5118 30438 5120 30490
rect 4874 30436 4880 30438
rect 4936 30436 4960 30438
rect 5016 30436 5040 30438
rect 5096 30436 5120 30438
rect 5176 30436 5182 30438
rect 4874 30427 5182 30436
rect 17328 30258 17356 30670
rect 17972 30598 18000 31368
rect 18248 30666 18276 31622
rect 18236 30660 18288 30666
rect 18236 30602 18288 30608
rect 17960 30592 18012 30598
rect 17960 30534 18012 30540
rect 17316 30252 17368 30258
rect 17316 30194 17368 30200
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 16856 29776 16908 29782
rect 16856 29718 16908 29724
rect 4874 29404 5182 29413
rect 4874 29402 4880 29404
rect 4936 29402 4960 29404
rect 5016 29402 5040 29404
rect 5096 29402 5120 29404
rect 5176 29402 5182 29404
rect 4936 29350 4938 29402
rect 5118 29350 5120 29402
rect 4874 29348 4880 29350
rect 4936 29348 4960 29350
rect 5016 29348 5040 29350
rect 5096 29348 5120 29350
rect 5176 29348 5182 29350
rect 4874 29339 5182 29348
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 4874 28316 5182 28325
rect 4874 28314 4880 28316
rect 4936 28314 4960 28316
rect 5016 28314 5040 28316
rect 5096 28314 5120 28316
rect 5176 28314 5182 28316
rect 4936 28262 4938 28314
rect 5118 28262 5120 28314
rect 4874 28260 4880 28262
rect 4936 28260 4960 28262
rect 5016 28260 5040 28262
rect 5096 28260 5120 28262
rect 5176 28260 5182 28262
rect 4874 28251 5182 28260
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 4874 27228 5182 27237
rect 4874 27226 4880 27228
rect 4936 27226 4960 27228
rect 5016 27226 5040 27228
rect 5096 27226 5120 27228
rect 5176 27226 5182 27228
rect 4936 27174 4938 27226
rect 5118 27174 5120 27226
rect 4874 27172 4880 27174
rect 4936 27172 4960 27174
rect 5016 27172 5040 27174
rect 5096 27172 5120 27174
rect 5176 27172 5182 27174
rect 4874 27163 5182 27172
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 4874 26140 5182 26149
rect 4874 26138 4880 26140
rect 4936 26138 4960 26140
rect 5016 26138 5040 26140
rect 5096 26138 5120 26140
rect 5176 26138 5182 26140
rect 4936 26086 4938 26138
rect 5118 26086 5120 26138
rect 4874 26084 4880 26086
rect 4936 26084 4960 26086
rect 5016 26084 5040 26086
rect 5096 26084 5120 26086
rect 5176 26084 5182 26086
rect 4874 26075 5182 26084
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 4874 25052 5182 25061
rect 4874 25050 4880 25052
rect 4936 25050 4960 25052
rect 5016 25050 5040 25052
rect 5096 25050 5120 25052
rect 5176 25050 5182 25052
rect 4936 24998 4938 25050
rect 5118 24998 5120 25050
rect 4874 24996 4880 24998
rect 4936 24996 4960 24998
rect 5016 24996 5040 24998
rect 5096 24996 5120 24998
rect 5176 24996 5182 24998
rect 4874 24987 5182 24996
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 4874 23964 5182 23973
rect 4874 23962 4880 23964
rect 4936 23962 4960 23964
rect 5016 23962 5040 23964
rect 5096 23962 5120 23964
rect 5176 23962 5182 23964
rect 4936 23910 4938 23962
rect 5118 23910 5120 23962
rect 4874 23908 4880 23910
rect 4936 23908 4960 23910
rect 5016 23908 5040 23910
rect 5096 23908 5120 23910
rect 5176 23908 5182 23910
rect 4874 23899 5182 23908
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 4874 22876 5182 22885
rect 4874 22874 4880 22876
rect 4936 22874 4960 22876
rect 5016 22874 5040 22876
rect 5096 22874 5120 22876
rect 5176 22874 5182 22876
rect 4936 22822 4938 22874
rect 5118 22822 5120 22874
rect 4874 22820 4880 22822
rect 4936 22820 4960 22822
rect 5016 22820 5040 22822
rect 5096 22820 5120 22822
rect 5176 22820 5182 22822
rect 4874 22811 5182 22820
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 4874 21788 5182 21797
rect 4874 21786 4880 21788
rect 4936 21786 4960 21788
rect 5016 21786 5040 21788
rect 5096 21786 5120 21788
rect 5176 21786 5182 21788
rect 4936 21734 4938 21786
rect 5118 21734 5120 21786
rect 4874 21732 4880 21734
rect 4936 21732 4960 21734
rect 5016 21732 5040 21734
rect 5096 21732 5120 21734
rect 5176 21732 5182 21734
rect 4874 21723 5182 21732
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 4874 20700 5182 20709
rect 4874 20698 4880 20700
rect 4936 20698 4960 20700
rect 5016 20698 5040 20700
rect 5096 20698 5120 20700
rect 5176 20698 5182 20700
rect 4936 20646 4938 20698
rect 5118 20646 5120 20698
rect 4874 20644 4880 20646
rect 4936 20644 4960 20646
rect 5016 20644 5040 20646
rect 5096 20644 5120 20646
rect 5176 20644 5182 20646
rect 4874 20635 5182 20644
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 15200 19848 15252 19854
rect 15200 19790 15252 19796
rect 848 19712 900 19718
rect 846 19680 848 19689
rect 900 19680 902 19689
rect 846 19615 902 19624
rect 4874 19612 5182 19621
rect 4874 19610 4880 19612
rect 4936 19610 4960 19612
rect 5016 19610 5040 19612
rect 5096 19610 5120 19612
rect 5176 19610 5182 19612
rect 4936 19558 4938 19610
rect 5118 19558 5120 19610
rect 4874 19556 4880 19558
rect 4936 19556 4960 19558
rect 5016 19556 5040 19558
rect 5096 19556 5120 19558
rect 5176 19556 5182 19558
rect 4874 19547 5182 19556
rect 15212 19514 15240 19790
rect 15200 19508 15252 19514
rect 15200 19450 15252 19456
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 15212 18834 15240 19450
rect 16120 19372 16172 19378
rect 16120 19314 16172 19320
rect 16672 19372 16724 19378
rect 16672 19314 16724 19320
rect 16132 18970 16160 19314
rect 16120 18964 16172 18970
rect 16120 18906 16172 18912
rect 15200 18828 15252 18834
rect 15200 18770 15252 18776
rect 4874 18524 5182 18533
rect 4874 18522 4880 18524
rect 4936 18522 4960 18524
rect 5016 18522 5040 18524
rect 5096 18522 5120 18524
rect 5176 18522 5182 18524
rect 4936 18470 4938 18522
rect 5118 18470 5120 18522
rect 4874 18468 4880 18470
rect 4936 18468 4960 18470
rect 5016 18468 5040 18470
rect 5096 18468 5120 18470
rect 5176 18468 5182 18470
rect 4874 18459 5182 18468
rect 16580 18284 16632 18290
rect 16580 18226 16632 18232
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 4874 17436 5182 17445
rect 4874 17434 4880 17436
rect 4936 17434 4960 17436
rect 5016 17434 5040 17436
rect 5096 17434 5120 17436
rect 5176 17434 5182 17436
rect 4936 17382 4938 17434
rect 5118 17382 5120 17434
rect 4874 17380 4880 17382
rect 4936 17380 4960 17382
rect 5016 17380 5040 17382
rect 5096 17380 5120 17382
rect 5176 17380 5182 17382
rect 4874 17371 5182 17380
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 4874 16348 5182 16357
rect 4874 16346 4880 16348
rect 4936 16346 4960 16348
rect 5016 16346 5040 16348
rect 5096 16346 5120 16348
rect 5176 16346 5182 16348
rect 4936 16294 4938 16346
rect 5118 16294 5120 16346
rect 4874 16292 4880 16294
rect 4936 16292 4960 16294
rect 5016 16292 5040 16294
rect 5096 16292 5120 16294
rect 5176 16292 5182 16294
rect 4874 16283 5182 16292
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 13268 15564 13320 15570
rect 13268 15506 13320 15512
rect 12624 15428 12676 15434
rect 12624 15370 12676 15376
rect 4874 15260 5182 15269
rect 4874 15258 4880 15260
rect 4936 15258 4960 15260
rect 5016 15258 5040 15260
rect 5096 15258 5120 15260
rect 5176 15258 5182 15260
rect 4936 15206 4938 15258
rect 5118 15206 5120 15258
rect 4874 15204 4880 15206
rect 4936 15204 4960 15206
rect 5016 15204 5040 15206
rect 5096 15204 5120 15206
rect 5176 15204 5182 15206
rect 4874 15195 5182 15204
rect 12636 15026 12664 15370
rect 12716 15360 12768 15366
rect 12716 15302 12768 15308
rect 12624 15020 12676 15026
rect 12624 14962 12676 14968
rect 12348 14816 12400 14822
rect 12348 14758 12400 14764
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 12360 14414 12388 14758
rect 12728 14482 12756 15302
rect 13280 15094 13308 15506
rect 14924 15496 14976 15502
rect 14924 15438 14976 15444
rect 13452 15428 13504 15434
rect 13452 15370 13504 15376
rect 13268 15088 13320 15094
rect 13268 15030 13320 15036
rect 12900 15020 12952 15026
rect 12900 14962 12952 14968
rect 12912 14618 12940 14962
rect 13464 14906 13492 15370
rect 14740 15020 14792 15026
rect 14740 14962 14792 14968
rect 13636 14952 13688 14958
rect 13464 14900 13636 14906
rect 13464 14894 13688 14900
rect 13464 14878 13676 14894
rect 12900 14612 12952 14618
rect 12900 14554 12952 14560
rect 13464 14482 13492 14878
rect 14752 14482 14780 14962
rect 14936 14822 14964 15438
rect 15108 15360 15160 15366
rect 15108 15302 15160 15308
rect 14924 14816 14976 14822
rect 14924 14758 14976 14764
rect 12716 14476 12768 14482
rect 12716 14418 12768 14424
rect 13176 14476 13228 14482
rect 13176 14418 13228 14424
rect 13452 14476 13504 14482
rect 13452 14418 13504 14424
rect 14740 14476 14792 14482
rect 14740 14418 14792 14424
rect 1216 14408 1268 14414
rect 1214 14376 1216 14385
rect 12348 14408 12400 14414
rect 1268 14376 1270 14385
rect 12348 14350 12400 14356
rect 1214 14311 1270 14320
rect 11704 14340 11756 14346
rect 11704 14282 11756 14288
rect 4874 14172 5182 14181
rect 4874 14170 4880 14172
rect 4936 14170 4960 14172
rect 5016 14170 5040 14172
rect 5096 14170 5120 14172
rect 5176 14170 5182 14172
rect 4936 14118 4938 14170
rect 5118 14118 5120 14170
rect 4874 14116 4880 14118
rect 4936 14116 4960 14118
rect 5016 14116 5040 14118
rect 5096 14116 5120 14118
rect 5176 14116 5182 14118
rect 4874 14107 5182 14116
rect 11716 14074 11744 14282
rect 12256 14272 12308 14278
rect 12256 14214 12308 14220
rect 11704 14068 11756 14074
rect 11704 14010 11756 14016
rect 12164 13864 12216 13870
rect 12164 13806 12216 13812
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 12176 13258 12204 13806
rect 12268 13394 12296 14214
rect 13188 14006 13216 14418
rect 13176 14000 13228 14006
rect 13176 13942 13228 13948
rect 13464 13530 13492 14418
rect 14752 13870 14780 14418
rect 13636 13864 13688 13870
rect 13636 13806 13688 13812
rect 14740 13864 14792 13870
rect 14740 13806 14792 13812
rect 13452 13524 13504 13530
rect 13452 13466 13504 13472
rect 12256 13388 12308 13394
rect 12256 13330 12308 13336
rect 13648 13258 13676 13806
rect 14752 13394 14780 13806
rect 14740 13388 14792 13394
rect 14740 13330 14792 13336
rect 14936 13326 14964 14758
rect 14924 13320 14976 13326
rect 14924 13262 14976 13268
rect 12164 13252 12216 13258
rect 12164 13194 12216 13200
rect 13636 13252 13688 13258
rect 13636 13194 13688 13200
rect 4874 13084 5182 13093
rect 4874 13082 4880 13084
rect 4936 13082 4960 13084
rect 5016 13082 5040 13084
rect 5096 13082 5120 13084
rect 5176 13082 5182 13084
rect 4936 13030 4938 13082
rect 5118 13030 5120 13082
rect 4874 13028 4880 13030
rect 4936 13028 4960 13030
rect 5016 13028 5040 13030
rect 5096 13028 5120 13030
rect 5176 13028 5182 13030
rect 4874 13019 5182 13028
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 12176 12306 12204 13194
rect 13648 12434 13676 13194
rect 15120 13190 15148 15302
rect 15476 14952 15528 14958
rect 15476 14894 15528 14900
rect 15200 14476 15252 14482
rect 15200 14418 15252 14424
rect 15212 13530 15240 14418
rect 15292 14408 15344 14414
rect 15292 14350 15344 14356
rect 15304 14074 15332 14350
rect 15488 14278 15516 14894
rect 16120 14816 16172 14822
rect 16120 14758 16172 14764
rect 15476 14272 15528 14278
rect 15476 14214 15528 14220
rect 15292 14068 15344 14074
rect 15292 14010 15344 14016
rect 15488 13938 15516 14214
rect 15476 13932 15528 13938
rect 15476 13874 15528 13880
rect 15200 13524 15252 13530
rect 15200 13466 15252 13472
rect 15660 13388 15712 13394
rect 15660 13330 15712 13336
rect 15108 13184 15160 13190
rect 15108 13126 15160 13132
rect 15384 12844 15436 12850
rect 15384 12786 15436 12792
rect 15396 12442 15424 12786
rect 13464 12406 13676 12434
rect 15384 12436 15436 12442
rect 12164 12300 12216 12306
rect 12164 12242 12216 12248
rect 4874 11996 5182 12005
rect 4874 11994 4880 11996
rect 4936 11994 4960 11996
rect 5016 11994 5040 11996
rect 5096 11994 5120 11996
rect 5176 11994 5182 11996
rect 4936 11942 4938 11994
rect 5118 11942 5120 11994
rect 4874 11940 4880 11942
rect 4936 11940 4960 11942
rect 5016 11940 5040 11942
rect 5096 11940 5120 11942
rect 5176 11940 5182 11942
rect 4874 11931 5182 11940
rect 12176 11762 12204 12242
rect 13464 12170 13492 12406
rect 15384 12378 15436 12384
rect 15672 12306 15700 13330
rect 16132 12434 16160 14758
rect 16592 13326 16620 18226
rect 16684 18154 16712 19314
rect 16868 18970 16896 29718
rect 18236 25696 18288 25702
rect 18236 25638 18288 25644
rect 17960 25356 18012 25362
rect 17960 25298 18012 25304
rect 17972 24818 18000 25298
rect 18248 24886 18276 25638
rect 18236 24880 18288 24886
rect 18236 24822 18288 24828
rect 17960 24812 18012 24818
rect 17960 24754 18012 24760
rect 17972 23118 18000 24754
rect 17960 23112 18012 23118
rect 17960 23054 18012 23060
rect 17972 22710 18000 23054
rect 17960 22704 18012 22710
rect 17960 22646 18012 22652
rect 18340 22642 18368 32166
rect 18604 31884 18656 31890
rect 18604 31826 18656 31832
rect 18420 31816 18472 31822
rect 18420 31758 18472 31764
rect 18432 31482 18460 31758
rect 18420 31476 18472 31482
rect 18420 31418 18472 31424
rect 18512 31136 18564 31142
rect 18512 31078 18564 31084
rect 18420 30864 18472 30870
rect 18420 30806 18472 30812
rect 18432 30326 18460 30806
rect 18524 30734 18552 31078
rect 18616 30938 18644 31826
rect 19260 31822 19288 32710
rect 19432 32020 19484 32026
rect 19432 31962 19484 31968
rect 19248 31816 19300 31822
rect 19248 31758 19300 31764
rect 19444 31278 19472 31962
rect 20640 31890 20668 32846
rect 22020 32774 22048 33458
rect 22008 32768 22060 32774
rect 22008 32710 22060 32716
rect 22112 32026 22140 34478
rect 22192 33856 22244 33862
rect 22192 33798 22244 33804
rect 22204 33522 22232 33798
rect 22284 33584 22336 33590
rect 22284 33526 22336 33532
rect 22192 33516 22244 33522
rect 22192 33458 22244 33464
rect 22296 32978 22324 33526
rect 22284 32972 22336 32978
rect 22284 32914 22336 32920
rect 22100 32020 22152 32026
rect 22100 31962 22152 31968
rect 20628 31884 20680 31890
rect 20628 31826 20680 31832
rect 20536 31748 20588 31754
rect 20536 31690 20588 31696
rect 19708 31680 19760 31686
rect 19708 31622 19760 31628
rect 19720 31521 19748 31622
rect 19706 31512 19762 31521
rect 19706 31447 19762 31456
rect 20548 31278 20576 31690
rect 21456 31680 21508 31686
rect 21456 31622 21508 31628
rect 21468 31346 21496 31622
rect 21456 31340 21508 31346
rect 21456 31282 21508 31288
rect 22008 31340 22060 31346
rect 22008 31282 22060 31288
rect 19432 31272 19484 31278
rect 19432 31214 19484 31220
rect 19800 31272 19852 31278
rect 19800 31214 19852 31220
rect 20536 31272 20588 31278
rect 20536 31214 20588 31220
rect 19432 31136 19484 31142
rect 19432 31078 19484 31084
rect 18604 30932 18656 30938
rect 18604 30874 18656 30880
rect 19444 30734 19472 31078
rect 18512 30728 18564 30734
rect 18512 30670 18564 30676
rect 19432 30728 19484 30734
rect 19432 30670 19484 30676
rect 18696 30592 18748 30598
rect 18696 30534 18748 30540
rect 18420 30320 18472 30326
rect 18420 30262 18472 30268
rect 18708 30190 18736 30534
rect 19812 30394 19840 31214
rect 21640 31204 21692 31210
rect 21824 31204 21876 31210
rect 21692 31164 21824 31192
rect 21640 31146 21692 31152
rect 21824 31146 21876 31152
rect 21916 31136 21968 31142
rect 21916 31078 21968 31084
rect 21928 30870 21956 31078
rect 22020 30938 22048 31282
rect 22008 30932 22060 30938
rect 22008 30874 22060 30880
rect 21916 30864 21968 30870
rect 21916 30806 21968 30812
rect 19800 30388 19852 30394
rect 19800 30330 19852 30336
rect 22112 30258 22140 31962
rect 22296 31754 22324 32914
rect 22284 31748 22336 31754
rect 22284 31690 22336 31696
rect 22376 31748 22428 31754
rect 22376 31690 22428 31696
rect 22388 31482 22416 31690
rect 22376 31476 22428 31482
rect 22376 31418 22428 31424
rect 22284 31408 22336 31414
rect 22204 31368 22284 31396
rect 22204 31210 22232 31368
rect 22284 31350 22336 31356
rect 22192 31204 22244 31210
rect 22192 31146 22244 31152
rect 22204 30734 22232 31146
rect 22192 30728 22244 30734
rect 22192 30670 22244 30676
rect 22480 30326 22508 35022
rect 22664 34610 22692 35022
rect 22652 34604 22704 34610
rect 22652 34546 22704 34552
rect 22560 33924 22612 33930
rect 22560 33866 22612 33872
rect 22572 33454 22600 33866
rect 22560 33448 22612 33454
rect 22560 33390 22612 33396
rect 22572 33114 22600 33390
rect 22560 33108 22612 33114
rect 22560 33050 22612 33056
rect 22560 31680 22612 31686
rect 22560 31622 22612 31628
rect 22572 31414 22600 31622
rect 22560 31408 22612 31414
rect 22560 31350 22612 31356
rect 22468 30320 22520 30326
rect 22468 30262 22520 30268
rect 22100 30252 22152 30258
rect 22100 30194 22152 30200
rect 18696 30184 18748 30190
rect 18696 30126 18748 30132
rect 22284 26036 22336 26042
rect 22284 25978 22336 25984
rect 20168 25968 20220 25974
rect 20168 25910 20220 25916
rect 19616 25900 19668 25906
rect 19616 25842 19668 25848
rect 19524 25288 19576 25294
rect 19524 25230 19576 25236
rect 19432 25220 19484 25226
rect 19432 25162 19484 25168
rect 19444 25129 19472 25162
rect 19430 25120 19486 25129
rect 19430 25055 19486 25064
rect 18512 24064 18564 24070
rect 18512 24006 18564 24012
rect 18524 23798 18552 24006
rect 18512 23792 18564 23798
rect 18512 23734 18564 23740
rect 19444 23712 19472 25055
rect 19536 24290 19564 25230
rect 19628 25226 19656 25842
rect 19800 25832 19852 25838
rect 19800 25774 19852 25780
rect 19616 25220 19668 25226
rect 19616 25162 19668 25168
rect 19708 25220 19760 25226
rect 19708 25162 19760 25168
rect 19628 24682 19656 25162
rect 19720 24886 19748 25162
rect 19812 24954 19840 25774
rect 20180 25294 20208 25910
rect 20536 25832 20588 25838
rect 20536 25774 20588 25780
rect 20548 25294 20576 25774
rect 21180 25696 21232 25702
rect 21180 25638 21232 25644
rect 22008 25696 22060 25702
rect 22008 25638 22060 25644
rect 21192 25294 21220 25638
rect 21548 25492 21600 25498
rect 21548 25434 21600 25440
rect 20168 25288 20220 25294
rect 20536 25288 20588 25294
rect 20220 25248 20300 25276
rect 20168 25230 20220 25236
rect 19800 24948 19852 24954
rect 19800 24890 19852 24896
rect 19708 24880 19760 24886
rect 19708 24822 19760 24828
rect 19892 24880 19944 24886
rect 19892 24822 19944 24828
rect 19616 24676 19668 24682
rect 19616 24618 19668 24624
rect 19536 24262 19840 24290
rect 19524 24200 19576 24206
rect 19524 24142 19576 24148
rect 19536 23866 19564 24142
rect 19524 23860 19576 23866
rect 19524 23802 19576 23808
rect 19812 23730 19840 24262
rect 19524 23724 19576 23730
rect 19444 23684 19524 23712
rect 19524 23666 19576 23672
rect 19800 23724 19852 23730
rect 19800 23666 19852 23672
rect 19248 23656 19300 23662
rect 19248 23598 19300 23604
rect 19260 23526 19288 23598
rect 19248 23520 19300 23526
rect 19248 23462 19300 23468
rect 19260 23186 19288 23462
rect 19248 23180 19300 23186
rect 19248 23122 19300 23128
rect 18604 23044 18656 23050
rect 19536 23032 19564 23666
rect 19616 23044 19668 23050
rect 19536 23004 19616 23032
rect 18604 22986 18656 22992
rect 19668 23004 19748 23032
rect 19616 22986 19668 22992
rect 18328 22636 18380 22642
rect 18328 22578 18380 22584
rect 18340 22094 18368 22578
rect 18616 22234 18644 22986
rect 19248 22704 19300 22710
rect 19248 22646 19300 22652
rect 18604 22228 18656 22234
rect 18604 22170 18656 22176
rect 18156 22066 18368 22094
rect 18156 19310 18184 22066
rect 18788 21344 18840 21350
rect 18788 21286 18840 21292
rect 18972 21344 19024 21350
rect 18972 21286 19024 21292
rect 18800 20398 18828 21286
rect 18984 21078 19012 21286
rect 18972 21072 19024 21078
rect 18972 21014 19024 21020
rect 19260 21010 19288 22646
rect 19616 22432 19668 22438
rect 19616 22374 19668 22380
rect 19628 22098 19656 22374
rect 19616 22092 19668 22098
rect 19616 22034 19668 22040
rect 19340 21956 19392 21962
rect 19340 21898 19392 21904
rect 19352 21350 19380 21898
rect 19432 21888 19484 21894
rect 19432 21830 19484 21836
rect 19444 21486 19472 21830
rect 19720 21672 19748 23004
rect 19812 22642 19840 23666
rect 19904 23338 19932 24822
rect 20076 24812 20128 24818
rect 19996 24772 20076 24800
rect 19996 24206 20024 24772
rect 20076 24754 20128 24760
rect 19984 24200 20036 24206
rect 19984 24142 20036 24148
rect 19996 23526 20024 24142
rect 20272 24070 20300 25248
rect 20536 25230 20588 25236
rect 20904 25288 20956 25294
rect 20904 25230 20956 25236
rect 21180 25288 21232 25294
rect 21180 25230 21232 25236
rect 20548 24818 20576 25230
rect 20916 24954 20944 25230
rect 20904 24948 20956 24954
rect 20904 24890 20956 24896
rect 20536 24812 20588 24818
rect 20536 24754 20588 24760
rect 20628 24676 20680 24682
rect 20628 24618 20680 24624
rect 20812 24676 20864 24682
rect 20812 24618 20864 24624
rect 20444 24608 20496 24614
rect 20444 24550 20496 24556
rect 20456 24410 20484 24550
rect 20444 24404 20496 24410
rect 20444 24346 20496 24352
rect 20260 24064 20312 24070
rect 20260 24006 20312 24012
rect 19984 23520 20036 23526
rect 20036 23480 20116 23508
rect 19984 23462 20036 23468
rect 19904 23310 20024 23338
rect 19892 22976 19944 22982
rect 19892 22918 19944 22924
rect 19904 22642 19932 22918
rect 19996 22642 20024 23310
rect 20088 22642 20116 23480
rect 19800 22636 19852 22642
rect 19800 22578 19852 22584
rect 19892 22636 19944 22642
rect 19892 22578 19944 22584
rect 19984 22636 20036 22642
rect 19984 22578 20036 22584
rect 20076 22636 20128 22642
rect 20076 22578 20128 22584
rect 19892 22024 19944 22030
rect 19890 21992 19892 22001
rect 19944 21992 19946 22001
rect 19890 21927 19946 21936
rect 19720 21644 19840 21672
rect 19708 21548 19760 21554
rect 19536 21508 19708 21536
rect 19432 21480 19484 21486
rect 19432 21422 19484 21428
rect 19340 21344 19392 21350
rect 19340 21286 19392 21292
rect 19248 21004 19300 21010
rect 19168 20964 19248 20992
rect 19168 20602 19196 20964
rect 19248 20946 19300 20952
rect 19156 20596 19208 20602
rect 19156 20538 19208 20544
rect 18788 20392 18840 20398
rect 18788 20334 18840 20340
rect 19536 20262 19564 21508
rect 19708 21490 19760 21496
rect 19812 20874 19840 21644
rect 19800 20868 19852 20874
rect 19800 20810 19852 20816
rect 19812 20618 19840 20810
rect 19807 20590 19840 20618
rect 19807 20505 19835 20590
rect 19798 20496 19854 20505
rect 19798 20431 19800 20440
rect 19852 20431 19854 20440
rect 19800 20402 19852 20408
rect 19524 20256 19576 20262
rect 19524 20198 19576 20204
rect 19340 19508 19392 19514
rect 19340 19450 19392 19456
rect 18144 19304 18196 19310
rect 18144 19246 18196 19252
rect 17592 19168 17644 19174
rect 17592 19110 17644 19116
rect 16856 18964 16908 18970
rect 16856 18906 16908 18912
rect 17604 18834 17632 19110
rect 17592 18828 17644 18834
rect 17592 18770 17644 18776
rect 16764 18760 16816 18766
rect 16764 18702 16816 18708
rect 17316 18760 17368 18766
rect 17316 18702 17368 18708
rect 16672 18148 16724 18154
rect 16672 18090 16724 18096
rect 16684 17678 16712 18090
rect 16672 17672 16724 17678
rect 16672 17614 16724 17620
rect 16684 17134 16712 17614
rect 16776 17338 16804 18702
rect 17328 18222 17356 18702
rect 17960 18624 18012 18630
rect 17960 18566 18012 18572
rect 17316 18216 17368 18222
rect 17316 18158 17368 18164
rect 16764 17332 16816 17338
rect 16764 17274 16816 17280
rect 17972 17270 18000 18566
rect 18156 18290 18184 19246
rect 19352 19242 19380 19450
rect 19536 19378 19564 20198
rect 19904 19530 19932 21927
rect 19996 21690 20024 22578
rect 20352 22568 20404 22574
rect 20456 22545 20484 24346
rect 20640 23730 20668 24618
rect 20824 23798 20852 24618
rect 21560 24274 21588 25434
rect 21824 25356 21876 25362
rect 21824 25298 21876 25304
rect 21730 25256 21786 25265
rect 21730 25191 21786 25200
rect 21744 24750 21772 25191
rect 21836 24750 21864 25298
rect 22020 25226 22048 25638
rect 22192 25492 22244 25498
rect 22192 25434 22244 25440
rect 22008 25220 22060 25226
rect 22008 25162 22060 25168
rect 21732 24744 21784 24750
rect 21732 24686 21784 24692
rect 21824 24744 21876 24750
rect 21824 24686 21876 24692
rect 22204 24596 22232 25434
rect 22112 24568 22232 24596
rect 21824 24336 21876 24342
rect 21824 24278 21876 24284
rect 21548 24268 21600 24274
rect 21548 24210 21600 24216
rect 20994 23896 21050 23905
rect 20994 23831 20996 23840
rect 21048 23831 21050 23840
rect 20996 23802 21048 23808
rect 20812 23792 20864 23798
rect 20812 23734 20864 23740
rect 20628 23724 20680 23730
rect 20628 23666 20680 23672
rect 21008 23322 21036 23802
rect 20996 23316 21048 23322
rect 20996 23258 21048 23264
rect 20352 22510 20404 22516
rect 20442 22536 20498 22545
rect 20074 22400 20130 22409
rect 20074 22335 20130 22344
rect 20088 21894 20116 22335
rect 20364 21978 20392 22510
rect 20442 22471 20498 22480
rect 20444 22432 20496 22438
rect 20444 22374 20496 22380
rect 20456 22234 20484 22374
rect 20444 22228 20496 22234
rect 20444 22170 20496 22176
rect 21008 22098 21036 23258
rect 21560 23186 21588 24210
rect 21836 24070 21864 24278
rect 22112 24138 22140 24568
rect 22296 24206 22324 25978
rect 22376 25900 22428 25906
rect 22376 25842 22428 25848
rect 22388 25498 22416 25842
rect 22376 25492 22428 25498
rect 22376 25434 22428 25440
rect 22376 25152 22428 25158
rect 22376 25094 22428 25100
rect 22388 24886 22416 25094
rect 22376 24880 22428 24886
rect 22480 24868 22508 30262
rect 22560 24880 22612 24886
rect 22480 24840 22560 24868
rect 22376 24822 22428 24828
rect 22560 24822 22612 24828
rect 22572 24410 22600 24822
rect 22560 24404 22612 24410
rect 22560 24346 22612 24352
rect 22374 24304 22430 24313
rect 22374 24239 22430 24248
rect 22560 24268 22612 24274
rect 22284 24200 22336 24206
rect 22284 24142 22336 24148
rect 22100 24132 22152 24138
rect 22100 24074 22152 24080
rect 21824 24064 21876 24070
rect 22112 24041 22140 24074
rect 22192 24064 22244 24070
rect 21824 24006 21876 24012
rect 22098 24032 22154 24041
rect 21548 23180 21600 23186
rect 21548 23122 21600 23128
rect 20996 22092 21048 22098
rect 20996 22034 21048 22040
rect 20272 21950 20392 21978
rect 20536 21956 20588 21962
rect 20076 21888 20128 21894
rect 20076 21830 20128 21836
rect 19984 21684 20036 21690
rect 19984 21626 20036 21632
rect 20168 21684 20220 21690
rect 20168 21626 20220 21632
rect 19984 21548 20036 21554
rect 19984 21490 20036 21496
rect 19996 21010 20024 21490
rect 20180 21146 20208 21626
rect 20272 21554 20300 21950
rect 20536 21898 20588 21904
rect 20904 21956 20956 21962
rect 20904 21898 20956 21904
rect 20352 21888 20404 21894
rect 20352 21830 20404 21836
rect 20260 21548 20312 21554
rect 20260 21490 20312 21496
rect 20272 21418 20300 21490
rect 20260 21412 20312 21418
rect 20260 21354 20312 21360
rect 20168 21140 20220 21146
rect 20168 21082 20220 21088
rect 19984 21004 20036 21010
rect 19984 20946 20036 20952
rect 19996 20777 20024 20946
rect 19982 20768 20038 20777
rect 19982 20703 20038 20712
rect 20364 20534 20392 21830
rect 20442 21720 20498 21729
rect 20442 21655 20444 21664
rect 20496 21655 20498 21664
rect 20444 21626 20496 21632
rect 20444 21548 20496 21554
rect 20548 21536 20576 21898
rect 20916 21690 20944 21898
rect 21560 21894 21588 23122
rect 21836 23118 21864 24006
rect 22192 24006 22244 24012
rect 22098 23967 22154 23976
rect 22100 23792 22152 23798
rect 22100 23734 22152 23740
rect 22008 23724 22060 23730
rect 22008 23666 22060 23672
rect 21824 23112 21876 23118
rect 21824 23054 21876 23060
rect 21836 22438 21864 23054
rect 22020 22778 22048 23666
rect 22112 23186 22140 23734
rect 22204 23322 22232 24006
rect 22296 23662 22324 24142
rect 22284 23656 22336 23662
rect 22284 23598 22336 23604
rect 22192 23316 22244 23322
rect 22192 23258 22244 23264
rect 22388 23186 22416 24239
rect 22560 24210 22612 24216
rect 22468 24200 22520 24206
rect 22468 24142 22520 24148
rect 22480 23322 22508 24142
rect 22572 23905 22600 24210
rect 22558 23896 22614 23905
rect 22558 23831 22614 23840
rect 22468 23316 22520 23322
rect 22468 23258 22520 23264
rect 22100 23180 22152 23186
rect 22100 23122 22152 23128
rect 22376 23180 22428 23186
rect 22376 23122 22428 23128
rect 22008 22772 22060 22778
rect 22008 22714 22060 22720
rect 22112 22710 22140 23122
rect 22192 22976 22244 22982
rect 22192 22918 22244 22924
rect 22100 22704 22152 22710
rect 22100 22646 22152 22652
rect 21824 22432 21876 22438
rect 21824 22374 21876 22380
rect 21548 21888 21600 21894
rect 21548 21830 21600 21836
rect 20904 21684 20956 21690
rect 20904 21626 20956 21632
rect 20496 21508 20576 21536
rect 20444 21490 20496 21496
rect 20456 20618 20484 21490
rect 21560 21350 21588 21830
rect 21548 21344 21600 21350
rect 21548 21286 21600 21292
rect 21836 20942 21864 22374
rect 22112 21078 22140 22646
rect 22204 22574 22232 22918
rect 22560 22704 22612 22710
rect 22560 22646 22612 22652
rect 22192 22568 22244 22574
rect 22192 22510 22244 22516
rect 22284 21888 22336 21894
rect 22284 21830 22336 21836
rect 22100 21072 22152 21078
rect 22100 21014 22152 21020
rect 21824 20936 21876 20942
rect 21824 20878 21876 20884
rect 20996 20800 21048 20806
rect 20994 20768 20996 20777
rect 21048 20768 21050 20777
rect 20994 20703 21050 20712
rect 20456 20602 20576 20618
rect 20456 20596 20588 20602
rect 20456 20590 20536 20596
rect 20352 20528 20404 20534
rect 20352 20470 20404 20476
rect 20456 20398 20484 20590
rect 20536 20538 20588 20544
rect 22112 20534 22140 21014
rect 22296 21010 22324 21830
rect 22376 21548 22428 21554
rect 22376 21490 22428 21496
rect 22284 21004 22336 21010
rect 22284 20946 22336 20952
rect 22388 20942 22416 21490
rect 22376 20936 22428 20942
rect 22376 20878 22428 20884
rect 22192 20800 22244 20806
rect 22192 20742 22244 20748
rect 22100 20528 22152 20534
rect 22100 20470 22152 20476
rect 22204 20398 22232 20742
rect 22572 20534 22600 22646
rect 22560 20528 22612 20534
rect 22558 20496 22560 20505
rect 22612 20496 22614 20505
rect 22558 20431 22614 20440
rect 20444 20392 20496 20398
rect 20444 20334 20496 20340
rect 22192 20392 22244 20398
rect 22192 20334 22244 20340
rect 19904 19502 20024 19530
rect 19892 19440 19944 19446
rect 19892 19382 19944 19388
rect 19524 19372 19576 19378
rect 19524 19314 19576 19320
rect 19616 19372 19668 19378
rect 19616 19314 19668 19320
rect 19800 19372 19852 19378
rect 19800 19314 19852 19320
rect 19340 19236 19392 19242
rect 19340 19178 19392 19184
rect 19248 19168 19300 19174
rect 19248 19110 19300 19116
rect 18144 18284 18196 18290
rect 18144 18226 18196 18232
rect 17960 17264 18012 17270
rect 17960 17206 18012 17212
rect 16672 17128 16724 17134
rect 16672 17070 16724 17076
rect 16684 16658 16712 17070
rect 16672 16652 16724 16658
rect 16672 16594 16724 16600
rect 16684 15162 16712 16594
rect 17972 16522 18000 17206
rect 19260 16998 19288 19110
rect 19536 18834 19564 19314
rect 19628 18902 19656 19314
rect 19616 18896 19668 18902
rect 19616 18838 19668 18844
rect 19524 18828 19576 18834
rect 19524 18770 19576 18776
rect 19812 18737 19840 19314
rect 19798 18728 19854 18737
rect 19524 18692 19576 18698
rect 19798 18663 19854 18672
rect 19524 18634 19576 18640
rect 19340 17128 19392 17134
rect 19340 17070 19392 17076
rect 19248 16992 19300 16998
rect 19248 16934 19300 16940
rect 18880 16584 18932 16590
rect 18880 16526 18932 16532
rect 18972 16584 19024 16590
rect 18972 16526 19024 16532
rect 17960 16516 18012 16522
rect 17960 16458 18012 16464
rect 16672 15156 16724 15162
rect 16672 15098 16724 15104
rect 17868 14952 17920 14958
rect 17868 14894 17920 14900
rect 17880 14482 17908 14894
rect 17316 14476 17368 14482
rect 17316 14418 17368 14424
rect 17868 14476 17920 14482
rect 17868 14418 17920 14424
rect 16764 14272 16816 14278
rect 16764 14214 16816 14220
rect 16776 13870 16804 14214
rect 16764 13864 16816 13870
rect 16764 13806 16816 13812
rect 16672 13388 16724 13394
rect 16672 13330 16724 13336
rect 16580 13320 16632 13326
rect 16580 13262 16632 13268
rect 16592 12986 16620 13262
rect 16580 12980 16632 12986
rect 16580 12922 16632 12928
rect 16684 12782 16712 13330
rect 16672 12776 16724 12782
rect 16672 12718 16724 12724
rect 16040 12406 16160 12434
rect 14740 12300 14792 12306
rect 14740 12242 14792 12248
rect 15660 12300 15712 12306
rect 15660 12242 15712 12248
rect 13452 12164 13504 12170
rect 13452 12106 13504 12112
rect 13464 11830 13492 12106
rect 14096 12096 14148 12102
rect 14096 12038 14148 12044
rect 13452 11824 13504 11830
rect 13452 11766 13504 11772
rect 12164 11756 12216 11762
rect 12164 11698 12216 11704
rect 12440 11688 12492 11694
rect 12440 11630 12492 11636
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 12452 11354 12480 11630
rect 14004 11552 14056 11558
rect 14004 11494 14056 11500
rect 12440 11348 12492 11354
rect 12440 11290 12492 11296
rect 13544 11212 13596 11218
rect 13544 11154 13596 11160
rect 4874 10908 5182 10917
rect 4874 10906 4880 10908
rect 4936 10906 4960 10908
rect 5016 10906 5040 10908
rect 5096 10906 5120 10908
rect 5176 10906 5182 10908
rect 4936 10854 4938 10906
rect 5118 10854 5120 10906
rect 4874 10852 4880 10854
rect 4936 10852 4960 10854
rect 5016 10852 5040 10854
rect 5096 10852 5120 10854
rect 5176 10852 5182 10854
rect 4874 10843 5182 10852
rect 13556 10810 13584 11154
rect 14016 11150 14044 11494
rect 14108 11150 14136 12038
rect 14752 11762 14780 12242
rect 14832 12232 14884 12238
rect 14832 12174 14884 12180
rect 15292 12232 15344 12238
rect 15292 12174 15344 12180
rect 14740 11756 14792 11762
rect 14740 11698 14792 11704
rect 14280 11688 14332 11694
rect 14280 11630 14332 11636
rect 14292 11150 14320 11630
rect 14752 11218 14780 11698
rect 14844 11354 14872 12174
rect 15304 12102 15332 12174
rect 15292 12096 15344 12102
rect 15292 12038 15344 12044
rect 14832 11348 14884 11354
rect 14832 11290 14884 11296
rect 15304 11286 15332 12038
rect 15476 11552 15528 11558
rect 15476 11494 15528 11500
rect 15292 11280 15344 11286
rect 15292 11222 15344 11228
rect 14740 11212 14792 11218
rect 14740 11154 14792 11160
rect 15488 11150 15516 11494
rect 15660 11348 15712 11354
rect 15660 11290 15712 11296
rect 14004 11144 14056 11150
rect 14004 11086 14056 11092
rect 14096 11144 14148 11150
rect 14096 11086 14148 11092
rect 14280 11144 14332 11150
rect 14280 11086 14332 11092
rect 15476 11144 15528 11150
rect 15476 11086 15528 11092
rect 15672 11014 15700 11290
rect 16040 11150 16068 12406
rect 16396 11552 16448 11558
rect 16396 11494 16448 11500
rect 16408 11354 16436 11494
rect 16684 11354 16712 12718
rect 16776 12238 16804 13806
rect 17328 13394 17356 14418
rect 17972 14346 18000 16458
rect 18892 15706 18920 16526
rect 18984 16454 19012 16526
rect 19352 16522 19380 17070
rect 19536 16658 19564 18634
rect 19616 18624 19668 18630
rect 19616 18566 19668 18572
rect 19708 18624 19760 18630
rect 19708 18566 19760 18572
rect 19628 18290 19656 18566
rect 19616 18284 19668 18290
rect 19616 18226 19668 18232
rect 19720 17218 19748 18566
rect 19628 17190 19748 17218
rect 19812 17202 19840 18663
rect 19904 18426 19932 19382
rect 19892 18420 19944 18426
rect 19892 18362 19944 18368
rect 19800 17196 19852 17202
rect 19524 16652 19576 16658
rect 19524 16594 19576 16600
rect 19340 16516 19392 16522
rect 19340 16458 19392 16464
rect 18972 16448 19024 16454
rect 18972 16390 19024 16396
rect 18984 16046 19012 16390
rect 19536 16250 19564 16594
rect 19628 16522 19656 17190
rect 19800 17138 19852 17144
rect 19708 17128 19760 17134
rect 19708 17070 19760 17076
rect 19720 16590 19748 17070
rect 19996 16640 20024 19502
rect 20076 19508 20128 19514
rect 20076 19450 20128 19456
rect 20088 19242 20116 19450
rect 20456 19446 20484 20334
rect 22664 19990 22692 34546
rect 23112 34536 23164 34542
rect 23112 34478 23164 34484
rect 23388 34536 23440 34542
rect 23388 34478 23440 34484
rect 23124 33998 23152 34478
rect 23112 33992 23164 33998
rect 23112 33934 23164 33940
rect 23400 33658 23428 34478
rect 23388 33652 23440 33658
rect 23388 33594 23440 33600
rect 23572 33312 23624 33318
rect 23572 33254 23624 33260
rect 23584 33046 23612 33254
rect 23768 33114 23796 35634
rect 25044 35624 25096 35630
rect 25044 35566 25096 35572
rect 24860 35080 24912 35086
rect 24860 35022 24912 35028
rect 24872 34746 24900 35022
rect 25056 34746 25084 35566
rect 25136 35488 25188 35494
rect 25136 35430 25188 35436
rect 24860 34740 24912 34746
rect 24860 34682 24912 34688
rect 25044 34740 25096 34746
rect 25044 34682 25096 34688
rect 24952 34400 25004 34406
rect 24952 34342 25004 34348
rect 24964 33590 24992 34342
rect 25056 33930 25084 34682
rect 25044 33924 25096 33930
rect 25044 33866 25096 33872
rect 24952 33584 25004 33590
rect 24952 33526 25004 33532
rect 25056 33522 25084 33866
rect 24860 33516 24912 33522
rect 24860 33458 24912 33464
rect 25044 33516 25096 33522
rect 25044 33458 25096 33464
rect 23756 33108 23808 33114
rect 23756 33050 23808 33056
rect 23572 33040 23624 33046
rect 23572 32982 23624 32988
rect 23584 32910 23612 32982
rect 23572 32904 23624 32910
rect 23572 32846 23624 32852
rect 23664 31884 23716 31890
rect 23664 31826 23716 31832
rect 23386 31512 23442 31521
rect 23386 31447 23442 31456
rect 23400 31414 23428 31447
rect 23388 31408 23440 31414
rect 23388 31350 23440 31356
rect 23676 31142 23704 31826
rect 23768 31754 23796 33050
rect 24872 32910 24900 33458
rect 23848 32904 23900 32910
rect 23848 32846 23900 32852
rect 24860 32904 24912 32910
rect 24860 32846 24912 32852
rect 23756 31748 23808 31754
rect 23756 31690 23808 31696
rect 23860 31482 23888 32846
rect 24584 32768 24636 32774
rect 24584 32710 24636 32716
rect 24596 32026 24624 32710
rect 24584 32020 24636 32026
rect 24584 31962 24636 31968
rect 24400 31680 24452 31686
rect 24400 31622 24452 31628
rect 23848 31476 23900 31482
rect 23848 31418 23900 31424
rect 22928 31136 22980 31142
rect 22928 31078 22980 31084
rect 23664 31136 23716 31142
rect 23664 31078 23716 31084
rect 22744 30864 22796 30870
rect 22744 30806 22796 30812
rect 22756 30598 22784 30806
rect 22940 30734 22968 31078
rect 24412 30734 24440 31622
rect 24860 31476 24912 31482
rect 24860 31418 24912 31424
rect 24676 31340 24728 31346
rect 24676 31282 24728 31288
rect 22928 30728 22980 30734
rect 22928 30670 22980 30676
rect 24400 30728 24452 30734
rect 24400 30670 24452 30676
rect 24688 30598 24716 31282
rect 24872 30666 24900 31418
rect 25044 30932 25096 30938
rect 25044 30874 25096 30880
rect 24860 30660 24912 30666
rect 24860 30602 24912 30608
rect 22744 30592 22796 30598
rect 22744 30534 22796 30540
rect 24676 30592 24728 30598
rect 24676 30534 24728 30540
rect 22756 29714 22784 30534
rect 24872 30394 24900 30602
rect 25056 30394 25084 30874
rect 24860 30388 24912 30394
rect 24860 30330 24912 30336
rect 25044 30388 25096 30394
rect 25044 30330 25096 30336
rect 22836 30184 22888 30190
rect 22836 30126 22888 30132
rect 22848 29850 22876 30126
rect 22836 29844 22888 29850
rect 22836 29786 22888 29792
rect 24872 29714 24900 30330
rect 22744 29708 22796 29714
rect 22744 29650 22796 29656
rect 24860 29708 24912 29714
rect 24860 29650 24912 29656
rect 22836 26920 22888 26926
rect 22836 26862 22888 26868
rect 23480 26920 23532 26926
rect 23480 26862 23532 26868
rect 22744 26240 22796 26246
rect 22744 26182 22796 26188
rect 22756 26042 22784 26182
rect 22744 26036 22796 26042
rect 22744 25978 22796 25984
rect 22756 25906 22784 25978
rect 22744 25900 22796 25906
rect 22744 25842 22796 25848
rect 22756 22234 22784 25842
rect 22848 24750 22876 26862
rect 23492 26586 23520 26862
rect 24952 26784 25004 26790
rect 24952 26726 25004 26732
rect 23480 26580 23532 26586
rect 23480 26522 23532 26528
rect 24964 26382 24992 26726
rect 24768 26376 24820 26382
rect 24768 26318 24820 26324
rect 24952 26376 25004 26382
rect 24952 26318 25004 26324
rect 25042 26344 25098 26353
rect 23296 25900 23348 25906
rect 23296 25842 23348 25848
rect 23480 25900 23532 25906
rect 23480 25842 23532 25848
rect 24124 25900 24176 25906
rect 24124 25842 24176 25848
rect 23020 25832 23072 25838
rect 23072 25792 23152 25820
rect 23020 25774 23072 25780
rect 23020 25220 23072 25226
rect 23020 25162 23072 25168
rect 23032 25129 23060 25162
rect 23018 25120 23074 25129
rect 23018 25055 23074 25064
rect 22836 24744 22888 24750
rect 22836 24686 22888 24692
rect 22848 24585 22876 24686
rect 23124 24682 23152 25792
rect 23308 25498 23336 25842
rect 23388 25832 23440 25838
rect 23388 25774 23440 25780
rect 23296 25492 23348 25498
rect 23296 25434 23348 25440
rect 23400 25362 23428 25774
rect 23388 25356 23440 25362
rect 23388 25298 23440 25304
rect 23492 25294 23520 25842
rect 23296 25288 23348 25294
rect 23294 25256 23296 25265
rect 23480 25288 23532 25294
rect 23348 25256 23350 25265
rect 23480 25230 23532 25236
rect 23294 25191 23350 25200
rect 23572 25220 23624 25226
rect 23572 25162 23624 25168
rect 23296 25152 23348 25158
rect 23296 25094 23348 25100
rect 23112 24676 23164 24682
rect 23112 24618 23164 24624
rect 23308 24614 23336 25094
rect 23584 24954 23612 25162
rect 23572 24948 23624 24954
rect 23572 24890 23624 24896
rect 23584 24614 23612 24890
rect 23296 24608 23348 24614
rect 22834 24576 22890 24585
rect 23296 24550 23348 24556
rect 23572 24608 23624 24614
rect 23572 24550 23624 24556
rect 22834 24511 22890 24520
rect 22848 23798 22876 24511
rect 22928 24404 22980 24410
rect 22928 24346 22980 24352
rect 23112 24404 23164 24410
rect 23112 24346 23164 24352
rect 22940 24313 22968 24346
rect 22926 24304 22982 24313
rect 22926 24239 22982 24248
rect 22928 24132 22980 24138
rect 22928 24074 22980 24080
rect 22940 23866 22968 24074
rect 23124 23866 23152 24346
rect 23296 24336 23348 24342
rect 23296 24278 23348 24284
rect 22928 23860 22980 23866
rect 22928 23802 22980 23808
rect 23112 23860 23164 23866
rect 23112 23802 23164 23808
rect 22836 23792 22888 23798
rect 22836 23734 22888 23740
rect 22836 23044 22888 23050
rect 22836 22986 22888 22992
rect 22848 22778 22876 22986
rect 22836 22772 22888 22778
rect 22836 22714 22888 22720
rect 22744 22228 22796 22234
rect 22744 22170 22796 22176
rect 23308 21894 23336 24278
rect 23584 24274 23612 24550
rect 23572 24268 23624 24274
rect 23572 24210 23624 24216
rect 23664 24200 23716 24206
rect 23664 24142 23716 24148
rect 23572 23724 23624 23730
rect 23572 23666 23624 23672
rect 23584 22094 23612 23666
rect 23676 23322 23704 24142
rect 23846 24032 23902 24041
rect 23846 23967 23902 23976
rect 23860 23730 23888 23967
rect 23756 23724 23808 23730
rect 23756 23666 23808 23672
rect 23848 23724 23900 23730
rect 23848 23666 23900 23672
rect 24032 23724 24084 23730
rect 24032 23666 24084 23672
rect 23664 23316 23716 23322
rect 23664 23258 23716 23264
rect 23664 22976 23716 22982
rect 23664 22918 23716 22924
rect 23676 22778 23704 22918
rect 23664 22772 23716 22778
rect 23664 22714 23716 22720
rect 23768 22642 23796 23666
rect 23756 22636 23808 22642
rect 23756 22578 23808 22584
rect 23584 22066 23704 22094
rect 23296 21888 23348 21894
rect 23296 21830 23348 21836
rect 23572 21684 23624 21690
rect 23572 21626 23624 21632
rect 23204 20868 23256 20874
rect 23204 20810 23256 20816
rect 23216 20505 23244 20810
rect 23202 20496 23258 20505
rect 23202 20431 23258 20440
rect 23584 20398 23612 21626
rect 23676 21486 23704 22066
rect 23860 21729 23888 23666
rect 24044 22982 24072 23666
rect 24032 22976 24084 22982
rect 24032 22918 24084 22924
rect 24032 21888 24084 21894
rect 24032 21830 24084 21836
rect 23846 21720 23902 21729
rect 23846 21655 23902 21664
rect 23860 21554 23888 21655
rect 23848 21548 23900 21554
rect 23848 21490 23900 21496
rect 23664 21480 23716 21486
rect 23716 21428 23980 21434
rect 23664 21422 23980 21428
rect 23676 21406 23980 21422
rect 23952 21350 23980 21406
rect 23848 21344 23900 21350
rect 23848 21286 23900 21292
rect 23940 21344 23992 21350
rect 23940 21286 23992 21292
rect 23664 20800 23716 20806
rect 23664 20742 23716 20748
rect 23676 20602 23704 20742
rect 23664 20596 23716 20602
rect 23664 20538 23716 20544
rect 23860 20466 23888 21286
rect 24044 20466 24072 21830
rect 24136 21554 24164 25842
rect 24780 25770 24808 26318
rect 24860 26240 24912 26246
rect 24860 26182 24912 26188
rect 24872 25770 24900 26182
rect 24768 25764 24820 25770
rect 24768 25706 24820 25712
rect 24860 25764 24912 25770
rect 24860 25706 24912 25712
rect 24964 25362 24992 26318
rect 25042 26279 25098 26288
rect 25056 25906 25084 26279
rect 25044 25900 25096 25906
rect 25044 25842 25096 25848
rect 25044 25424 25096 25430
rect 25044 25366 25096 25372
rect 24952 25356 25004 25362
rect 24952 25298 25004 25304
rect 24216 25152 24268 25158
rect 24216 25094 24268 25100
rect 24228 21962 24256 25094
rect 25056 24290 25084 25366
rect 25148 24410 25176 35430
rect 25240 33114 25268 35770
rect 26700 35760 26752 35766
rect 26700 35702 26752 35708
rect 29276 35760 29328 35766
rect 29276 35702 29328 35708
rect 25320 35624 25372 35630
rect 25320 35566 25372 35572
rect 25332 35290 25360 35566
rect 25320 35284 25372 35290
rect 25320 35226 25372 35232
rect 25688 35080 25740 35086
rect 25688 35022 25740 35028
rect 25872 35080 25924 35086
rect 25872 35022 25924 35028
rect 26056 35080 26108 35086
rect 26056 35022 26108 35028
rect 26332 35080 26384 35086
rect 26332 35022 26384 35028
rect 25700 34678 25728 35022
rect 25688 34672 25740 34678
rect 25688 34614 25740 34620
rect 25780 34196 25832 34202
rect 25780 34138 25832 34144
rect 25792 33998 25820 34138
rect 25780 33992 25832 33998
rect 25700 33952 25780 33980
rect 25320 33448 25372 33454
rect 25320 33390 25372 33396
rect 25332 33114 25360 33390
rect 25228 33108 25280 33114
rect 25228 33050 25280 33056
rect 25320 33108 25372 33114
rect 25320 33050 25372 33056
rect 25240 30054 25268 33050
rect 25700 33046 25728 33952
rect 25780 33934 25832 33940
rect 25884 33862 25912 35022
rect 26068 34542 26096 35022
rect 26056 34536 26108 34542
rect 26056 34478 26108 34484
rect 26240 34128 26292 34134
rect 26240 34070 26292 34076
rect 25872 33856 25924 33862
rect 25872 33798 25924 33804
rect 25688 33040 25740 33046
rect 25688 32982 25740 32988
rect 25884 32774 25912 33798
rect 25964 33312 26016 33318
rect 25964 33254 26016 33260
rect 25976 32910 26004 33254
rect 26252 32978 26280 34070
rect 26344 33998 26372 35022
rect 26424 35012 26476 35018
rect 26424 34954 26476 34960
rect 26436 34610 26464 34954
rect 26608 34944 26660 34950
rect 26608 34886 26660 34892
rect 26424 34604 26476 34610
rect 26424 34546 26476 34552
rect 26620 34542 26648 34886
rect 26608 34536 26660 34542
rect 26608 34478 26660 34484
rect 26712 34406 26740 35702
rect 28816 35692 28868 35698
rect 28816 35634 28868 35640
rect 27804 35624 27856 35630
rect 27804 35566 27856 35572
rect 26792 35488 26844 35494
rect 26792 35430 26844 35436
rect 26804 35018 26832 35430
rect 27816 35154 27844 35566
rect 28828 35290 28856 35634
rect 28816 35284 28868 35290
rect 28816 35226 28868 35232
rect 27804 35148 27856 35154
rect 27804 35090 27856 35096
rect 28816 35148 28868 35154
rect 28816 35090 28868 35096
rect 26792 35012 26844 35018
rect 26792 34954 26844 34960
rect 26804 34610 26832 34954
rect 27068 34944 27120 34950
rect 27068 34886 27120 34892
rect 27080 34678 27108 34886
rect 27816 34746 27844 35090
rect 27804 34740 27856 34746
rect 27804 34682 27856 34688
rect 27068 34672 27120 34678
rect 27068 34614 27120 34620
rect 26792 34604 26844 34610
rect 26792 34546 26844 34552
rect 26804 34406 26832 34546
rect 26700 34400 26752 34406
rect 26700 34342 26752 34348
rect 26792 34400 26844 34406
rect 26792 34342 26844 34348
rect 27252 34400 27304 34406
rect 27252 34342 27304 34348
rect 26332 33992 26384 33998
rect 26332 33934 26384 33940
rect 26516 33992 26568 33998
rect 26516 33934 26568 33940
rect 26332 33856 26384 33862
rect 26332 33798 26384 33804
rect 26344 33114 26372 33798
rect 26528 33640 26556 33934
rect 26608 33652 26660 33658
rect 26528 33612 26608 33640
rect 26332 33108 26384 33114
rect 26332 33050 26384 33056
rect 26240 32972 26292 32978
rect 26240 32914 26292 32920
rect 25964 32904 26016 32910
rect 25964 32846 26016 32852
rect 25872 32768 25924 32774
rect 25872 32710 25924 32716
rect 26344 32434 26372 33050
rect 26332 32428 26384 32434
rect 26332 32370 26384 32376
rect 26528 32366 26556 33612
rect 26608 33594 26660 33600
rect 26712 33590 26740 34342
rect 27160 33992 27212 33998
rect 27160 33934 27212 33940
rect 26700 33584 26752 33590
rect 26700 33526 26752 33532
rect 26712 32858 26740 33526
rect 27172 33318 27200 33934
rect 27264 33658 27292 34342
rect 27344 33856 27396 33862
rect 27344 33798 27396 33804
rect 27252 33652 27304 33658
rect 27252 33594 27304 33600
rect 27356 33590 27384 33798
rect 27344 33584 27396 33590
rect 27344 33526 27396 33532
rect 27816 33522 27844 34682
rect 28828 34610 28856 35090
rect 29288 35018 29316 35702
rect 29564 35290 29592 35974
rect 29748 35834 29776 36042
rect 29736 35828 29788 35834
rect 29736 35770 29788 35776
rect 31680 35290 31708 37198
rect 32232 36922 32260 39200
rect 32876 36922 32904 39200
rect 33520 36922 33548 39200
rect 34164 36922 34192 39200
rect 34808 36922 34836 39200
rect 34934 37564 35242 37573
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37499 35242 37508
rect 35452 36922 35480 39200
rect 35594 37020 35902 37029
rect 35594 37018 35600 37020
rect 35656 37018 35680 37020
rect 35736 37018 35760 37020
rect 35816 37018 35840 37020
rect 35896 37018 35902 37020
rect 35656 36966 35658 37018
rect 35838 36966 35840 37018
rect 35594 36964 35600 36966
rect 35656 36964 35680 36966
rect 35736 36964 35760 36966
rect 35816 36964 35840 36966
rect 35896 36964 35902 36966
rect 35594 36955 35902 36964
rect 36096 36922 36124 39200
rect 36740 36922 36768 39200
rect 37384 36922 37412 39200
rect 38028 36922 38056 39200
rect 38672 36922 38700 39200
rect 39316 36922 39344 39200
rect 39960 36922 39988 39200
rect 40604 36922 40632 39200
rect 41248 36922 41276 39200
rect 41892 36922 41920 39200
rect 42536 36922 42564 39200
rect 43180 36922 43208 39200
rect 43824 36922 43852 39200
rect 44468 36922 44496 39200
rect 45112 36922 45140 39200
rect 45756 36922 45784 39200
rect 46400 36922 46428 39200
rect 47044 36922 47072 39200
rect 47688 36922 47716 39200
rect 32220 36916 32272 36922
rect 32220 36858 32272 36864
rect 32864 36916 32916 36922
rect 32864 36858 32916 36864
rect 33508 36916 33560 36922
rect 33508 36858 33560 36864
rect 34152 36916 34204 36922
rect 34152 36858 34204 36864
rect 34796 36916 34848 36922
rect 34796 36858 34848 36864
rect 35440 36916 35492 36922
rect 35440 36858 35492 36864
rect 36084 36916 36136 36922
rect 36084 36858 36136 36864
rect 36728 36916 36780 36922
rect 36728 36858 36780 36864
rect 37372 36916 37424 36922
rect 37372 36858 37424 36864
rect 38016 36916 38068 36922
rect 38016 36858 38068 36864
rect 38660 36916 38712 36922
rect 38660 36858 38712 36864
rect 39304 36916 39356 36922
rect 39304 36858 39356 36864
rect 39948 36916 40000 36922
rect 39948 36858 40000 36864
rect 40592 36916 40644 36922
rect 40592 36858 40644 36864
rect 41236 36916 41288 36922
rect 41236 36858 41288 36864
rect 41880 36916 41932 36922
rect 41880 36858 41932 36864
rect 42524 36916 42576 36922
rect 42524 36858 42576 36864
rect 43168 36916 43220 36922
rect 43168 36858 43220 36864
rect 43812 36916 43864 36922
rect 43812 36858 43864 36864
rect 44456 36916 44508 36922
rect 44456 36858 44508 36864
rect 45100 36916 45152 36922
rect 45100 36858 45152 36864
rect 45744 36916 45796 36922
rect 45744 36858 45796 36864
rect 46388 36916 46440 36922
rect 46388 36858 46440 36864
rect 47032 36916 47084 36922
rect 47032 36858 47084 36864
rect 47676 36916 47728 36922
rect 47676 36858 47728 36864
rect 32220 36780 32272 36786
rect 32220 36722 32272 36728
rect 35348 36780 35400 36786
rect 35348 36722 35400 36728
rect 37372 36780 37424 36786
rect 37372 36722 37424 36728
rect 42524 36780 42576 36786
rect 42524 36722 42576 36728
rect 46204 36780 46256 36786
rect 46204 36722 46256 36728
rect 32232 36378 32260 36722
rect 34934 36476 35242 36485
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36411 35242 36420
rect 35360 36378 35388 36722
rect 37384 36378 37412 36722
rect 42536 36378 42564 36722
rect 46216 36378 46244 36722
rect 32220 36372 32272 36378
rect 32220 36314 32272 36320
rect 35348 36372 35400 36378
rect 35348 36314 35400 36320
rect 37372 36372 37424 36378
rect 37372 36314 37424 36320
rect 42524 36372 42576 36378
rect 42524 36314 42576 36320
rect 46204 36372 46256 36378
rect 46204 36314 46256 36320
rect 33324 36032 33376 36038
rect 33324 35974 33376 35980
rect 29552 35284 29604 35290
rect 29552 35226 29604 35232
rect 31668 35284 31720 35290
rect 31668 35226 31720 35232
rect 30380 35080 30432 35086
rect 30380 35022 30432 35028
rect 30656 35080 30708 35086
rect 30656 35022 30708 35028
rect 31852 35080 31904 35086
rect 31852 35022 31904 35028
rect 29276 35012 29328 35018
rect 29276 34954 29328 34960
rect 29184 34944 29236 34950
rect 29184 34886 29236 34892
rect 28816 34604 28868 34610
rect 28816 34546 28868 34552
rect 27804 33516 27856 33522
rect 27804 33458 27856 33464
rect 27160 33312 27212 33318
rect 27160 33254 27212 33260
rect 27816 32978 27844 33458
rect 27804 32972 27856 32978
rect 27804 32914 27856 32920
rect 26712 32842 26832 32858
rect 26712 32836 26844 32842
rect 26712 32830 26792 32836
rect 26792 32778 26844 32784
rect 27528 32836 27580 32842
rect 27528 32778 27580 32784
rect 28908 32836 28960 32842
rect 28908 32778 28960 32784
rect 26804 32570 26832 32778
rect 27160 32768 27212 32774
rect 27160 32710 27212 32716
rect 26792 32564 26844 32570
rect 26792 32506 26844 32512
rect 27172 32434 27200 32710
rect 27540 32570 27568 32778
rect 27252 32564 27304 32570
rect 27252 32506 27304 32512
rect 27528 32564 27580 32570
rect 27528 32506 27580 32512
rect 27160 32428 27212 32434
rect 27160 32370 27212 32376
rect 26516 32360 26568 32366
rect 26516 32302 26568 32308
rect 25596 31884 25648 31890
rect 25596 31826 25648 31832
rect 25412 31816 25464 31822
rect 25412 31758 25464 31764
rect 25424 31210 25452 31758
rect 25412 31204 25464 31210
rect 25412 31146 25464 31152
rect 25504 31136 25556 31142
rect 25504 31078 25556 31084
rect 25516 30734 25544 31078
rect 25608 30802 25636 31826
rect 26240 31816 26292 31822
rect 26240 31758 26292 31764
rect 25688 31340 25740 31346
rect 25688 31282 25740 31288
rect 25700 30938 25728 31282
rect 25688 30932 25740 30938
rect 25688 30874 25740 30880
rect 25596 30796 25648 30802
rect 25596 30738 25648 30744
rect 25504 30728 25556 30734
rect 25504 30670 25556 30676
rect 26252 30326 26280 31758
rect 26332 31272 26384 31278
rect 26332 31214 26384 31220
rect 26344 30938 26372 31214
rect 26332 30932 26384 30938
rect 26332 30874 26384 30880
rect 26240 30320 26292 30326
rect 26240 30262 26292 30268
rect 25228 30048 25280 30054
rect 25228 29990 25280 29996
rect 25240 29782 25268 29990
rect 25228 29776 25280 29782
rect 25228 29718 25280 29724
rect 27172 29578 27200 32370
rect 27264 31754 27292 32506
rect 28920 32026 28948 32778
rect 28908 32020 28960 32026
rect 28908 31962 28960 31968
rect 29000 31884 29052 31890
rect 29000 31826 29052 31832
rect 27264 31726 27476 31754
rect 27448 31482 27476 31726
rect 27436 31476 27488 31482
rect 27436 31418 27488 31424
rect 27448 30666 27476 31418
rect 29012 31414 29040 31826
rect 29000 31408 29052 31414
rect 29000 31350 29052 31356
rect 29012 30802 29040 31350
rect 29000 30796 29052 30802
rect 29000 30738 29052 30744
rect 27436 30660 27488 30666
rect 27436 30602 27488 30608
rect 27448 30394 27476 30602
rect 27436 30388 27488 30394
rect 27436 30330 27488 30336
rect 27160 29572 27212 29578
rect 27160 29514 27212 29520
rect 27172 29306 27200 29514
rect 27160 29300 27212 29306
rect 27160 29242 27212 29248
rect 26516 29096 26568 29102
rect 26516 29038 26568 29044
rect 25964 28960 26016 28966
rect 25964 28902 26016 28908
rect 25872 28620 25924 28626
rect 25872 28562 25924 28568
rect 25884 26926 25912 28562
rect 25976 28490 26004 28902
rect 26528 28762 26556 29038
rect 27448 29034 27476 30330
rect 28264 30184 28316 30190
rect 28264 30126 28316 30132
rect 28276 29102 28304 30126
rect 28816 29844 28868 29850
rect 28816 29786 28868 29792
rect 28632 29504 28684 29510
rect 28632 29446 28684 29452
rect 28264 29096 28316 29102
rect 28078 29064 28134 29073
rect 27436 29028 27488 29034
rect 28264 29038 28316 29044
rect 28078 28999 28080 29008
rect 27436 28970 27488 28976
rect 28132 28999 28134 29008
rect 28080 28970 28132 28976
rect 26516 28756 26568 28762
rect 26516 28698 26568 28704
rect 27448 28490 27476 28970
rect 25964 28484 26016 28490
rect 25964 28426 26016 28432
rect 27436 28484 27488 28490
rect 27436 28426 27488 28432
rect 27448 28218 27476 28426
rect 27436 28212 27488 28218
rect 27436 28154 27488 28160
rect 28276 28014 28304 29038
rect 28644 28150 28672 29446
rect 28828 28762 28856 29786
rect 29092 29776 29144 29782
rect 29092 29718 29144 29724
rect 29104 29238 29132 29718
rect 29092 29232 29144 29238
rect 29092 29174 29144 29180
rect 28816 28756 28868 28762
rect 28816 28698 28868 28704
rect 28632 28144 28684 28150
rect 28632 28086 28684 28092
rect 28264 28008 28316 28014
rect 28264 27950 28316 27956
rect 28276 27690 28304 27950
rect 28276 27662 28396 27690
rect 25320 26920 25372 26926
rect 25320 26862 25372 26868
rect 25872 26920 25924 26926
rect 25872 26862 25924 26868
rect 27620 26920 27672 26926
rect 27620 26862 27672 26868
rect 25332 26602 25360 26862
rect 25884 26790 25912 26862
rect 25872 26784 25924 26790
rect 25872 26726 25924 26732
rect 26792 26784 26844 26790
rect 26792 26726 26844 26732
rect 25240 26586 25360 26602
rect 25228 26580 25360 26586
rect 25280 26574 25360 26580
rect 25228 26522 25280 26528
rect 25240 26450 25544 26466
rect 25228 26444 25556 26450
rect 25280 26438 25504 26444
rect 25228 26386 25280 26392
rect 25504 26386 25556 26392
rect 25320 26376 25372 26382
rect 25320 26318 25372 26324
rect 25228 26240 25280 26246
rect 25228 26182 25280 26188
rect 25240 25906 25268 26182
rect 25228 25900 25280 25906
rect 25228 25842 25280 25848
rect 25240 25430 25268 25842
rect 25332 25770 25360 26318
rect 25320 25764 25372 25770
rect 25320 25706 25372 25712
rect 25516 25702 25544 26386
rect 25964 26376 26016 26382
rect 25962 26344 25964 26353
rect 26332 26376 26384 26382
rect 26016 26344 26018 26353
rect 26332 26318 26384 26324
rect 25962 26279 26018 26288
rect 26240 26308 26292 26314
rect 26240 26250 26292 26256
rect 26252 25838 26280 26250
rect 26240 25832 26292 25838
rect 26240 25774 26292 25780
rect 25412 25696 25464 25702
rect 25412 25638 25464 25644
rect 25504 25696 25556 25702
rect 25504 25638 25556 25644
rect 26148 25696 26200 25702
rect 26148 25638 26200 25644
rect 25228 25424 25280 25430
rect 25228 25366 25280 25372
rect 25228 25288 25280 25294
rect 25228 25230 25280 25236
rect 25136 24404 25188 24410
rect 25136 24346 25188 24352
rect 25240 24290 25268 25230
rect 25424 25226 25452 25638
rect 25688 25356 25740 25362
rect 25688 25298 25740 25304
rect 25412 25220 25464 25226
rect 25412 25162 25464 25168
rect 25700 24886 25728 25298
rect 26056 25152 26108 25158
rect 26056 25094 26108 25100
rect 25596 24880 25648 24886
rect 25318 24848 25374 24857
rect 25596 24822 25648 24828
rect 25688 24880 25740 24886
rect 25688 24822 25740 24828
rect 25318 24783 25320 24792
rect 25372 24783 25374 24792
rect 25320 24754 25372 24760
rect 25332 24614 25360 24754
rect 25608 24732 25636 24822
rect 25792 24818 26004 24834
rect 26068 24818 26096 25094
rect 25792 24812 26016 24818
rect 25792 24806 25964 24812
rect 25792 24732 25820 24806
rect 25964 24754 26016 24760
rect 26056 24812 26108 24818
rect 26056 24754 26108 24760
rect 25608 24704 25820 24732
rect 25412 24676 25464 24682
rect 25412 24618 25464 24624
rect 25320 24608 25372 24614
rect 25320 24550 25372 24556
rect 24872 24262 25084 24290
rect 25148 24262 25268 24290
rect 25320 24336 25372 24342
rect 25320 24278 25372 24284
rect 24872 23050 24900 24262
rect 25044 24200 25096 24206
rect 25044 24142 25096 24148
rect 24952 24064 25004 24070
rect 24952 24006 25004 24012
rect 24860 23044 24912 23050
rect 24860 22986 24912 22992
rect 24860 22228 24912 22234
rect 24860 22170 24912 22176
rect 24216 21956 24268 21962
rect 24268 21916 24348 21944
rect 24216 21898 24268 21904
rect 24124 21548 24176 21554
rect 24124 21490 24176 21496
rect 24136 21078 24164 21490
rect 24124 21072 24176 21078
rect 24124 21014 24176 21020
rect 24124 20868 24176 20874
rect 24124 20810 24176 20816
rect 24136 20466 24164 20810
rect 23848 20460 23900 20466
rect 23848 20402 23900 20408
rect 24032 20460 24084 20466
rect 24032 20402 24084 20408
rect 24124 20460 24176 20466
rect 24124 20402 24176 20408
rect 23572 20392 23624 20398
rect 23572 20334 23624 20340
rect 22652 19984 22704 19990
rect 22652 19926 22704 19932
rect 20444 19440 20496 19446
rect 20444 19382 20496 19388
rect 22192 19372 22244 19378
rect 21836 19320 22192 19334
rect 21836 19314 22244 19320
rect 22376 19372 22428 19378
rect 22376 19314 22428 19320
rect 23020 19372 23072 19378
rect 23020 19314 23072 19320
rect 23112 19372 23164 19378
rect 23112 19314 23164 19320
rect 23296 19372 23348 19378
rect 23296 19314 23348 19320
rect 21836 19306 22232 19314
rect 20076 19236 20128 19242
rect 20076 19178 20128 19184
rect 20076 18896 20128 18902
rect 20074 18864 20076 18873
rect 20128 18864 20130 18873
rect 20074 18799 20130 18808
rect 20260 18624 20312 18630
rect 20260 18566 20312 18572
rect 20272 18290 20300 18566
rect 21836 18426 21864 19306
rect 21916 19168 21968 19174
rect 21916 19110 21968 19116
rect 22100 19168 22152 19174
rect 22100 19110 22152 19116
rect 21928 18834 21956 19110
rect 21916 18828 21968 18834
rect 21916 18770 21968 18776
rect 21916 18692 21968 18698
rect 21916 18634 21968 18640
rect 21824 18420 21876 18426
rect 21824 18362 21876 18368
rect 20534 18320 20590 18329
rect 20260 18284 20312 18290
rect 20534 18255 20536 18264
rect 20260 18226 20312 18232
rect 20588 18255 20590 18264
rect 20536 18226 20588 18232
rect 20628 18216 20680 18222
rect 20628 18158 20680 18164
rect 20352 17196 20404 17202
rect 20352 17138 20404 17144
rect 20168 17128 20220 17134
rect 20168 17070 20220 17076
rect 19904 16612 20024 16640
rect 19708 16584 19760 16590
rect 19708 16526 19760 16532
rect 19616 16516 19668 16522
rect 19616 16458 19668 16464
rect 19524 16244 19576 16250
rect 19524 16186 19576 16192
rect 19524 16108 19576 16114
rect 19628 16096 19656 16458
rect 19720 16114 19748 16526
rect 19800 16244 19852 16250
rect 19800 16186 19852 16192
rect 19576 16068 19656 16096
rect 19524 16050 19576 16056
rect 18972 16040 19024 16046
rect 18972 15982 19024 15988
rect 18880 15700 18932 15706
rect 18880 15642 18932 15648
rect 18144 15360 18196 15366
rect 18144 15302 18196 15308
rect 18156 15094 18184 15302
rect 18052 15088 18104 15094
rect 18052 15030 18104 15036
rect 18144 15088 18196 15094
rect 18144 15030 18196 15036
rect 18064 14482 18092 15030
rect 19628 14958 19656 16068
rect 19708 16108 19760 16114
rect 19708 16050 19760 16056
rect 19720 15026 19748 16050
rect 19812 15502 19840 16186
rect 19800 15496 19852 15502
rect 19800 15438 19852 15444
rect 19708 15020 19760 15026
rect 19708 14962 19760 14968
rect 19616 14952 19668 14958
rect 19616 14894 19668 14900
rect 19812 14890 19840 15438
rect 19800 14884 19852 14890
rect 19800 14826 19852 14832
rect 19812 14634 19840 14826
rect 19720 14618 19840 14634
rect 19708 14612 19840 14618
rect 19760 14606 19840 14612
rect 19708 14554 19760 14560
rect 18052 14476 18104 14482
rect 18052 14418 18104 14424
rect 17960 14340 18012 14346
rect 17960 14282 18012 14288
rect 17972 13394 18000 14282
rect 18064 14074 18092 14418
rect 19432 14340 19484 14346
rect 19432 14282 19484 14288
rect 18144 14272 18196 14278
rect 18144 14214 18196 14220
rect 19156 14272 19208 14278
rect 19156 14214 19208 14220
rect 18052 14068 18104 14074
rect 18052 14010 18104 14016
rect 18156 13938 18184 14214
rect 19168 13938 19196 14214
rect 19444 14074 19472 14282
rect 19904 14278 19932 16612
rect 19984 16516 20036 16522
rect 19984 16458 20036 16464
rect 19996 15638 20024 16458
rect 20180 16046 20208 17070
rect 20364 16590 20392 17138
rect 20352 16584 20404 16590
rect 20352 16526 20404 16532
rect 20260 16244 20312 16250
rect 20260 16186 20312 16192
rect 20168 16040 20220 16046
rect 20168 15982 20220 15988
rect 20076 15972 20128 15978
rect 20076 15914 20128 15920
rect 20088 15706 20116 15914
rect 20076 15700 20128 15706
rect 20076 15642 20128 15648
rect 20168 15700 20220 15706
rect 20168 15642 20220 15648
rect 19984 15632 20036 15638
rect 19984 15574 20036 15580
rect 19996 15094 20024 15574
rect 20076 15496 20128 15502
rect 20076 15438 20128 15444
rect 20088 15162 20116 15438
rect 20076 15156 20128 15162
rect 20076 15098 20128 15104
rect 19984 15088 20036 15094
rect 19984 15030 20036 15036
rect 20180 15026 20208 15642
rect 20272 15502 20300 16186
rect 20260 15496 20312 15502
rect 20260 15438 20312 15444
rect 20364 15065 20392 16526
rect 20350 15056 20406 15065
rect 20168 15020 20220 15026
rect 20168 14962 20220 14968
rect 20260 15020 20312 15026
rect 20640 15026 20668 18158
rect 21640 17264 21692 17270
rect 21640 17206 21692 17212
rect 20812 16516 20864 16522
rect 20812 16458 20864 16464
rect 20824 16250 20852 16458
rect 21652 16250 21680 17206
rect 21928 16590 21956 18634
rect 22112 18154 22140 19110
rect 22192 18760 22244 18766
rect 22192 18702 22244 18708
rect 22100 18148 22152 18154
rect 22100 18090 22152 18096
rect 22112 17882 22140 18090
rect 22100 17876 22152 17882
rect 22100 17818 22152 17824
rect 22204 16658 22232 18702
rect 22388 18630 22416 19314
rect 23032 19174 23060 19314
rect 22560 19168 22612 19174
rect 22560 19110 22612 19116
rect 23020 19168 23072 19174
rect 23020 19110 23072 19116
rect 22572 18834 22600 19110
rect 22926 18864 22982 18873
rect 22560 18828 22612 18834
rect 22926 18799 22982 18808
rect 23020 18828 23072 18834
rect 22560 18770 22612 18776
rect 22376 18624 22428 18630
rect 22376 18566 22428 18572
rect 22466 18320 22522 18329
rect 22376 18284 22428 18290
rect 22466 18255 22468 18264
rect 22376 18226 22428 18232
rect 22520 18255 22522 18264
rect 22468 18226 22520 18232
rect 22388 18086 22416 18226
rect 22376 18080 22428 18086
rect 22376 18022 22428 18028
rect 22284 17264 22336 17270
rect 22284 17206 22336 17212
rect 22192 16652 22244 16658
rect 22192 16594 22244 16600
rect 21916 16584 21968 16590
rect 21916 16526 21968 16532
rect 20812 16244 20864 16250
rect 20812 16186 20864 16192
rect 21640 16244 21692 16250
rect 21640 16186 21692 16192
rect 21652 16046 21680 16186
rect 21640 16040 21692 16046
rect 21640 15982 21692 15988
rect 21548 15972 21600 15978
rect 21548 15914 21600 15920
rect 21560 15570 21588 15914
rect 21548 15564 21600 15570
rect 21548 15506 21600 15512
rect 20720 15360 20772 15366
rect 20720 15302 20772 15308
rect 21732 15360 21784 15366
rect 21732 15302 21784 15308
rect 20350 14991 20352 15000
rect 20260 14962 20312 14968
rect 20404 14991 20406 15000
rect 20628 15020 20680 15026
rect 20352 14962 20404 14968
rect 20628 14962 20680 14968
rect 20272 14618 20300 14962
rect 20444 14816 20496 14822
rect 20444 14758 20496 14764
rect 20260 14612 20312 14618
rect 20260 14554 20312 14560
rect 20456 14346 20484 14758
rect 20640 14482 20668 14962
rect 20732 14482 20760 15302
rect 21744 14482 21772 15302
rect 21928 15026 21956 16526
rect 22192 16448 22244 16454
rect 22296 16436 22324 17206
rect 22744 16992 22796 16998
rect 22744 16934 22796 16940
rect 22756 16794 22784 16934
rect 22744 16788 22796 16794
rect 22744 16730 22796 16736
rect 22244 16408 22324 16436
rect 22192 16390 22244 16396
rect 22296 16114 22324 16408
rect 22376 16448 22428 16454
rect 22376 16390 22428 16396
rect 22388 16250 22416 16390
rect 22376 16244 22428 16250
rect 22376 16186 22428 16192
rect 22192 16108 22244 16114
rect 22192 16050 22244 16056
rect 22284 16108 22336 16114
rect 22284 16050 22336 16056
rect 22468 16108 22520 16114
rect 22468 16050 22520 16056
rect 22204 15706 22232 16050
rect 22480 15978 22508 16050
rect 22940 15994 22968 18799
rect 23020 18770 23072 18776
rect 23032 18426 23060 18770
rect 23124 18426 23152 19314
rect 23308 18834 23336 19314
rect 23296 18828 23348 18834
rect 23296 18770 23348 18776
rect 23848 18624 23900 18630
rect 23848 18566 23900 18572
rect 23020 18420 23072 18426
rect 23020 18362 23072 18368
rect 23112 18420 23164 18426
rect 23112 18362 23164 18368
rect 23860 18290 23888 18566
rect 23572 18284 23624 18290
rect 23572 18226 23624 18232
rect 23848 18284 23900 18290
rect 23848 18226 23900 18232
rect 23296 18216 23348 18222
rect 23296 18158 23348 18164
rect 23112 17876 23164 17882
rect 23112 17818 23164 17824
rect 23020 17128 23072 17134
rect 23020 17070 23072 17076
rect 23032 16794 23060 17070
rect 23124 16998 23152 17818
rect 23204 17196 23256 17202
rect 23204 17138 23256 17144
rect 23112 16992 23164 16998
rect 23112 16934 23164 16940
rect 23020 16788 23072 16794
rect 23020 16730 23072 16736
rect 23032 16182 23060 16730
rect 23020 16176 23072 16182
rect 23020 16118 23072 16124
rect 22468 15972 22520 15978
rect 22468 15914 22520 15920
rect 22836 15972 22888 15978
rect 22940 15966 23060 15994
rect 22836 15914 22888 15920
rect 22192 15700 22244 15706
rect 22192 15642 22244 15648
rect 22560 15700 22612 15706
rect 22560 15642 22612 15648
rect 22192 15496 22244 15502
rect 22192 15438 22244 15444
rect 22376 15496 22428 15502
rect 22376 15438 22428 15444
rect 22100 15360 22152 15366
rect 22100 15302 22152 15308
rect 21916 15020 21968 15026
rect 21916 14962 21968 14968
rect 20628 14476 20680 14482
rect 20628 14418 20680 14424
rect 20720 14476 20772 14482
rect 20720 14418 20772 14424
rect 21732 14476 21784 14482
rect 21732 14418 21784 14424
rect 20444 14340 20496 14346
rect 20444 14282 20496 14288
rect 19892 14272 19944 14278
rect 19892 14214 19944 14220
rect 19432 14068 19484 14074
rect 19432 14010 19484 14016
rect 18144 13932 18196 13938
rect 18144 13874 18196 13880
rect 19156 13932 19208 13938
rect 19156 13874 19208 13880
rect 20260 13932 20312 13938
rect 20260 13874 20312 13880
rect 19340 13864 19392 13870
rect 20272 13841 20300 13874
rect 19340 13806 19392 13812
rect 20258 13832 20314 13841
rect 17316 13388 17368 13394
rect 17316 13330 17368 13336
rect 17960 13388 18012 13394
rect 17960 13330 18012 13336
rect 16856 13320 16908 13326
rect 16856 13262 16908 13268
rect 17040 13320 17092 13326
rect 17040 13262 17092 13268
rect 17224 13320 17276 13326
rect 17224 13262 17276 13268
rect 16868 12986 16896 13262
rect 17052 13190 17080 13262
rect 17040 13184 17092 13190
rect 17040 13126 17092 13132
rect 16856 12980 16908 12986
rect 16856 12922 16908 12928
rect 17052 12442 17080 13126
rect 17236 12986 17264 13262
rect 17328 13258 17356 13330
rect 17316 13252 17368 13258
rect 17316 13194 17368 13200
rect 17224 12980 17276 12986
rect 17224 12922 17276 12928
rect 17328 12850 17356 13194
rect 17960 13184 18012 13190
rect 17960 13126 18012 13132
rect 19248 13184 19300 13190
rect 19248 13126 19300 13132
rect 17316 12844 17368 12850
rect 17316 12786 17368 12792
rect 17040 12436 17092 12442
rect 17040 12378 17092 12384
rect 16764 12232 16816 12238
rect 16764 12174 16816 12180
rect 16948 12164 17000 12170
rect 16948 12106 17000 12112
rect 16396 11348 16448 11354
rect 16396 11290 16448 11296
rect 16672 11348 16724 11354
rect 16672 11290 16724 11296
rect 16960 11150 16988 12106
rect 17328 11762 17356 12786
rect 17972 12374 18000 13126
rect 19260 12918 19288 13126
rect 18420 12912 18472 12918
rect 18420 12854 18472 12860
rect 19248 12912 19300 12918
rect 19248 12854 19300 12860
rect 17960 12368 18012 12374
rect 17960 12310 18012 12316
rect 18432 12238 18460 12854
rect 19248 12368 19300 12374
rect 19248 12310 19300 12316
rect 19260 12238 19288 12310
rect 18420 12232 18472 12238
rect 18420 12174 18472 12180
rect 19248 12232 19300 12238
rect 19248 12174 19300 12180
rect 17500 12096 17552 12102
rect 17500 12038 17552 12044
rect 17868 12096 17920 12102
rect 17868 12038 17920 12044
rect 17512 11898 17540 12038
rect 17500 11892 17552 11898
rect 17500 11834 17552 11840
rect 17316 11756 17368 11762
rect 17316 11698 17368 11704
rect 17224 11280 17276 11286
rect 17224 11222 17276 11228
rect 16028 11144 16080 11150
rect 16028 11086 16080 11092
rect 16948 11144 17000 11150
rect 16948 11086 17000 11092
rect 15844 11076 15896 11082
rect 15844 11018 15896 11024
rect 15568 11008 15620 11014
rect 15568 10950 15620 10956
rect 15660 11008 15712 11014
rect 15660 10950 15712 10956
rect 13544 10804 13596 10810
rect 13544 10746 13596 10752
rect 13452 10464 13504 10470
rect 13452 10406 13504 10412
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 12348 9988 12400 9994
rect 12348 9930 12400 9936
rect 4874 9820 5182 9829
rect 4874 9818 4880 9820
rect 4936 9818 4960 9820
rect 5016 9818 5040 9820
rect 5096 9818 5120 9820
rect 5176 9818 5182 9820
rect 4936 9766 4938 9818
rect 5118 9766 5120 9818
rect 4874 9764 4880 9766
rect 4936 9764 4960 9766
rect 5016 9764 5040 9766
rect 5096 9764 5120 9766
rect 5176 9764 5182 9766
rect 4874 9755 5182 9764
rect 12360 9518 12388 9930
rect 13464 9654 13492 10406
rect 13556 10198 13584 10746
rect 13912 10736 13964 10742
rect 13912 10678 13964 10684
rect 13924 10198 13952 10678
rect 14832 10668 14884 10674
rect 14832 10610 14884 10616
rect 14096 10532 14148 10538
rect 14096 10474 14148 10480
rect 13544 10192 13596 10198
rect 13544 10134 13596 10140
rect 13912 10192 13964 10198
rect 13912 10134 13964 10140
rect 13924 9994 13952 10134
rect 14108 10062 14136 10474
rect 14844 10470 14872 10610
rect 15580 10538 15608 10950
rect 15672 10674 15700 10950
rect 15856 10742 15884 11018
rect 17132 11008 17184 11014
rect 17132 10950 17184 10956
rect 17144 10810 17172 10950
rect 17132 10804 17184 10810
rect 17132 10746 17184 10752
rect 15844 10736 15896 10742
rect 15844 10678 15896 10684
rect 15660 10668 15712 10674
rect 15660 10610 15712 10616
rect 16120 10600 16172 10606
rect 16120 10542 16172 10548
rect 15568 10532 15620 10538
rect 15568 10474 15620 10480
rect 14832 10464 14884 10470
rect 14832 10406 14884 10412
rect 14096 10056 14148 10062
rect 14096 9998 14148 10004
rect 13728 9988 13780 9994
rect 13728 9930 13780 9936
rect 13912 9988 13964 9994
rect 13912 9930 13964 9936
rect 13452 9648 13504 9654
rect 13452 9590 13504 9596
rect 13740 9518 13768 9930
rect 14844 9926 14872 10406
rect 16132 10062 16160 10542
rect 16120 10056 16172 10062
rect 16120 9998 16172 10004
rect 16856 9988 16908 9994
rect 16856 9930 16908 9936
rect 14832 9920 14884 9926
rect 14832 9862 14884 9868
rect 16764 9920 16816 9926
rect 16764 9862 16816 9868
rect 14844 9722 14872 9862
rect 14832 9716 14884 9722
rect 14832 9658 14884 9664
rect 15476 9648 15528 9654
rect 15476 9590 15528 9596
rect 12348 9512 12400 9518
rect 12348 9454 12400 9460
rect 12440 9512 12492 9518
rect 12440 9454 12492 9460
rect 13728 9512 13780 9518
rect 13728 9454 13780 9460
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 4874 8732 5182 8741
rect 4874 8730 4880 8732
rect 4936 8730 4960 8732
rect 5016 8730 5040 8732
rect 5096 8730 5120 8732
rect 5176 8730 5182 8732
rect 4936 8678 4938 8730
rect 5118 8678 5120 8730
rect 4874 8676 4880 8678
rect 4936 8676 4960 8678
rect 5016 8676 5040 8678
rect 5096 8676 5120 8678
rect 5176 8676 5182 8678
rect 4874 8667 5182 8676
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 12452 7954 12480 9454
rect 12072 7948 12124 7954
rect 12072 7890 12124 7896
rect 12440 7948 12492 7954
rect 12440 7890 12492 7896
rect 4874 7644 5182 7653
rect 4874 7642 4880 7644
rect 4936 7642 4960 7644
rect 5016 7642 5040 7644
rect 5096 7642 5120 7644
rect 5176 7642 5182 7644
rect 4936 7590 4938 7642
rect 5118 7590 5120 7642
rect 4874 7588 4880 7590
rect 4936 7588 4960 7590
rect 5016 7588 5040 7590
rect 5096 7588 5120 7590
rect 5176 7588 5182 7590
rect 4874 7579 5182 7588
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 4874 6556 5182 6565
rect 4874 6554 4880 6556
rect 4936 6554 4960 6556
rect 5016 6554 5040 6556
rect 5096 6554 5120 6556
rect 5176 6554 5182 6556
rect 4936 6502 4938 6554
rect 5118 6502 5120 6554
rect 4874 6500 4880 6502
rect 4936 6500 4960 6502
rect 5016 6500 5040 6502
rect 5096 6500 5120 6502
rect 5176 6500 5182 6502
rect 4874 6491 5182 6500
rect 12084 6254 12112 7890
rect 13740 7818 13768 9454
rect 15292 8492 15344 8498
rect 15292 8434 15344 8440
rect 15304 7936 15332 8434
rect 15384 7948 15436 7954
rect 15304 7908 15384 7936
rect 12440 7812 12492 7818
rect 12440 7754 12492 7760
rect 13728 7812 13780 7818
rect 13728 7754 13780 7760
rect 14372 7812 14424 7818
rect 14372 7754 14424 7760
rect 12452 7342 12480 7754
rect 12440 7336 12492 7342
rect 12440 7278 12492 7284
rect 12900 7336 12952 7342
rect 12900 7278 12952 7284
rect 12912 6474 12940 7278
rect 12912 6458 13032 6474
rect 12912 6452 13044 6458
rect 12912 6446 12992 6452
rect 12072 6248 12124 6254
rect 12072 6190 12124 6196
rect 12348 6112 12400 6118
rect 12348 6054 12400 6060
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 4874 5468 5182 5477
rect 4874 5466 4880 5468
rect 4936 5466 4960 5468
rect 5016 5466 5040 5468
rect 5096 5466 5120 5468
rect 5176 5466 5182 5468
rect 4936 5414 4938 5466
rect 5118 5414 5120 5466
rect 4874 5412 4880 5414
rect 4936 5412 4960 5414
rect 5016 5412 5040 5414
rect 5096 5412 5120 5414
rect 5176 5412 5182 5414
rect 4874 5403 5182 5412
rect 12360 5234 12388 6054
rect 12912 5710 12940 6446
rect 12992 6394 13044 6400
rect 13636 6384 13688 6390
rect 13556 6344 13636 6372
rect 12992 6248 13044 6254
rect 12992 6190 13044 6196
rect 13004 5914 13032 6190
rect 12992 5908 13044 5914
rect 12992 5850 13044 5856
rect 12900 5704 12952 5710
rect 12900 5646 12952 5652
rect 13556 5302 13584 6344
rect 13740 6372 13768 7754
rect 14004 7744 14056 7750
rect 14004 7686 14056 7692
rect 14016 7410 14044 7686
rect 14384 7546 14412 7754
rect 14372 7540 14424 7546
rect 14372 7482 14424 7488
rect 15304 7478 15332 7908
rect 15384 7890 15436 7896
rect 15488 7886 15516 9590
rect 16776 9586 16804 9862
rect 16868 9722 16896 9930
rect 16856 9716 16908 9722
rect 16856 9658 16908 9664
rect 16764 9580 16816 9586
rect 16764 9522 16816 9528
rect 16948 9580 17000 9586
rect 16948 9522 17000 9528
rect 16672 8968 16724 8974
rect 16672 8910 16724 8916
rect 15844 8492 15896 8498
rect 15844 8434 15896 8440
rect 16028 8492 16080 8498
rect 16028 8434 16080 8440
rect 15476 7880 15528 7886
rect 15476 7822 15528 7828
rect 15856 7750 15884 8434
rect 15936 8424 15988 8430
rect 15936 8366 15988 8372
rect 15948 7936 15976 8366
rect 16040 8090 16068 8434
rect 16684 8430 16712 8910
rect 16672 8424 16724 8430
rect 16672 8366 16724 8372
rect 16120 8288 16172 8294
rect 16120 8230 16172 8236
rect 16028 8084 16080 8090
rect 16028 8026 16080 8032
rect 15948 7908 16068 7936
rect 16040 7750 16068 7908
rect 15844 7744 15896 7750
rect 15844 7686 15896 7692
rect 16028 7744 16080 7750
rect 16028 7686 16080 7692
rect 15292 7472 15344 7478
rect 15292 7414 15344 7420
rect 14004 7404 14056 7410
rect 14004 7346 14056 7352
rect 14740 6792 14792 6798
rect 14740 6734 14792 6740
rect 14096 6656 14148 6662
rect 14096 6598 14148 6604
rect 13688 6344 13768 6372
rect 13636 6326 13688 6332
rect 14108 6322 14136 6598
rect 14752 6458 14780 6734
rect 14924 6656 14976 6662
rect 14924 6598 14976 6604
rect 14740 6452 14792 6458
rect 14740 6394 14792 6400
rect 14936 6390 14964 6598
rect 14924 6384 14976 6390
rect 14924 6326 14976 6332
rect 14004 6316 14056 6322
rect 14004 6258 14056 6264
rect 14096 6316 14148 6322
rect 14096 6258 14148 6264
rect 14556 6316 14608 6322
rect 14556 6258 14608 6264
rect 14832 6316 14884 6322
rect 14832 6258 14884 6264
rect 13912 6112 13964 6118
rect 13912 6054 13964 6060
rect 13924 5710 13952 6054
rect 14016 5710 14044 6258
rect 14280 6112 14332 6118
rect 14280 6054 14332 6060
rect 14292 5710 14320 6054
rect 14568 5914 14596 6258
rect 14740 6180 14792 6186
rect 14740 6122 14792 6128
rect 14556 5908 14608 5914
rect 14556 5850 14608 5856
rect 13912 5704 13964 5710
rect 13912 5646 13964 5652
rect 14004 5704 14056 5710
rect 14004 5646 14056 5652
rect 14280 5704 14332 5710
rect 14280 5646 14332 5652
rect 14752 5642 14780 6122
rect 14844 5914 14872 6258
rect 14832 5908 14884 5914
rect 14832 5850 14884 5856
rect 14556 5636 14608 5642
rect 14556 5578 14608 5584
rect 14740 5636 14792 5642
rect 14740 5578 14792 5584
rect 13820 5568 13872 5574
rect 13820 5510 13872 5516
rect 13544 5296 13596 5302
rect 13544 5238 13596 5244
rect 12348 5228 12400 5234
rect 12348 5170 12400 5176
rect 13832 5166 13860 5510
rect 14568 5370 14596 5578
rect 14752 5370 14780 5578
rect 15304 5370 15332 7414
rect 15856 7274 15884 7686
rect 15844 7268 15896 7274
rect 15844 7210 15896 7216
rect 15856 6934 15884 7210
rect 15844 6928 15896 6934
rect 15844 6870 15896 6876
rect 16040 6662 16068 7686
rect 16132 7410 16160 8230
rect 16212 8016 16264 8022
rect 16212 7958 16264 7964
rect 16684 7970 16712 8366
rect 16224 7410 16252 7958
rect 16488 7948 16540 7954
rect 16684 7942 16804 7970
rect 16488 7890 16540 7896
rect 16500 7410 16528 7890
rect 16672 7880 16724 7886
rect 16672 7822 16724 7828
rect 16684 7546 16712 7822
rect 16672 7540 16724 7546
rect 16672 7482 16724 7488
rect 16580 7472 16632 7478
rect 16580 7414 16632 7420
rect 16120 7404 16172 7410
rect 16120 7346 16172 7352
rect 16212 7404 16264 7410
rect 16212 7346 16264 7352
rect 16488 7404 16540 7410
rect 16488 7346 16540 7352
rect 16500 6866 16528 7346
rect 16592 6866 16620 7414
rect 16776 7206 16804 7942
rect 16856 7880 16908 7886
rect 16856 7822 16908 7828
rect 16764 7200 16816 7206
rect 16764 7142 16816 7148
rect 16488 6860 16540 6866
rect 16488 6802 16540 6808
rect 16580 6860 16632 6866
rect 16580 6802 16632 6808
rect 16776 6798 16804 7142
rect 16764 6792 16816 6798
rect 16764 6734 16816 6740
rect 16028 6656 16080 6662
rect 16028 6598 16080 6604
rect 16868 6322 16896 7822
rect 16960 7750 16988 9522
rect 17236 7886 17264 11222
rect 17880 11218 17908 12038
rect 19260 11898 19288 12174
rect 19248 11892 19300 11898
rect 19248 11834 19300 11840
rect 18236 11280 18288 11286
rect 18236 11222 18288 11228
rect 17868 11212 17920 11218
rect 17868 11154 17920 11160
rect 17316 11144 17368 11150
rect 17316 11086 17368 11092
rect 17328 10266 17356 11086
rect 17960 11008 18012 11014
rect 17960 10950 18012 10956
rect 17972 10742 18000 10950
rect 17960 10736 18012 10742
rect 17960 10678 18012 10684
rect 17972 10266 18000 10678
rect 18248 10674 18276 11222
rect 19248 11008 19300 11014
rect 19248 10950 19300 10956
rect 18052 10668 18104 10674
rect 18052 10610 18104 10616
rect 18236 10668 18288 10674
rect 18236 10610 18288 10616
rect 17316 10260 17368 10266
rect 17316 10202 17368 10208
rect 17960 10260 18012 10266
rect 17960 10202 18012 10208
rect 18064 10198 18092 10610
rect 19260 10606 19288 10950
rect 18328 10600 18380 10606
rect 18328 10542 18380 10548
rect 19248 10600 19300 10606
rect 19248 10542 19300 10548
rect 18052 10192 18104 10198
rect 18052 10134 18104 10140
rect 18340 10130 18368 10542
rect 18328 10124 18380 10130
rect 18328 10066 18380 10072
rect 17684 9920 17736 9926
rect 17684 9862 17736 9868
rect 17696 8566 17724 9862
rect 18144 8832 18196 8838
rect 18144 8774 18196 8780
rect 17684 8560 17736 8566
rect 17684 8502 17736 8508
rect 17696 7954 17724 8502
rect 18052 8424 18104 8430
rect 18052 8366 18104 8372
rect 17684 7948 17736 7954
rect 17684 7890 17736 7896
rect 17224 7880 17276 7886
rect 17224 7822 17276 7828
rect 16948 7744 17000 7750
rect 16948 7686 17000 7692
rect 17592 7744 17644 7750
rect 17592 7686 17644 7692
rect 16960 7342 16988 7686
rect 17604 7410 17632 7686
rect 18064 7546 18092 8366
rect 18156 7886 18184 8774
rect 18340 8634 18368 10066
rect 18328 8628 18380 8634
rect 18328 8570 18380 8576
rect 18340 8480 18368 8570
rect 18420 8492 18472 8498
rect 18340 8452 18420 8480
rect 18420 8434 18472 8440
rect 18144 7880 18196 7886
rect 18144 7822 18196 7828
rect 18052 7540 18104 7546
rect 18052 7482 18104 7488
rect 17408 7404 17460 7410
rect 17408 7346 17460 7352
rect 17592 7404 17644 7410
rect 17592 7346 17644 7352
rect 16948 7336 17000 7342
rect 17000 7284 17172 7290
rect 16948 7278 17172 7284
rect 16960 7274 17172 7278
rect 16960 7268 17184 7274
rect 16960 7262 17132 7268
rect 15384 6316 15436 6322
rect 15384 6258 15436 6264
rect 16856 6316 16908 6322
rect 16856 6258 16908 6264
rect 15396 5846 15424 6258
rect 15844 6248 15896 6254
rect 15844 6190 15896 6196
rect 15752 6112 15804 6118
rect 15752 6054 15804 6060
rect 15384 5840 15436 5846
rect 15384 5782 15436 5788
rect 15764 5778 15792 6054
rect 15856 5778 15884 6190
rect 15752 5772 15804 5778
rect 15752 5714 15804 5720
rect 15844 5772 15896 5778
rect 15844 5714 15896 5720
rect 16960 5710 16988 7262
rect 17132 7210 17184 7216
rect 17420 6730 17448 7346
rect 17684 6792 17736 6798
rect 17684 6734 17736 6740
rect 17408 6724 17460 6730
rect 17408 6666 17460 6672
rect 17420 6322 17448 6666
rect 17408 6316 17460 6322
rect 17408 6258 17460 6264
rect 17696 6254 17724 6734
rect 18144 6656 18196 6662
rect 18144 6598 18196 6604
rect 17684 6248 17736 6254
rect 17684 6190 17736 6196
rect 17500 6112 17552 6118
rect 17500 6054 17552 6060
rect 16580 5704 16632 5710
rect 16580 5646 16632 5652
rect 16948 5704 17000 5710
rect 16948 5646 17000 5652
rect 16488 5636 16540 5642
rect 16488 5578 16540 5584
rect 16212 5568 16264 5574
rect 16212 5510 16264 5516
rect 14556 5364 14608 5370
rect 14556 5306 14608 5312
rect 14740 5364 14792 5370
rect 14740 5306 14792 5312
rect 15292 5364 15344 5370
rect 15292 5306 15344 5312
rect 15568 5364 15620 5370
rect 15568 5306 15620 5312
rect 13820 5160 13872 5166
rect 13820 5102 13872 5108
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 15580 4690 15608 5306
rect 16224 5302 16252 5510
rect 16212 5296 16264 5302
rect 16212 5238 16264 5244
rect 16500 5250 16528 5578
rect 16592 5370 16620 5646
rect 17512 5642 17540 6054
rect 18156 5914 18184 6598
rect 19156 6248 19208 6254
rect 19156 6190 19208 6196
rect 19168 5914 19196 6190
rect 18144 5908 18196 5914
rect 18144 5850 18196 5856
rect 19156 5908 19208 5914
rect 19156 5850 19208 5856
rect 17776 5704 17828 5710
rect 17776 5646 17828 5652
rect 16856 5636 16908 5642
rect 16856 5578 16908 5584
rect 17500 5636 17552 5642
rect 17500 5578 17552 5584
rect 16580 5364 16632 5370
rect 16580 5306 16632 5312
rect 16500 5234 16620 5250
rect 16868 5234 16896 5578
rect 16500 5228 16632 5234
rect 16500 5222 16580 5228
rect 16580 5170 16632 5176
rect 16856 5228 16908 5234
rect 16856 5170 16908 5176
rect 17316 5228 17368 5234
rect 17316 5170 17368 5176
rect 16120 5160 16172 5166
rect 16120 5102 16172 5108
rect 15568 4684 15620 4690
rect 15568 4626 15620 4632
rect 16132 4554 16160 5102
rect 16120 4548 16172 4554
rect 16120 4490 16172 4496
rect 17328 4486 17356 5170
rect 17788 4826 17816 5646
rect 17776 4820 17828 4826
rect 17776 4762 17828 4768
rect 16672 4480 16724 4486
rect 16672 4422 16724 4428
rect 17316 4480 17368 4486
rect 17316 4422 17368 4428
rect 4874 4380 5182 4389
rect 4874 4378 4880 4380
rect 4936 4378 4960 4380
rect 5016 4378 5040 4380
rect 5096 4378 5120 4380
rect 5176 4378 5182 4380
rect 4936 4326 4938 4378
rect 5118 4326 5120 4378
rect 4874 4324 4880 4326
rect 4936 4324 4960 4326
rect 5016 4324 5040 4326
rect 5096 4324 5120 4326
rect 5176 4324 5182 4326
rect 4874 4315 5182 4324
rect 16684 4146 16712 4422
rect 17328 4146 17356 4422
rect 16672 4140 16724 4146
rect 16672 4082 16724 4088
rect 17316 4140 17368 4146
rect 17316 4082 17368 4088
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 4874 3292 5182 3301
rect 4874 3290 4880 3292
rect 4936 3290 4960 3292
rect 5016 3290 5040 3292
rect 5096 3290 5120 3292
rect 5176 3290 5182 3292
rect 4936 3238 4938 3290
rect 5118 3238 5120 3290
rect 4874 3236 4880 3238
rect 4936 3236 4960 3238
rect 5016 3236 5040 3238
rect 5096 3236 5120 3238
rect 5176 3236 5182 3238
rect 4874 3227 5182 3236
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 19352 2650 19380 13806
rect 20258 13767 20314 13776
rect 19984 13728 20036 13734
rect 19984 13670 20036 13676
rect 19800 12844 19852 12850
rect 19800 12786 19852 12792
rect 19616 12640 19668 12646
rect 19616 12582 19668 12588
rect 19708 12640 19760 12646
rect 19708 12582 19760 12588
rect 19628 11830 19656 12582
rect 19720 12238 19748 12582
rect 19812 12442 19840 12786
rect 19800 12436 19852 12442
rect 19800 12378 19852 12384
rect 19708 12232 19760 12238
rect 19708 12174 19760 12180
rect 19616 11824 19668 11830
rect 19616 11766 19668 11772
rect 19892 11144 19944 11150
rect 19892 11086 19944 11092
rect 19904 10470 19932 11086
rect 19996 10742 20024 13670
rect 20640 13326 20668 14418
rect 21456 14408 21508 14414
rect 21456 14350 21508 14356
rect 21468 13938 21496 14350
rect 21928 14328 21956 14962
rect 22008 14340 22060 14346
rect 21928 14300 22008 14328
rect 22008 14282 22060 14288
rect 22112 14006 22140 15302
rect 22204 15162 22232 15438
rect 22388 15162 22416 15438
rect 22192 15156 22244 15162
rect 22192 15098 22244 15104
rect 22376 15156 22428 15162
rect 22376 15098 22428 15104
rect 22572 15026 22600 15642
rect 22848 15065 22876 15914
rect 22928 15496 22980 15502
rect 22928 15438 22980 15444
rect 22834 15056 22890 15065
rect 22560 15020 22612 15026
rect 22560 14962 22612 14968
rect 22744 15020 22796 15026
rect 22834 14991 22836 15000
rect 22744 14962 22796 14968
rect 22888 14991 22890 15000
rect 22836 14962 22888 14968
rect 22756 14890 22784 14962
rect 22744 14884 22796 14890
rect 22744 14826 22796 14832
rect 22940 14618 22968 15438
rect 23032 15026 23060 15966
rect 23124 15502 23152 16934
rect 23216 16250 23244 17138
rect 23204 16244 23256 16250
rect 23204 16186 23256 16192
rect 23308 16114 23336 18158
rect 23584 18086 23612 18226
rect 23572 18080 23624 18086
rect 24320 18034 24348 21916
rect 24400 21616 24452 21622
rect 24584 21616 24636 21622
rect 24452 21564 24584 21570
rect 24400 21558 24636 21564
rect 24412 21542 24624 21558
rect 24872 21554 24900 22170
rect 24860 21548 24912 21554
rect 24412 18766 24440 21542
rect 24860 21490 24912 21496
rect 24584 21344 24636 21350
rect 24584 21286 24636 21292
rect 24596 20942 24624 21286
rect 24584 20936 24636 20942
rect 24584 20878 24636 20884
rect 24860 20868 24912 20874
rect 24860 20810 24912 20816
rect 24872 20777 24900 20810
rect 24858 20768 24914 20777
rect 24858 20703 24914 20712
rect 24768 20256 24820 20262
rect 24768 20198 24820 20204
rect 24780 19446 24808 20198
rect 24872 19854 24900 20703
rect 24860 19848 24912 19854
rect 24860 19790 24912 19796
rect 24768 19440 24820 19446
rect 24768 19382 24820 19388
rect 24584 19304 24636 19310
rect 24584 19246 24636 19252
rect 24596 19145 24624 19246
rect 24582 19136 24638 19145
rect 24582 19071 24638 19080
rect 24858 19136 24914 19145
rect 24858 19071 24914 19080
rect 24400 18760 24452 18766
rect 24400 18702 24452 18708
rect 24768 18692 24820 18698
rect 24768 18634 24820 18640
rect 24584 18624 24636 18630
rect 24584 18566 24636 18572
rect 24596 18154 24624 18566
rect 24676 18420 24728 18426
rect 24676 18362 24728 18368
rect 24584 18148 24636 18154
rect 24584 18090 24636 18096
rect 23572 18022 23624 18028
rect 23296 16108 23348 16114
rect 23216 16068 23296 16096
rect 23112 15496 23164 15502
rect 23112 15438 23164 15444
rect 23124 15162 23152 15438
rect 23216 15162 23244 16068
rect 23296 16050 23348 16056
rect 23480 16108 23532 16114
rect 23584 16096 23612 18022
rect 23952 18006 24348 18034
rect 23664 17060 23716 17066
rect 23664 17002 23716 17008
rect 23676 16454 23704 17002
rect 23664 16448 23716 16454
rect 23664 16390 23716 16396
rect 23676 16114 23704 16390
rect 23532 16068 23612 16096
rect 23664 16108 23716 16114
rect 23480 16050 23532 16056
rect 23664 16050 23716 16056
rect 23848 16108 23900 16114
rect 23848 16050 23900 16056
rect 23492 15706 23520 16050
rect 23756 15972 23808 15978
rect 23756 15914 23808 15920
rect 23480 15700 23532 15706
rect 23480 15642 23532 15648
rect 23294 15600 23350 15609
rect 23294 15535 23350 15544
rect 23308 15434 23336 15535
rect 23388 15496 23440 15502
rect 23388 15438 23440 15444
rect 23296 15428 23348 15434
rect 23296 15370 23348 15376
rect 23112 15156 23164 15162
rect 23112 15098 23164 15104
rect 23204 15156 23256 15162
rect 23204 15098 23256 15104
rect 23020 15020 23072 15026
rect 23020 14962 23072 14968
rect 22928 14612 22980 14618
rect 22928 14554 22980 14560
rect 23124 14550 23152 15098
rect 23112 14544 23164 14550
rect 23112 14486 23164 14492
rect 23216 14414 23244 15098
rect 23400 14890 23428 15438
rect 23492 15366 23520 15642
rect 23572 15564 23624 15570
rect 23572 15506 23624 15512
rect 23480 15360 23532 15366
rect 23480 15302 23532 15308
rect 23388 14884 23440 14890
rect 23388 14826 23440 14832
rect 23204 14408 23256 14414
rect 23204 14350 23256 14356
rect 22192 14340 22244 14346
rect 22192 14282 22244 14288
rect 22204 14006 22232 14282
rect 22100 14000 22152 14006
rect 22100 13942 22152 13948
rect 22192 14000 22244 14006
rect 22192 13942 22244 13948
rect 21456 13932 21508 13938
rect 21456 13874 21508 13880
rect 20628 13320 20680 13326
rect 20628 13262 20680 13268
rect 21088 12776 21140 12782
rect 21088 12718 21140 12724
rect 20904 12096 20956 12102
rect 21100 12050 21128 12718
rect 22204 12170 22232 13942
rect 23400 13802 23428 14826
rect 23492 14278 23520 15302
rect 23584 14414 23612 15506
rect 23572 14408 23624 14414
rect 23572 14350 23624 14356
rect 23768 14346 23796 15914
rect 23860 15570 23888 16050
rect 23848 15564 23900 15570
rect 23848 15506 23900 15512
rect 23756 14340 23808 14346
rect 23756 14282 23808 14288
rect 23480 14272 23532 14278
rect 23480 14214 23532 14220
rect 23848 13932 23900 13938
rect 23848 13874 23900 13880
rect 23388 13796 23440 13802
rect 23388 13738 23440 13744
rect 23860 13394 23888 13874
rect 23848 13388 23900 13394
rect 23848 13330 23900 13336
rect 23952 13326 23980 18006
rect 24596 17882 24624 18090
rect 24584 17876 24636 17882
rect 24584 17818 24636 17824
rect 24596 17202 24624 17818
rect 24688 17270 24716 18362
rect 24780 18358 24808 18634
rect 24768 18352 24820 18358
rect 24768 18294 24820 18300
rect 24676 17264 24728 17270
rect 24676 17206 24728 17212
rect 24032 17196 24084 17202
rect 24032 17138 24084 17144
rect 24584 17196 24636 17202
rect 24584 17138 24636 17144
rect 24044 15570 24072 17138
rect 24216 16992 24268 16998
rect 24216 16934 24268 16940
rect 24400 16992 24452 16998
rect 24400 16934 24452 16940
rect 24674 16960 24730 16969
rect 24124 16652 24176 16658
rect 24124 16594 24176 16600
rect 24032 15564 24084 15570
rect 24032 15506 24084 15512
rect 24136 15434 24164 16594
rect 24228 15706 24256 16934
rect 24412 16590 24440 16934
rect 24674 16895 24730 16904
rect 24400 16584 24452 16590
rect 24400 16526 24452 16532
rect 24492 16584 24544 16590
rect 24492 16526 24544 16532
rect 24400 16448 24452 16454
rect 24400 16390 24452 16396
rect 24216 15700 24268 15706
rect 24216 15642 24268 15648
rect 24124 15428 24176 15434
rect 24124 15370 24176 15376
rect 24136 15026 24164 15370
rect 24124 15020 24176 15026
rect 24124 14962 24176 14968
rect 24136 14006 24164 14962
rect 24216 14408 24268 14414
rect 24216 14350 24268 14356
rect 24124 14000 24176 14006
rect 24124 13942 24176 13948
rect 24228 13938 24256 14350
rect 24308 14272 24360 14278
rect 24308 14214 24360 14220
rect 24320 13938 24348 14214
rect 24412 13938 24440 16390
rect 24504 15638 24532 16526
rect 24584 16516 24636 16522
rect 24584 16458 24636 16464
rect 24596 15910 24624 16458
rect 24688 16182 24716 16895
rect 24676 16176 24728 16182
rect 24676 16118 24728 16124
rect 24768 16108 24820 16114
rect 24768 16050 24820 16056
rect 24780 15910 24808 16050
rect 24584 15904 24636 15910
rect 24584 15846 24636 15852
rect 24768 15904 24820 15910
rect 24768 15846 24820 15852
rect 24872 15706 24900 19071
rect 24964 18834 24992 24006
rect 25056 23866 25084 24142
rect 25044 23860 25096 23866
rect 25044 23802 25096 23808
rect 25148 22094 25176 24262
rect 25228 24200 25280 24206
rect 25228 24142 25280 24148
rect 25240 23866 25268 24142
rect 25228 23860 25280 23866
rect 25228 23802 25280 23808
rect 25332 23730 25360 24278
rect 25424 24206 25452 24618
rect 25504 24608 25556 24614
rect 25504 24550 25556 24556
rect 25516 24206 25544 24550
rect 25412 24200 25464 24206
rect 25412 24142 25464 24148
rect 25504 24200 25556 24206
rect 25504 24142 25556 24148
rect 25608 24070 25636 24704
rect 25964 24676 26016 24682
rect 25964 24618 26016 24624
rect 25778 24440 25834 24449
rect 25778 24375 25834 24384
rect 25792 24206 25820 24375
rect 25780 24200 25832 24206
rect 25780 24142 25832 24148
rect 25596 24064 25648 24070
rect 25410 24032 25466 24041
rect 25596 24006 25648 24012
rect 25688 24064 25740 24070
rect 25688 24006 25740 24012
rect 25410 23967 25466 23976
rect 25320 23724 25372 23730
rect 25320 23666 25372 23672
rect 25320 23520 25372 23526
rect 25320 23462 25372 23468
rect 25056 22066 25176 22094
rect 25056 19854 25084 22066
rect 25228 20460 25280 20466
rect 25228 20402 25280 20408
rect 25136 20392 25188 20398
rect 25136 20334 25188 20340
rect 25148 20074 25176 20334
rect 25240 20262 25268 20402
rect 25228 20256 25280 20262
rect 25228 20198 25280 20204
rect 25148 20046 25268 20074
rect 25044 19848 25096 19854
rect 25044 19790 25096 19796
rect 25136 19780 25188 19786
rect 25136 19722 25188 19728
rect 25044 19168 25096 19174
rect 25044 19110 25096 19116
rect 24952 18828 25004 18834
rect 24952 18770 25004 18776
rect 24964 18426 24992 18770
rect 25056 18766 25084 19110
rect 25148 19009 25176 19722
rect 25134 19000 25190 19009
rect 25134 18935 25190 18944
rect 25148 18902 25176 18935
rect 25136 18896 25188 18902
rect 25136 18838 25188 18844
rect 25044 18760 25096 18766
rect 25044 18702 25096 18708
rect 25136 18692 25188 18698
rect 25136 18634 25188 18640
rect 25044 18624 25096 18630
rect 25044 18566 25096 18572
rect 24952 18420 25004 18426
rect 24952 18362 25004 18368
rect 25056 18222 25084 18566
rect 25148 18290 25176 18634
rect 25136 18284 25188 18290
rect 25136 18226 25188 18232
rect 25044 18216 25096 18222
rect 25044 18158 25096 18164
rect 25056 17610 25084 18158
rect 25044 17604 25096 17610
rect 25044 17546 25096 17552
rect 25240 17218 25268 20046
rect 25332 19938 25360 23462
rect 25424 20602 25452 23967
rect 25594 23896 25650 23905
rect 25594 23831 25650 23840
rect 25608 23798 25636 23831
rect 25596 23792 25648 23798
rect 25596 23734 25648 23740
rect 25700 23730 25728 24006
rect 25688 23724 25740 23730
rect 25688 23666 25740 23672
rect 25596 22636 25648 22642
rect 25596 22578 25648 22584
rect 25608 22234 25636 22578
rect 25596 22228 25648 22234
rect 25596 22170 25648 22176
rect 25596 21344 25648 21350
rect 25596 21286 25648 21292
rect 25504 21004 25556 21010
rect 25504 20946 25556 20952
rect 25412 20596 25464 20602
rect 25412 20538 25464 20544
rect 25516 20466 25544 20946
rect 25608 20874 25636 21286
rect 25596 20868 25648 20874
rect 25596 20810 25648 20816
rect 25412 20460 25464 20466
rect 25412 20402 25464 20408
rect 25504 20460 25556 20466
rect 25504 20402 25556 20408
rect 25424 20058 25452 20402
rect 25596 20256 25648 20262
rect 25596 20198 25648 20204
rect 25412 20052 25464 20058
rect 25412 19994 25464 20000
rect 25332 19910 25452 19938
rect 25320 19848 25372 19854
rect 25320 19790 25372 19796
rect 25332 18970 25360 19790
rect 25320 18964 25372 18970
rect 25320 18906 25372 18912
rect 25424 18766 25452 19910
rect 25504 19916 25556 19922
rect 25504 19858 25556 19864
rect 25412 18760 25464 18766
rect 25412 18702 25464 18708
rect 25424 18601 25452 18702
rect 25410 18592 25466 18601
rect 25410 18527 25466 18536
rect 24952 17196 25004 17202
rect 24952 17138 25004 17144
rect 25148 17190 25268 17218
rect 24964 16250 24992 17138
rect 25044 16788 25096 16794
rect 25044 16730 25096 16736
rect 25056 16697 25084 16730
rect 25042 16688 25098 16697
rect 25042 16623 25098 16632
rect 25044 16584 25096 16590
rect 25042 16552 25044 16561
rect 25096 16552 25098 16561
rect 25042 16487 25098 16496
rect 24952 16244 25004 16250
rect 24952 16186 25004 16192
rect 25056 16114 25084 16487
rect 25148 16250 25176 17190
rect 25228 17128 25280 17134
rect 25228 17070 25280 17076
rect 25240 16726 25268 17070
rect 25412 16992 25464 16998
rect 25412 16934 25464 16940
rect 25318 16824 25374 16833
rect 25318 16759 25320 16768
rect 25372 16759 25374 16768
rect 25320 16730 25372 16736
rect 25228 16720 25280 16726
rect 25228 16662 25280 16668
rect 25320 16584 25372 16590
rect 25320 16526 25372 16532
rect 25136 16244 25188 16250
rect 25136 16186 25188 16192
rect 25044 16108 25096 16114
rect 25044 16050 25096 16056
rect 25148 16046 25176 16186
rect 25136 16040 25188 16046
rect 25136 15982 25188 15988
rect 24676 15700 24728 15706
rect 24676 15642 24728 15648
rect 24860 15700 24912 15706
rect 24860 15642 24912 15648
rect 24492 15632 24544 15638
rect 24492 15574 24544 15580
rect 24492 15496 24544 15502
rect 24492 15438 24544 15444
rect 24216 13932 24268 13938
rect 24216 13874 24268 13880
rect 24308 13932 24360 13938
rect 24308 13874 24360 13880
rect 24400 13932 24452 13938
rect 24400 13874 24452 13880
rect 23940 13320 23992 13326
rect 23940 13262 23992 13268
rect 24228 12918 24256 13874
rect 24320 13530 24348 13874
rect 24308 13524 24360 13530
rect 24308 13466 24360 13472
rect 24412 13326 24440 13874
rect 24504 13870 24532 15438
rect 24688 14414 24716 15642
rect 24768 15564 24820 15570
rect 24768 15506 24820 15512
rect 24780 14618 24808 15506
rect 24860 15020 24912 15026
rect 24860 14962 24912 14968
rect 24768 14612 24820 14618
rect 24768 14554 24820 14560
rect 24676 14408 24728 14414
rect 24676 14350 24728 14356
rect 24584 14068 24636 14074
rect 24584 14010 24636 14016
rect 24492 13864 24544 13870
rect 24492 13806 24544 13812
rect 24400 13320 24452 13326
rect 24400 13262 24452 13268
rect 24412 12986 24440 13262
rect 24596 12986 24624 14010
rect 24780 13954 24808 14554
rect 24688 13938 24808 13954
rect 24872 13938 24900 14962
rect 25332 14958 25360 16526
rect 25424 16454 25452 16934
rect 25516 16522 25544 19858
rect 25608 19281 25636 20198
rect 25700 20058 25728 23666
rect 25792 22094 25820 24142
rect 25872 24132 25924 24138
rect 25872 24074 25924 24080
rect 25884 23633 25912 24074
rect 25870 23624 25926 23633
rect 25870 23559 25926 23568
rect 25976 23526 26004 24618
rect 26056 24336 26108 24342
rect 26056 24278 26108 24284
rect 25964 23520 26016 23526
rect 25964 23462 26016 23468
rect 26068 23066 26096 24278
rect 26160 23304 26188 25638
rect 26252 25430 26280 25774
rect 26240 25424 26292 25430
rect 26240 25366 26292 25372
rect 26344 24954 26372 26318
rect 26804 26314 26832 26726
rect 26792 26308 26844 26314
rect 26792 26250 26844 26256
rect 26516 25968 26568 25974
rect 26516 25910 26568 25916
rect 26332 24948 26384 24954
rect 26332 24890 26384 24896
rect 26332 24608 26384 24614
rect 26332 24550 26384 24556
rect 26344 24313 26372 24550
rect 26528 24449 26556 25910
rect 27632 25906 27660 26862
rect 28368 26790 28396 27662
rect 28908 27124 28960 27130
rect 28908 27066 28960 27072
rect 28356 26784 28408 26790
rect 28356 26726 28408 26732
rect 28632 26784 28684 26790
rect 28632 26726 28684 26732
rect 27988 26512 28040 26518
rect 27988 26454 28040 26460
rect 27804 26444 27856 26450
rect 27804 26386 27856 26392
rect 27712 26376 27764 26382
rect 27710 26344 27712 26353
rect 27764 26344 27766 26353
rect 27710 26279 27766 26288
rect 27712 26240 27764 26246
rect 27712 26182 27764 26188
rect 27620 25900 27672 25906
rect 27620 25842 27672 25848
rect 26976 25832 27028 25838
rect 26976 25774 27028 25780
rect 26514 24440 26570 24449
rect 26514 24375 26516 24384
rect 26568 24375 26570 24384
rect 26516 24346 26568 24352
rect 26330 24304 26386 24313
rect 26330 24239 26386 24248
rect 26424 24268 26476 24274
rect 26424 24210 26476 24216
rect 26330 24168 26386 24177
rect 26330 24103 26332 24112
rect 26384 24103 26386 24112
rect 26332 24074 26384 24080
rect 26436 23798 26464 24210
rect 26988 24206 27016 25774
rect 27724 25226 27752 26182
rect 27816 25974 27844 26386
rect 27804 25968 27856 25974
rect 27804 25910 27856 25916
rect 28000 25906 28028 26454
rect 28368 26314 28396 26726
rect 28446 26344 28502 26353
rect 28356 26308 28408 26314
rect 28446 26279 28502 26288
rect 28356 26250 28408 26256
rect 28368 25906 28396 26250
rect 27988 25900 28040 25906
rect 27988 25842 28040 25848
rect 28356 25900 28408 25906
rect 28356 25842 28408 25848
rect 28460 25294 28488 26279
rect 28540 26240 28592 26246
rect 28540 26182 28592 26188
rect 28552 25974 28580 26182
rect 28540 25968 28592 25974
rect 28540 25910 28592 25916
rect 28644 25838 28672 26726
rect 28816 26376 28868 26382
rect 28816 26318 28868 26324
rect 28632 25832 28684 25838
rect 28632 25774 28684 25780
rect 28356 25288 28408 25294
rect 28356 25230 28408 25236
rect 28448 25288 28500 25294
rect 28448 25230 28500 25236
rect 27712 25220 27764 25226
rect 27712 25162 27764 25168
rect 27344 25152 27396 25158
rect 27344 25094 27396 25100
rect 26976 24200 27028 24206
rect 26976 24142 27028 24148
rect 26608 23860 26660 23866
rect 26608 23802 26660 23808
rect 26424 23792 26476 23798
rect 26424 23734 26476 23740
rect 26160 23276 26280 23304
rect 26068 23038 26188 23066
rect 26056 22976 26108 22982
rect 26056 22918 26108 22924
rect 25872 22500 25924 22506
rect 25872 22442 25924 22448
rect 25884 22234 25912 22442
rect 25872 22228 25924 22234
rect 25872 22170 25924 22176
rect 25792 22066 26004 22094
rect 25872 21480 25924 21486
rect 25872 21422 25924 21428
rect 25884 21146 25912 21422
rect 25872 21140 25924 21146
rect 25872 21082 25924 21088
rect 25884 20806 25912 21082
rect 25872 20800 25924 20806
rect 25872 20742 25924 20748
rect 25688 20052 25740 20058
rect 25688 19994 25740 20000
rect 25700 19786 25728 19994
rect 25688 19780 25740 19786
rect 25688 19722 25740 19728
rect 25700 19514 25728 19722
rect 25688 19508 25740 19514
rect 25688 19450 25740 19456
rect 25884 19334 25912 20742
rect 25792 19306 25912 19334
rect 25594 19272 25650 19281
rect 25594 19207 25650 19216
rect 25792 19122 25820 19306
rect 25872 19236 25924 19242
rect 25872 19178 25924 19184
rect 25884 19145 25912 19178
rect 25976 19174 26004 22066
rect 26068 21690 26096 22918
rect 26056 21684 26108 21690
rect 26056 21626 26108 21632
rect 26068 21010 26096 21626
rect 26056 21004 26108 21010
rect 26056 20946 26108 20952
rect 26160 20584 26188 23038
rect 26252 22506 26280 23276
rect 26332 22976 26384 22982
rect 26332 22918 26384 22924
rect 26344 22710 26372 22918
rect 26332 22704 26384 22710
rect 26332 22646 26384 22652
rect 26240 22500 26292 22506
rect 26240 22442 26292 22448
rect 26252 21418 26280 22442
rect 26332 22432 26384 22438
rect 26332 22374 26384 22380
rect 26344 22234 26372 22374
rect 26332 22228 26384 22234
rect 26332 22170 26384 22176
rect 26620 22094 26648 23802
rect 26700 23724 26752 23730
rect 26700 23666 26752 23672
rect 26712 23254 26740 23666
rect 26700 23248 26752 23254
rect 26700 23190 26752 23196
rect 26988 22642 27016 24142
rect 27068 23792 27120 23798
rect 27066 23760 27068 23769
rect 27120 23760 27122 23769
rect 27066 23695 27122 23704
rect 26976 22636 27028 22642
rect 26976 22578 27028 22584
rect 26528 22066 26648 22094
rect 26240 21412 26292 21418
rect 26240 21354 26292 21360
rect 26252 21078 26280 21354
rect 26332 21344 26384 21350
rect 26332 21286 26384 21292
rect 26240 21072 26292 21078
rect 26240 21014 26292 21020
rect 26160 20556 26280 20584
rect 26146 20496 26202 20505
rect 26146 20431 26148 20440
rect 26200 20431 26202 20440
rect 26148 20402 26200 20408
rect 26056 20256 26108 20262
rect 26056 20198 26108 20204
rect 26068 20058 26096 20198
rect 26056 20052 26108 20058
rect 26056 19994 26108 20000
rect 26252 19938 26280 20556
rect 26344 20534 26372 21286
rect 26332 20528 26384 20534
rect 26332 20470 26384 20476
rect 26528 20330 26556 22066
rect 26608 21548 26660 21554
rect 26608 21490 26660 21496
rect 26620 21146 26648 21490
rect 26608 21140 26660 21146
rect 26608 21082 26660 21088
rect 26700 20596 26752 20602
rect 26700 20538 26752 20544
rect 26516 20324 26568 20330
rect 26516 20266 26568 20272
rect 26608 20256 26660 20262
rect 26608 20198 26660 20204
rect 26068 19910 26280 19938
rect 26424 19984 26476 19990
rect 26424 19926 26476 19932
rect 26068 19334 26096 19910
rect 26332 19848 26384 19854
rect 26252 19808 26332 19836
rect 26252 19514 26280 19808
rect 26332 19790 26384 19796
rect 26436 19718 26464 19926
rect 26620 19922 26648 20198
rect 26608 19916 26660 19922
rect 26608 19858 26660 19864
rect 26608 19780 26660 19786
rect 26608 19722 26660 19728
rect 26332 19712 26384 19718
rect 26332 19654 26384 19660
rect 26424 19712 26476 19718
rect 26424 19654 26476 19660
rect 26148 19508 26200 19514
rect 26148 19450 26200 19456
rect 26240 19508 26292 19514
rect 26240 19450 26292 19456
rect 26160 19394 26188 19450
rect 26160 19366 26280 19394
rect 26068 19306 26188 19334
rect 25964 19168 26016 19174
rect 25744 19094 25820 19122
rect 25870 19136 25926 19145
rect 25744 18952 25772 19094
rect 25964 19110 26016 19116
rect 25870 19071 25926 19080
rect 25700 18924 25772 18952
rect 25700 18884 25728 18924
rect 25608 18856 25728 18884
rect 25608 18714 25636 18856
rect 26160 18816 26188 19306
rect 26069 18788 26188 18816
rect 25872 18760 25924 18766
rect 25608 18708 25872 18714
rect 26069 18748 26097 18788
rect 25608 18702 25924 18708
rect 25976 18720 26097 18748
rect 26146 18728 26202 18737
rect 25608 18686 25912 18702
rect 25792 17882 25820 18686
rect 25976 18630 26004 18720
rect 26146 18663 26202 18672
rect 26160 18630 26188 18663
rect 25964 18624 26016 18630
rect 25964 18566 26016 18572
rect 26148 18624 26200 18630
rect 26148 18566 26200 18572
rect 25976 18068 26004 18566
rect 26056 18080 26108 18086
rect 25976 18040 26056 18068
rect 26056 18022 26108 18028
rect 25780 17876 25832 17882
rect 25780 17818 25832 17824
rect 25872 16992 25924 16998
rect 25872 16934 25924 16940
rect 25884 16794 25912 16934
rect 25872 16788 25924 16794
rect 25872 16730 25924 16736
rect 25964 16788 26016 16794
rect 25964 16730 26016 16736
rect 25976 16674 26004 16730
rect 25700 16646 26004 16674
rect 25700 16590 25728 16646
rect 25688 16584 25740 16590
rect 25688 16526 25740 16532
rect 25872 16584 25924 16590
rect 25872 16526 25924 16532
rect 25504 16516 25556 16522
rect 25504 16458 25556 16464
rect 25884 16454 25912 16526
rect 25412 16448 25464 16454
rect 25412 16390 25464 16396
rect 25872 16448 25924 16454
rect 25872 16390 25924 16396
rect 25872 16108 25924 16114
rect 25872 16050 25924 16056
rect 25688 15496 25740 15502
rect 25688 15438 25740 15444
rect 25700 15162 25728 15438
rect 25688 15156 25740 15162
rect 25688 15098 25740 15104
rect 25884 15094 25912 16050
rect 26068 15910 26096 18022
rect 26148 17808 26200 17814
rect 26148 17750 26200 17756
rect 26160 15910 26188 17750
rect 26252 17270 26280 19366
rect 26344 18986 26372 19654
rect 26516 19372 26568 19378
rect 26516 19314 26568 19320
rect 26528 19145 26556 19314
rect 26620 19310 26648 19722
rect 26608 19304 26660 19310
rect 26608 19246 26660 19252
rect 26514 19136 26570 19145
rect 26514 19071 26570 19080
rect 26606 19000 26662 19009
rect 26344 18958 26556 18986
rect 26344 18698 26372 18958
rect 26422 18864 26478 18873
rect 26422 18799 26478 18808
rect 26436 18766 26464 18799
rect 26424 18760 26476 18766
rect 26424 18702 26476 18708
rect 26332 18692 26384 18698
rect 26332 18634 26384 18640
rect 26424 18624 26476 18630
rect 26424 18566 26476 18572
rect 26436 17678 26464 18566
rect 26528 18358 26556 18958
rect 26606 18935 26662 18944
rect 26620 18834 26648 18935
rect 26608 18828 26660 18834
rect 26608 18770 26660 18776
rect 26608 18624 26660 18630
rect 26608 18566 26660 18572
rect 26516 18352 26568 18358
rect 26516 18294 26568 18300
rect 26516 18216 26568 18222
rect 26516 18158 26568 18164
rect 26528 17882 26556 18158
rect 26516 17876 26568 17882
rect 26516 17818 26568 17824
rect 26620 17746 26648 18566
rect 26608 17740 26660 17746
rect 26608 17682 26660 17688
rect 26332 17672 26384 17678
rect 26332 17614 26384 17620
rect 26424 17672 26476 17678
rect 26424 17614 26476 17620
rect 26240 17264 26292 17270
rect 26240 17206 26292 17212
rect 26344 17218 26372 17614
rect 26252 16590 26280 17206
rect 26344 17190 26464 17218
rect 26436 17134 26464 17190
rect 26332 17128 26384 17134
rect 26330 17096 26332 17105
rect 26424 17128 26476 17134
rect 26384 17096 26386 17105
rect 26424 17070 26476 17076
rect 26330 17031 26386 17040
rect 26436 16980 26464 17070
rect 26344 16952 26464 16980
rect 26240 16584 26292 16590
rect 26240 16526 26292 16532
rect 26056 15904 26108 15910
rect 26056 15846 26108 15852
rect 26148 15904 26200 15910
rect 26148 15846 26200 15852
rect 25964 15428 26016 15434
rect 25964 15370 26016 15376
rect 25976 15094 26004 15370
rect 26160 15162 26188 15846
rect 26344 15638 26372 16952
rect 26422 16688 26478 16697
rect 26712 16674 26740 20538
rect 26976 20528 27028 20534
rect 26976 20470 27028 20476
rect 26988 19938 27016 20470
rect 27080 20262 27108 23695
rect 27356 23225 27384 25094
rect 27436 24812 27488 24818
rect 27436 24754 27488 24760
rect 27448 24342 27476 24754
rect 27528 24744 27580 24750
rect 27528 24686 27580 24692
rect 27540 24585 27568 24686
rect 27526 24576 27582 24585
rect 27526 24511 27582 24520
rect 27436 24336 27488 24342
rect 27436 24278 27488 24284
rect 27724 23730 27752 25162
rect 28172 25152 28224 25158
rect 28172 25094 28224 25100
rect 27804 24744 27856 24750
rect 27804 24686 27856 24692
rect 27816 24410 27844 24686
rect 27804 24404 27856 24410
rect 27804 24346 27856 24352
rect 28080 24268 28132 24274
rect 28080 24210 28132 24216
rect 27896 24064 27948 24070
rect 27896 24006 27948 24012
rect 27436 23724 27488 23730
rect 27436 23666 27488 23672
rect 27712 23724 27764 23730
rect 27712 23666 27764 23672
rect 27804 23724 27856 23730
rect 27804 23666 27856 23672
rect 27342 23216 27398 23225
rect 27342 23151 27398 23160
rect 27160 20936 27212 20942
rect 27160 20878 27212 20884
rect 27068 20256 27120 20262
rect 27068 20198 27120 20204
rect 27080 20058 27108 20198
rect 27068 20052 27120 20058
rect 27068 19994 27120 20000
rect 26988 19910 27108 19938
rect 26884 19508 26936 19514
rect 26884 19450 26936 19456
rect 26792 18624 26844 18630
rect 26790 18592 26792 18601
rect 26844 18592 26846 18601
rect 26790 18527 26846 18536
rect 26804 17338 26832 18527
rect 26792 17332 26844 17338
rect 26792 17274 26844 17280
rect 26896 16794 26924 19450
rect 26974 19272 27030 19281
rect 26974 19207 27030 19216
rect 26988 19174 27016 19207
rect 26976 19168 27028 19174
rect 26976 19110 27028 19116
rect 26974 19000 27030 19009
rect 26974 18935 26976 18944
rect 27028 18935 27030 18944
rect 26976 18906 27028 18912
rect 26974 18728 27030 18737
rect 26974 18663 27030 18672
rect 26988 18630 27016 18663
rect 26976 18624 27028 18630
rect 26976 18566 27028 18572
rect 26976 18216 27028 18222
rect 26976 18158 27028 18164
rect 26884 16788 26936 16794
rect 26884 16730 26936 16736
rect 26422 16623 26424 16632
rect 26476 16623 26478 16632
rect 26620 16646 26740 16674
rect 26988 16658 27016 18158
rect 26976 16652 27028 16658
rect 26424 16594 26476 16600
rect 26424 16108 26476 16114
rect 26620 16096 26648 16646
rect 26976 16594 27028 16600
rect 26792 16584 26844 16590
rect 26792 16526 26844 16532
rect 26476 16068 26648 16096
rect 26424 16050 26476 16056
rect 26516 15972 26568 15978
rect 26516 15914 26568 15920
rect 26332 15632 26384 15638
rect 26332 15574 26384 15580
rect 26240 15360 26292 15366
rect 26240 15302 26292 15308
rect 26148 15156 26200 15162
rect 26148 15098 26200 15104
rect 25872 15088 25924 15094
rect 25872 15030 25924 15036
rect 25964 15088 26016 15094
rect 25964 15030 26016 15036
rect 25320 14952 25372 14958
rect 25320 14894 25372 14900
rect 25884 14822 25912 15030
rect 25872 14816 25924 14822
rect 25872 14758 25924 14764
rect 25964 14340 26016 14346
rect 25964 14282 26016 14288
rect 25596 14000 25648 14006
rect 25596 13942 25648 13948
rect 24676 13932 24808 13938
rect 24728 13926 24808 13932
rect 24860 13932 24912 13938
rect 24676 13874 24728 13880
rect 24860 13874 24912 13880
rect 24400 12980 24452 12986
rect 24400 12922 24452 12928
rect 24584 12980 24636 12986
rect 24584 12922 24636 12928
rect 24216 12912 24268 12918
rect 24216 12854 24268 12860
rect 24596 12306 24624 12922
rect 24768 12776 24820 12782
rect 24768 12718 24820 12724
rect 24584 12300 24636 12306
rect 24584 12242 24636 12248
rect 22192 12164 22244 12170
rect 22192 12106 22244 12112
rect 20956 12044 21128 12050
rect 20904 12038 21128 12044
rect 20916 12022 21128 12038
rect 21100 11694 21128 12022
rect 22204 11830 22232 12106
rect 24780 12102 24808 12718
rect 24872 12442 24900 13874
rect 25608 12986 25636 13942
rect 25780 13728 25832 13734
rect 25780 13670 25832 13676
rect 25596 12980 25648 12986
rect 25596 12922 25648 12928
rect 25792 12850 25820 13670
rect 25976 12850 26004 14282
rect 26160 14278 26188 15098
rect 26252 14482 26280 15302
rect 26240 14476 26292 14482
rect 26240 14418 26292 14424
rect 26344 14346 26372 15574
rect 26528 15570 26556 15914
rect 26620 15706 26648 16068
rect 26700 16040 26752 16046
rect 26700 15982 26752 15988
rect 26608 15700 26660 15706
rect 26608 15642 26660 15648
rect 26712 15638 26740 15982
rect 26804 15978 26832 16526
rect 26884 16448 26936 16454
rect 26884 16390 26936 16396
rect 26896 16046 26924 16390
rect 26884 16040 26936 16046
rect 26884 15982 26936 15988
rect 26792 15972 26844 15978
rect 26792 15914 26844 15920
rect 26700 15632 26752 15638
rect 26700 15574 26752 15580
rect 26516 15564 26568 15570
rect 26516 15506 26568 15512
rect 26332 14340 26384 14346
rect 26332 14282 26384 14288
rect 26528 14278 26556 15506
rect 26700 15428 26752 15434
rect 26700 15370 26752 15376
rect 26712 14618 26740 15370
rect 26792 14884 26844 14890
rect 26792 14826 26844 14832
rect 26700 14612 26752 14618
rect 26700 14554 26752 14560
rect 26148 14272 26200 14278
rect 26148 14214 26200 14220
rect 26516 14272 26568 14278
rect 26516 14214 26568 14220
rect 26160 12918 26188 14214
rect 26804 13870 26832 14826
rect 26988 14482 27016 16594
rect 27080 14482 27108 19910
rect 27172 14822 27200 20878
rect 27356 20602 27384 23151
rect 27448 22778 27476 23666
rect 27816 23633 27844 23666
rect 27802 23624 27858 23633
rect 27802 23559 27858 23568
rect 27528 23112 27580 23118
rect 27528 23054 27580 23060
rect 27436 22772 27488 22778
rect 27436 22714 27488 22720
rect 27540 22098 27568 23054
rect 27528 22092 27580 22098
rect 27528 22034 27580 22040
rect 27434 21992 27490 22001
rect 27434 21927 27436 21936
rect 27488 21927 27490 21936
rect 27436 21898 27488 21904
rect 27540 21622 27568 22034
rect 27528 21616 27580 21622
rect 27528 21558 27580 21564
rect 27540 21010 27568 21558
rect 27712 21480 27764 21486
rect 27712 21422 27764 21428
rect 27528 21004 27580 21010
rect 27528 20946 27580 20952
rect 27540 20754 27568 20946
rect 27724 20806 27752 21422
rect 27804 20868 27856 20874
rect 27804 20810 27856 20816
rect 27712 20800 27764 20806
rect 27540 20726 27660 20754
rect 27712 20742 27764 20748
rect 27344 20596 27396 20602
rect 27344 20538 27396 20544
rect 27252 19304 27304 19310
rect 27252 19246 27304 19252
rect 27264 19009 27292 19246
rect 27250 19000 27306 19009
rect 27250 18935 27306 18944
rect 27342 18864 27398 18873
rect 27632 18834 27660 20726
rect 27724 20466 27752 20742
rect 27712 20460 27764 20466
rect 27712 20402 27764 20408
rect 27724 19922 27752 20402
rect 27816 20398 27844 20810
rect 27804 20392 27856 20398
rect 27804 20334 27856 20340
rect 27712 19916 27764 19922
rect 27712 19858 27764 19864
rect 27908 19786 27936 24006
rect 28092 23798 28120 24210
rect 28184 24206 28212 25094
rect 28368 24750 28396 25230
rect 28356 24744 28408 24750
rect 28356 24686 28408 24692
rect 28368 24274 28396 24686
rect 28460 24449 28488 25230
rect 28644 25226 28672 25774
rect 28724 25696 28776 25702
rect 28724 25638 28776 25644
rect 28632 25220 28684 25226
rect 28632 25162 28684 25168
rect 28736 25106 28764 25638
rect 28828 25498 28856 26318
rect 28920 25974 28948 27066
rect 29092 26580 29144 26586
rect 29092 26522 29144 26528
rect 28908 25968 28960 25974
rect 28908 25910 28960 25916
rect 28816 25492 28868 25498
rect 28816 25434 28868 25440
rect 28816 25288 28868 25294
rect 28816 25230 28868 25236
rect 28828 25106 28856 25230
rect 28552 25078 28856 25106
rect 28446 24440 28502 24449
rect 28446 24375 28502 24384
rect 28356 24268 28408 24274
rect 28356 24210 28408 24216
rect 28172 24200 28224 24206
rect 28172 24142 28224 24148
rect 28080 23792 28132 23798
rect 28080 23734 28132 23740
rect 28264 23724 28316 23730
rect 28448 23724 28500 23730
rect 28316 23684 28448 23712
rect 28264 23666 28316 23672
rect 28448 23666 28500 23672
rect 27988 23656 28040 23662
rect 27988 23598 28040 23604
rect 28000 22982 28028 23598
rect 28356 23588 28408 23594
rect 28356 23530 28408 23536
rect 28080 23044 28132 23050
rect 28080 22986 28132 22992
rect 27988 22976 28040 22982
rect 27988 22918 28040 22924
rect 28000 22166 28028 22918
rect 28092 22778 28120 22986
rect 28080 22772 28132 22778
rect 28080 22714 28132 22720
rect 28368 22642 28396 23530
rect 28448 23520 28500 23526
rect 28448 23462 28500 23468
rect 28460 23050 28488 23462
rect 28448 23044 28500 23050
rect 28448 22986 28500 22992
rect 28552 22710 28580 25078
rect 28920 24818 28948 25910
rect 28998 25256 29054 25265
rect 28998 25191 29054 25200
rect 28908 24812 28960 24818
rect 28908 24754 28960 24760
rect 28814 24440 28870 24449
rect 28814 24375 28870 24384
rect 28828 24206 28856 24375
rect 28816 24200 28868 24206
rect 28736 24160 28816 24188
rect 28632 23520 28684 23526
rect 28632 23462 28684 23468
rect 28540 22704 28592 22710
rect 28540 22646 28592 22652
rect 28264 22636 28316 22642
rect 28264 22578 28316 22584
rect 28356 22636 28408 22642
rect 28356 22578 28408 22584
rect 28448 22636 28500 22642
rect 28448 22578 28500 22584
rect 28172 22228 28224 22234
rect 28172 22170 28224 22176
rect 27988 22160 28040 22166
rect 27988 22102 28040 22108
rect 27988 21956 28040 21962
rect 27988 21898 28040 21904
rect 28000 21690 28028 21898
rect 27988 21684 28040 21690
rect 27988 21626 28040 21632
rect 27896 19780 27948 19786
rect 27896 19722 27948 19728
rect 28184 19514 28212 22170
rect 28172 19508 28224 19514
rect 28172 19450 28224 19456
rect 28276 19242 28304 22578
rect 28264 19236 28316 19242
rect 28184 19196 28264 19224
rect 27342 18799 27398 18808
rect 27620 18828 27672 18834
rect 27356 18766 27384 18799
rect 27620 18770 27672 18776
rect 27344 18760 27396 18766
rect 27396 18720 27568 18748
rect 27344 18702 27396 18708
rect 27344 18624 27396 18630
rect 27344 18566 27396 18572
rect 27252 16992 27304 16998
rect 27252 16934 27304 16940
rect 27264 16658 27292 16934
rect 27252 16652 27304 16658
rect 27252 16594 27304 16600
rect 27356 16182 27384 18566
rect 27344 16176 27396 16182
rect 27344 16118 27396 16124
rect 27356 15434 27384 16118
rect 27540 16114 27568 18720
rect 27988 18692 28040 18698
rect 27988 18634 28040 18640
rect 28000 18290 28028 18634
rect 28184 18290 28212 19196
rect 28264 19178 28316 19184
rect 28264 18624 28316 18630
rect 28264 18566 28316 18572
rect 28276 18290 28304 18566
rect 27988 18284 28040 18290
rect 27988 18226 28040 18232
rect 28172 18284 28224 18290
rect 28172 18226 28224 18232
rect 28264 18284 28316 18290
rect 28264 18226 28316 18232
rect 27896 17196 27948 17202
rect 27896 17138 27948 17144
rect 27804 17128 27856 17134
rect 27804 17070 27856 17076
rect 27816 16969 27844 17070
rect 27802 16960 27858 16969
rect 27802 16895 27858 16904
rect 27816 16794 27844 16895
rect 27804 16788 27856 16794
rect 27804 16730 27856 16736
rect 27528 16108 27580 16114
rect 27528 16050 27580 16056
rect 27908 15910 27936 17138
rect 28356 16584 28408 16590
rect 28356 16526 28408 16532
rect 27896 15904 27948 15910
rect 27896 15846 27948 15852
rect 27988 15904 28040 15910
rect 27988 15846 28040 15852
rect 28000 15609 28028 15846
rect 27710 15600 27766 15609
rect 27710 15535 27766 15544
rect 27986 15600 28042 15609
rect 27986 15535 28042 15544
rect 27344 15428 27396 15434
rect 27344 15370 27396 15376
rect 27160 14816 27212 14822
rect 27160 14758 27212 14764
rect 26976 14476 27028 14482
rect 26976 14418 27028 14424
rect 27068 14476 27120 14482
rect 27068 14418 27120 14424
rect 26988 14074 27016 14418
rect 27172 14414 27200 14758
rect 27160 14408 27212 14414
rect 27160 14350 27212 14356
rect 26976 14068 27028 14074
rect 26976 14010 27028 14016
rect 26792 13864 26844 13870
rect 26792 13806 26844 13812
rect 26424 13388 26476 13394
rect 26424 13330 26476 13336
rect 26238 13016 26294 13025
rect 26238 12951 26294 12960
rect 26148 12912 26200 12918
rect 26148 12854 26200 12860
rect 25780 12844 25832 12850
rect 25780 12786 25832 12792
rect 25964 12844 26016 12850
rect 25964 12786 26016 12792
rect 24860 12436 24912 12442
rect 24860 12378 24912 12384
rect 26252 12102 26280 12951
rect 26332 12844 26384 12850
rect 26332 12786 26384 12792
rect 26344 12374 26372 12786
rect 26436 12434 26464 13330
rect 26516 13184 26568 13190
rect 26516 13126 26568 13132
rect 26528 12986 26556 13126
rect 26516 12980 26568 12986
rect 26516 12922 26568 12928
rect 26804 12782 26832 13806
rect 27160 13388 27212 13394
rect 27160 13330 27212 13336
rect 26792 12776 26844 12782
rect 26792 12718 26844 12724
rect 26608 12708 26660 12714
rect 26608 12650 26660 12656
rect 26436 12406 26556 12434
rect 26332 12368 26384 12374
rect 26332 12310 26384 12316
rect 24768 12096 24820 12102
rect 24768 12038 24820 12044
rect 26240 12096 26292 12102
rect 26240 12038 26292 12044
rect 22192 11824 22244 11830
rect 22192 11766 22244 11772
rect 21088 11688 21140 11694
rect 21088 11630 21140 11636
rect 22468 11688 22520 11694
rect 22468 11630 22520 11636
rect 20168 11552 20220 11558
rect 20168 11494 20220 11500
rect 22008 11552 22060 11558
rect 22008 11494 22060 11500
rect 20076 11008 20128 11014
rect 20076 10950 20128 10956
rect 19984 10736 20036 10742
rect 19984 10678 20036 10684
rect 19892 10464 19944 10470
rect 19892 10406 19944 10412
rect 19996 10062 20024 10678
rect 20088 10062 20116 10950
rect 20180 10810 20208 11494
rect 21364 11212 21416 11218
rect 21364 11154 21416 11160
rect 20720 11144 20772 11150
rect 20720 11086 20772 11092
rect 20168 10804 20220 10810
rect 20168 10746 20220 10752
rect 20732 10674 20760 11086
rect 21376 10674 21404 11154
rect 22020 11150 22048 11494
rect 22480 11354 22508 11630
rect 22468 11348 22520 11354
rect 22468 11290 22520 11296
rect 22008 11144 22060 11150
rect 22008 11086 22060 11092
rect 22480 10810 22508 11290
rect 22560 11280 22612 11286
rect 22560 11222 22612 11228
rect 22468 10804 22520 10810
rect 22468 10746 22520 10752
rect 22100 10736 22152 10742
rect 22100 10678 22152 10684
rect 20720 10668 20772 10674
rect 20720 10610 20772 10616
rect 21364 10668 21416 10674
rect 21364 10610 21416 10616
rect 20260 10532 20312 10538
rect 20260 10474 20312 10480
rect 20272 10062 20300 10474
rect 19984 10056 20036 10062
rect 19984 9998 20036 10004
rect 20076 10056 20128 10062
rect 20076 9998 20128 10004
rect 20260 10056 20312 10062
rect 20260 9998 20312 10004
rect 19996 8906 20024 9998
rect 21376 9926 21404 10610
rect 22008 10532 22060 10538
rect 22008 10474 22060 10480
rect 21640 10464 21692 10470
rect 21640 10406 21692 10412
rect 21652 10198 21680 10406
rect 22020 10266 22048 10474
rect 22008 10260 22060 10266
rect 22008 10202 22060 10208
rect 21640 10192 21692 10198
rect 21640 10134 21692 10140
rect 22112 9994 22140 10678
rect 22572 10266 22600 11222
rect 24952 11144 25004 11150
rect 24952 11086 25004 11092
rect 22928 11076 22980 11082
rect 22928 11018 22980 11024
rect 22940 10742 22968 11018
rect 22928 10736 22980 10742
rect 22928 10678 22980 10684
rect 22836 10600 22888 10606
rect 22836 10542 22888 10548
rect 22848 10266 22876 10542
rect 22560 10260 22612 10266
rect 22560 10202 22612 10208
rect 22836 10260 22888 10266
rect 22836 10202 22888 10208
rect 22572 10062 22600 10202
rect 22560 10056 22612 10062
rect 22560 9998 22612 10004
rect 22100 9988 22152 9994
rect 22100 9930 22152 9936
rect 21364 9920 21416 9926
rect 21364 9862 21416 9868
rect 22376 9920 22428 9926
rect 22376 9862 22428 9868
rect 21376 9466 21404 9862
rect 21824 9580 21876 9586
rect 21824 9522 21876 9528
rect 21916 9580 21968 9586
rect 21916 9522 21968 9528
rect 21192 9438 21404 9466
rect 21732 9512 21784 9518
rect 21732 9454 21784 9460
rect 21192 9178 21220 9438
rect 21180 9172 21232 9178
rect 21180 9114 21232 9120
rect 21744 9110 21772 9454
rect 21732 9104 21784 9110
rect 21732 9046 21784 9052
rect 21744 8906 21772 9046
rect 21836 8906 21864 9522
rect 21928 9178 21956 9522
rect 21916 9172 21968 9178
rect 21916 9114 21968 9120
rect 22388 9110 22416 9862
rect 22468 9376 22520 9382
rect 22468 9318 22520 9324
rect 22376 9104 22428 9110
rect 22376 9046 22428 9052
rect 19984 8900 20036 8906
rect 19984 8842 20036 8848
rect 21548 8900 21600 8906
rect 21548 8842 21600 8848
rect 21732 8900 21784 8906
rect 21732 8842 21784 8848
rect 21824 8900 21876 8906
rect 21824 8842 21876 8848
rect 20720 8832 20772 8838
rect 20720 8774 20772 8780
rect 21088 8832 21140 8838
rect 21088 8774 21140 8780
rect 21364 8832 21416 8838
rect 21364 8774 21416 8780
rect 20732 8498 20760 8774
rect 20720 8492 20772 8498
rect 20720 8434 20772 8440
rect 19432 8424 19484 8430
rect 19432 8366 19484 8372
rect 19444 8090 19472 8366
rect 19432 8084 19484 8090
rect 19432 8026 19484 8032
rect 21100 7954 21128 8774
rect 21180 8628 21232 8634
rect 21180 8570 21232 8576
rect 21088 7948 21140 7954
rect 21088 7890 21140 7896
rect 21100 7546 21128 7890
rect 21192 7818 21220 8570
rect 21376 8294 21404 8774
rect 21560 8498 21588 8842
rect 21732 8560 21784 8566
rect 21732 8502 21784 8508
rect 21548 8492 21600 8498
rect 21548 8434 21600 8440
rect 21364 8288 21416 8294
rect 21364 8230 21416 8236
rect 21560 7954 21588 8434
rect 21744 8090 21772 8502
rect 21836 8430 21864 8842
rect 22480 8498 22508 9318
rect 22940 8566 22968 10678
rect 24964 10606 24992 11086
rect 26528 10674 26556 12406
rect 26620 12238 26648 12650
rect 26792 12436 26844 12442
rect 26792 12378 26844 12384
rect 26700 12300 26752 12306
rect 26700 12242 26752 12248
rect 26608 12232 26660 12238
rect 26608 12174 26660 12180
rect 26712 11898 26740 12242
rect 26804 11914 26832 12378
rect 26884 12368 26936 12374
rect 26884 12310 26936 12316
rect 26896 12102 26924 12310
rect 27172 12238 27200 13330
rect 27618 13016 27674 13025
rect 27618 12951 27620 12960
rect 27672 12951 27674 12960
rect 27620 12922 27672 12928
rect 27252 12640 27304 12646
rect 27252 12582 27304 12588
rect 27160 12232 27212 12238
rect 27160 12174 27212 12180
rect 26884 12096 26936 12102
rect 26884 12038 26936 12044
rect 26976 12096 27028 12102
rect 26976 12038 27028 12044
rect 26988 11914 27016 12038
rect 26700 11892 26752 11898
rect 26700 11834 26752 11840
rect 26804 11886 27016 11914
rect 27264 11898 27292 12582
rect 27344 12300 27396 12306
rect 27344 12242 27396 12248
rect 27252 11892 27304 11898
rect 26700 11756 26752 11762
rect 26700 11698 26752 11704
rect 26712 11121 26740 11698
rect 26698 11112 26754 11121
rect 26698 11047 26754 11056
rect 26712 10810 26740 11047
rect 26700 10804 26752 10810
rect 26700 10746 26752 10752
rect 26608 10736 26660 10742
rect 26608 10678 26660 10684
rect 26516 10668 26568 10674
rect 26516 10610 26568 10616
rect 23940 10600 23992 10606
rect 23940 10542 23992 10548
rect 24952 10600 25004 10606
rect 24952 10542 25004 10548
rect 25872 10600 25924 10606
rect 25872 10542 25924 10548
rect 23112 10124 23164 10130
rect 23112 10066 23164 10072
rect 23020 10056 23072 10062
rect 23020 9998 23072 10004
rect 23032 9450 23060 9998
rect 23020 9444 23072 9450
rect 23020 9386 23072 9392
rect 22928 8560 22980 8566
rect 22928 8502 22980 8508
rect 22468 8492 22520 8498
rect 22468 8434 22520 8440
rect 21824 8424 21876 8430
rect 21824 8366 21876 8372
rect 21836 8090 21864 8366
rect 22940 8362 22968 8502
rect 22928 8356 22980 8362
rect 22928 8298 22980 8304
rect 21732 8084 21784 8090
rect 21732 8026 21784 8032
rect 21824 8084 21876 8090
rect 21824 8026 21876 8032
rect 21548 7948 21600 7954
rect 21548 7890 21600 7896
rect 21180 7812 21232 7818
rect 21180 7754 21232 7760
rect 21364 7744 21416 7750
rect 21364 7686 21416 7692
rect 21088 7540 21140 7546
rect 21088 7482 21140 7488
rect 21376 7410 21404 7686
rect 20352 7404 20404 7410
rect 20352 7346 20404 7352
rect 20444 7404 20496 7410
rect 20444 7346 20496 7352
rect 20536 7404 20588 7410
rect 20536 7346 20588 7352
rect 21364 7404 21416 7410
rect 21364 7346 21416 7352
rect 20260 7336 20312 7342
rect 20260 7278 20312 7284
rect 20272 6798 20300 7278
rect 20260 6792 20312 6798
rect 20260 6734 20312 6740
rect 20364 6730 20392 7346
rect 20352 6724 20404 6730
rect 20352 6666 20404 6672
rect 20456 6458 20484 7346
rect 20548 6798 20576 7346
rect 20720 7268 20772 7274
rect 20720 7210 20772 7216
rect 20732 6866 20760 7210
rect 21272 7200 21324 7206
rect 21272 7142 21324 7148
rect 20720 6860 20772 6866
rect 20720 6802 20772 6808
rect 20536 6792 20588 6798
rect 20536 6734 20588 6740
rect 20444 6452 20496 6458
rect 20444 6394 20496 6400
rect 19984 6384 20036 6390
rect 19984 6326 20036 6332
rect 19708 6180 19760 6186
rect 19708 6122 19760 6128
rect 19720 5794 19748 6122
rect 19628 5778 19748 5794
rect 19996 5778 20024 6326
rect 20548 5914 20576 6734
rect 20628 6656 20680 6662
rect 20628 6598 20680 6604
rect 20640 6390 20668 6598
rect 20732 6458 20760 6802
rect 20812 6792 20864 6798
rect 20812 6734 20864 6740
rect 20720 6452 20772 6458
rect 20720 6394 20772 6400
rect 20628 6384 20680 6390
rect 20628 6326 20680 6332
rect 20628 6248 20680 6254
rect 20732 6236 20760 6394
rect 20824 6322 20852 6734
rect 20904 6656 20956 6662
rect 20904 6598 20956 6604
rect 20812 6316 20864 6322
rect 20812 6258 20864 6264
rect 20680 6208 20760 6236
rect 20628 6190 20680 6196
rect 20916 6186 20944 6598
rect 20996 6384 21048 6390
rect 20996 6326 21048 6332
rect 20904 6180 20956 6186
rect 20904 6122 20956 6128
rect 20536 5908 20588 5914
rect 20536 5850 20588 5856
rect 19616 5772 19748 5778
rect 19668 5766 19748 5772
rect 19616 5714 19668 5720
rect 19432 5636 19484 5642
rect 19432 5578 19484 5584
rect 19444 5370 19472 5578
rect 19432 5364 19484 5370
rect 19432 5306 19484 5312
rect 19720 4078 19748 5766
rect 19984 5772 20036 5778
rect 19984 5714 20036 5720
rect 19996 5642 20024 5714
rect 19984 5636 20036 5642
rect 19984 5578 20036 5584
rect 20548 5234 20576 5850
rect 21008 5778 21036 6326
rect 21088 6112 21140 6118
rect 21088 6054 21140 6060
rect 21100 5778 21128 6054
rect 20720 5772 20772 5778
rect 20720 5714 20772 5720
rect 20996 5772 21048 5778
rect 20996 5714 21048 5720
rect 21088 5772 21140 5778
rect 21088 5714 21140 5720
rect 20536 5228 20588 5234
rect 20536 5170 20588 5176
rect 19984 4480 20036 4486
rect 19984 4422 20036 4428
rect 19996 4214 20024 4422
rect 20732 4214 20760 5714
rect 21284 5710 21312 7142
rect 21376 6866 21404 7346
rect 21364 6860 21416 6866
rect 21364 6802 21416 6808
rect 21744 6798 21772 8026
rect 22008 7336 22060 7342
rect 22008 7278 22060 7284
rect 22020 6798 22048 7278
rect 22940 6866 22968 8298
rect 23124 7410 23152 10066
rect 23664 9920 23716 9926
rect 23664 9862 23716 9868
rect 23296 9716 23348 9722
rect 23296 9658 23348 9664
rect 23308 7546 23336 9658
rect 23480 9512 23532 9518
rect 23480 9454 23532 9460
rect 23492 8634 23520 9454
rect 23676 9042 23704 9862
rect 23664 9036 23716 9042
rect 23664 8978 23716 8984
rect 23952 8974 23980 10542
rect 25884 10266 25912 10542
rect 25872 10260 25924 10266
rect 25872 10202 25924 10208
rect 23940 8968 23992 8974
rect 23940 8910 23992 8916
rect 23480 8628 23532 8634
rect 23480 8570 23532 8576
rect 23952 8294 23980 8910
rect 26620 8566 26648 10678
rect 26608 8560 26660 8566
rect 26608 8502 26660 8508
rect 25320 8424 25372 8430
rect 25320 8366 25372 8372
rect 23940 8288 23992 8294
rect 23940 8230 23992 8236
rect 23296 7540 23348 7546
rect 23296 7482 23348 7488
rect 23020 7404 23072 7410
rect 23020 7346 23072 7352
rect 23112 7404 23164 7410
rect 23112 7346 23164 7352
rect 22928 6860 22980 6866
rect 22928 6802 22980 6808
rect 21732 6792 21784 6798
rect 21732 6734 21784 6740
rect 22008 6792 22060 6798
rect 22008 6734 22060 6740
rect 21916 6724 21968 6730
rect 21916 6666 21968 6672
rect 21364 6452 21416 6458
rect 21364 6394 21416 6400
rect 21376 6254 21404 6394
rect 21928 6390 21956 6666
rect 21916 6384 21968 6390
rect 21916 6326 21968 6332
rect 21364 6248 21416 6254
rect 21364 6190 21416 6196
rect 21364 6112 21416 6118
rect 21364 6054 21416 6060
rect 21376 5914 21404 6054
rect 21364 5908 21416 5914
rect 21364 5850 21416 5856
rect 21272 5704 21324 5710
rect 21272 5646 21324 5652
rect 21916 4684 21968 4690
rect 21916 4626 21968 4632
rect 21180 4480 21232 4486
rect 21180 4422 21232 4428
rect 19984 4208 20036 4214
rect 19984 4150 20036 4156
rect 20720 4208 20772 4214
rect 20720 4150 20772 4156
rect 19708 4072 19760 4078
rect 19708 4014 19760 4020
rect 19720 3602 19748 4014
rect 19708 3596 19760 3602
rect 19708 3538 19760 3544
rect 20732 3466 20760 4150
rect 19984 3460 20036 3466
rect 19984 3402 20036 3408
rect 20720 3460 20772 3466
rect 20720 3402 20772 3408
rect 19996 3194 20024 3402
rect 19984 3188 20036 3194
rect 19984 3130 20036 3136
rect 21192 2990 21220 4422
rect 21928 4078 21956 4626
rect 21364 4072 21416 4078
rect 21364 4014 21416 4020
rect 21916 4072 21968 4078
rect 21916 4014 21968 4020
rect 21376 3942 21404 4014
rect 22020 4010 22048 6734
rect 22940 6730 22968 6802
rect 22928 6724 22980 6730
rect 22928 6666 22980 6672
rect 23032 6662 23060 7346
rect 23124 7274 23152 7346
rect 23952 7342 23980 8230
rect 25332 8090 25360 8366
rect 25320 8084 25372 8090
rect 25320 8026 25372 8032
rect 26148 7744 26200 7750
rect 26148 7686 26200 7692
rect 23940 7336 23992 7342
rect 23940 7278 23992 7284
rect 23112 7268 23164 7274
rect 23112 7210 23164 7216
rect 23020 6656 23072 6662
rect 23020 6598 23072 6604
rect 22928 4548 22980 4554
rect 22928 4490 22980 4496
rect 22940 4146 22968 4490
rect 23124 4146 23152 7210
rect 23848 7200 23900 7206
rect 23848 7142 23900 7148
rect 25964 7200 26016 7206
rect 25964 7142 26016 7148
rect 23860 7002 23888 7142
rect 25976 7002 26004 7142
rect 23848 6996 23900 7002
rect 23848 6938 23900 6944
rect 25964 6996 26016 7002
rect 25964 6938 26016 6944
rect 23572 6860 23624 6866
rect 23572 6802 23624 6808
rect 23584 6254 23612 6802
rect 26056 6724 26108 6730
rect 26056 6666 26108 6672
rect 23296 6248 23348 6254
rect 23296 6190 23348 6196
rect 23572 6248 23624 6254
rect 23572 6190 23624 6196
rect 23308 5914 23336 6190
rect 23296 5908 23348 5914
rect 23296 5850 23348 5856
rect 23584 5302 23612 6190
rect 24768 5704 24820 5710
rect 24768 5646 24820 5652
rect 24780 5370 24808 5646
rect 24768 5364 24820 5370
rect 24768 5306 24820 5312
rect 23572 5296 23624 5302
rect 23572 5238 23624 5244
rect 23940 5160 23992 5166
rect 23940 5102 23992 5108
rect 23952 4826 23980 5102
rect 23940 4820 23992 4826
rect 23940 4762 23992 4768
rect 24780 4690 24808 5306
rect 26068 5302 26096 6666
rect 26056 5296 26108 5302
rect 26056 5238 26108 5244
rect 24768 4684 24820 4690
rect 24768 4626 24820 4632
rect 23388 4548 23440 4554
rect 23388 4490 23440 4496
rect 24676 4548 24728 4554
rect 24676 4490 24728 4496
rect 23204 4480 23256 4486
rect 23204 4422 23256 4428
rect 23216 4282 23244 4422
rect 23204 4276 23256 4282
rect 23204 4218 23256 4224
rect 22560 4140 22612 4146
rect 22560 4082 22612 4088
rect 22928 4140 22980 4146
rect 22928 4082 22980 4088
rect 23112 4140 23164 4146
rect 23112 4082 23164 4088
rect 22008 4004 22060 4010
rect 22008 3946 22060 3952
rect 21364 3936 21416 3942
rect 21364 3878 21416 3884
rect 21548 3936 21600 3942
rect 21548 3878 21600 3884
rect 21180 2984 21232 2990
rect 21180 2926 21232 2932
rect 19340 2644 19392 2650
rect 19340 2586 19392 2592
rect 21376 2378 21404 3878
rect 21560 2990 21588 3878
rect 21824 3460 21876 3466
rect 21824 3402 21876 3408
rect 21836 2990 21864 3402
rect 21916 3392 21968 3398
rect 21916 3334 21968 3340
rect 21928 3058 21956 3334
rect 22572 3194 22600 4082
rect 22836 3936 22888 3942
rect 22836 3878 22888 3884
rect 22652 3392 22704 3398
rect 22652 3334 22704 3340
rect 22192 3188 22244 3194
rect 22192 3130 22244 3136
rect 22560 3188 22612 3194
rect 22560 3130 22612 3136
rect 21916 3052 21968 3058
rect 21916 2994 21968 3000
rect 21548 2984 21600 2990
rect 21548 2926 21600 2932
rect 21824 2984 21876 2990
rect 21824 2926 21876 2932
rect 21836 2514 21864 2926
rect 22204 2922 22232 3130
rect 22664 3126 22692 3334
rect 22848 3126 22876 3878
rect 22940 3466 22968 4082
rect 23400 4078 23428 4490
rect 23480 4208 23532 4214
rect 23480 4150 23532 4156
rect 23388 4072 23440 4078
rect 23388 4014 23440 4020
rect 23296 3936 23348 3942
rect 23296 3878 23348 3884
rect 22928 3460 22980 3466
rect 22928 3402 22980 3408
rect 22652 3120 22704 3126
rect 22652 3062 22704 3068
rect 22836 3120 22888 3126
rect 22836 3062 22888 3068
rect 22192 2916 22244 2922
rect 22192 2858 22244 2864
rect 21824 2508 21876 2514
rect 21824 2450 21876 2456
rect 22204 2446 22232 2858
rect 22560 2576 22612 2582
rect 22560 2518 22612 2524
rect 22192 2440 22244 2446
rect 22192 2382 22244 2388
rect 21364 2372 21416 2378
rect 21364 2314 21416 2320
rect 19340 2304 19392 2310
rect 19340 2246 19392 2252
rect 20628 2304 20680 2310
rect 20628 2246 20680 2252
rect 21272 2304 21324 2310
rect 21272 2246 21324 2252
rect 4874 2204 5182 2213
rect 4874 2202 4880 2204
rect 4936 2202 4960 2204
rect 5016 2202 5040 2204
rect 5096 2202 5120 2204
rect 5176 2202 5182 2204
rect 4936 2150 4938 2202
rect 5118 2150 5120 2202
rect 4874 2148 4880 2150
rect 4936 2148 4960 2150
rect 5016 2148 5040 2150
rect 5096 2148 5120 2150
rect 5176 2148 5182 2150
rect 4874 2139 5182 2148
rect 19352 800 19380 2246
rect 20640 800 20668 2246
rect 21284 800 21312 2246
rect 22572 800 22600 2518
rect 22664 2378 22692 3062
rect 22940 2990 22968 3402
rect 23308 3398 23336 3878
rect 23400 3534 23428 4014
rect 23492 3670 23520 4150
rect 23756 4072 23808 4078
rect 23756 4014 23808 4020
rect 23480 3664 23532 3670
rect 23480 3606 23532 3612
rect 23388 3528 23440 3534
rect 23388 3470 23440 3476
rect 23296 3392 23348 3398
rect 23296 3334 23348 3340
rect 23388 3392 23440 3398
rect 23388 3334 23440 3340
rect 23308 3194 23336 3334
rect 23296 3188 23348 3194
rect 23296 3130 23348 3136
rect 22928 2984 22980 2990
rect 22928 2926 22980 2932
rect 23296 2984 23348 2990
rect 23296 2926 23348 2932
rect 23308 2514 23336 2926
rect 23400 2922 23428 3334
rect 23768 3194 23796 4014
rect 24688 3738 24716 4490
rect 24676 3732 24728 3738
rect 24676 3674 24728 3680
rect 24780 3602 24808 4626
rect 26068 4554 26096 5238
rect 26160 4826 26188 7686
rect 26620 7342 26648 8502
rect 26804 7954 26832 11886
rect 27252 11834 27304 11840
rect 27252 10668 27304 10674
rect 27252 10610 27304 10616
rect 27264 10470 27292 10610
rect 27252 10464 27304 10470
rect 27252 10406 27304 10412
rect 27356 10062 27384 12242
rect 27620 12096 27672 12102
rect 27620 12038 27672 12044
rect 27632 11558 27660 12038
rect 27620 11552 27672 11558
rect 27620 11494 27672 11500
rect 27632 11082 27660 11494
rect 27620 11076 27672 11082
rect 27620 11018 27672 11024
rect 27632 10198 27660 11018
rect 27724 10266 27752 15535
rect 28368 14618 28396 16526
rect 28356 14612 28408 14618
rect 28356 14554 28408 14560
rect 28368 14346 28396 14554
rect 28356 14340 28408 14346
rect 28356 14282 28408 14288
rect 28368 14006 28396 14282
rect 28356 14000 28408 14006
rect 28356 13942 28408 13948
rect 27988 13456 28040 13462
rect 27988 13398 28040 13404
rect 28000 13326 28028 13398
rect 27988 13320 28040 13326
rect 27988 13262 28040 13268
rect 28000 12442 28028 13262
rect 27988 12436 28040 12442
rect 27988 12378 28040 12384
rect 28356 11756 28408 11762
rect 28356 11698 28408 11704
rect 27988 11552 28040 11558
rect 27988 11494 28040 11500
rect 27896 11076 27948 11082
rect 27896 11018 27948 11024
rect 27908 10810 27936 11018
rect 27896 10804 27948 10810
rect 27896 10746 27948 10752
rect 28000 10674 28028 11494
rect 28368 11150 28396 11698
rect 28356 11144 28408 11150
rect 28356 11086 28408 11092
rect 28368 10674 28396 11086
rect 28460 10810 28488 22578
rect 28644 22094 28672 23462
rect 28552 22066 28672 22094
rect 28552 22030 28580 22066
rect 28540 22024 28592 22030
rect 28540 21966 28592 21972
rect 28644 21622 28672 22066
rect 28736 21894 28764 24160
rect 28816 24142 28868 24148
rect 28920 23712 28948 24754
rect 29012 24614 29040 25191
rect 29000 24608 29052 24614
rect 29000 24550 29052 24556
rect 29104 24206 29132 26522
rect 29196 24449 29224 34886
rect 30392 34678 30420 35022
rect 30380 34672 30432 34678
rect 30380 34614 30432 34620
rect 30288 34060 30340 34066
rect 30288 34002 30340 34008
rect 29368 32292 29420 32298
rect 29368 32234 29420 32240
rect 29380 31822 29408 32234
rect 29920 32224 29972 32230
rect 29920 32166 29972 32172
rect 30104 32224 30156 32230
rect 30104 32166 30156 32172
rect 29932 32026 29960 32166
rect 29920 32020 29972 32026
rect 29920 31962 29972 31968
rect 29368 31816 29420 31822
rect 29368 31758 29420 31764
rect 30116 31754 30144 32166
rect 30300 31754 30328 34002
rect 30392 33590 30420 34614
rect 30472 34536 30524 34542
rect 30472 34478 30524 34484
rect 30484 34202 30512 34478
rect 30472 34196 30524 34202
rect 30472 34138 30524 34144
rect 30668 34134 30696 35022
rect 31208 34944 31260 34950
rect 31208 34886 31260 34892
rect 30656 34128 30708 34134
rect 30656 34070 30708 34076
rect 31116 34128 31168 34134
rect 31116 34070 31168 34076
rect 31128 33998 31156 34070
rect 31220 34066 31248 34886
rect 31864 34202 31892 35022
rect 32312 34536 32364 34542
rect 32312 34478 32364 34484
rect 33232 34536 33284 34542
rect 33232 34478 33284 34484
rect 32128 34400 32180 34406
rect 32128 34342 32180 34348
rect 31852 34196 31904 34202
rect 31852 34138 31904 34144
rect 31208 34060 31260 34066
rect 31208 34002 31260 34008
rect 32036 34060 32088 34066
rect 32036 34002 32088 34008
rect 30656 33992 30708 33998
rect 30656 33934 30708 33940
rect 31116 33992 31168 33998
rect 31116 33934 31168 33940
rect 30380 33584 30432 33590
rect 30380 33526 30432 33532
rect 30104 31748 30156 31754
rect 30104 31690 30156 31696
rect 30208 31726 30328 31754
rect 29368 31680 29420 31686
rect 29368 31622 29420 31628
rect 29380 31278 29408 31622
rect 29552 31476 29604 31482
rect 29552 31418 29604 31424
rect 29368 31272 29420 31278
rect 29368 31214 29420 31220
rect 29276 29640 29328 29646
rect 29276 29582 29328 29588
rect 29288 28558 29316 29582
rect 29276 28552 29328 28558
rect 29276 28494 29328 28500
rect 29564 27402 29592 31418
rect 30116 30938 30144 31690
rect 30208 31482 30236 31726
rect 30196 31476 30248 31482
rect 30196 31418 30248 31424
rect 30392 31346 30420 33526
rect 30668 33386 30696 33934
rect 31668 33924 31720 33930
rect 31668 33866 31720 33872
rect 31116 33516 31168 33522
rect 31116 33458 31168 33464
rect 30656 33380 30708 33386
rect 30656 33322 30708 33328
rect 30564 33312 30616 33318
rect 30564 33254 30616 33260
rect 30576 32910 30604 33254
rect 30668 32910 30696 33322
rect 31128 33114 31156 33458
rect 31680 33454 31708 33866
rect 32048 33658 32076 34002
rect 32140 33998 32168 34342
rect 32128 33992 32180 33998
rect 32128 33934 32180 33940
rect 32036 33652 32088 33658
rect 32036 33594 32088 33600
rect 31668 33448 31720 33454
rect 31668 33390 31720 33396
rect 31116 33108 31168 33114
rect 31116 33050 31168 33056
rect 30564 32904 30616 32910
rect 30564 32846 30616 32852
rect 30656 32904 30708 32910
rect 30656 32846 30708 32852
rect 30840 32768 30892 32774
rect 30840 32710 30892 32716
rect 30472 32564 30524 32570
rect 30472 32506 30524 32512
rect 30484 32434 30512 32506
rect 30852 32502 30880 32710
rect 30840 32496 30892 32502
rect 30840 32438 30892 32444
rect 30472 32428 30524 32434
rect 30472 32370 30524 32376
rect 30564 32428 30616 32434
rect 30564 32370 30616 32376
rect 30380 31340 30432 31346
rect 30380 31282 30432 31288
rect 30104 30932 30156 30938
rect 30104 30874 30156 30880
rect 30484 30734 30512 32370
rect 30576 31686 30604 32370
rect 31300 32360 31352 32366
rect 31300 32302 31352 32308
rect 31312 32026 31340 32302
rect 31300 32020 31352 32026
rect 31300 31962 31352 31968
rect 32324 31822 32352 34478
rect 33244 34202 33272 34478
rect 32680 34196 32732 34202
rect 32680 34138 32732 34144
rect 33232 34196 33284 34202
rect 33232 34138 33284 34144
rect 32692 33998 32720 34138
rect 33048 34060 33100 34066
rect 33048 34002 33100 34008
rect 32680 33992 32732 33998
rect 32680 33934 32732 33940
rect 32772 33992 32824 33998
rect 32772 33934 32824 33940
rect 32784 33862 32812 33934
rect 32772 33856 32824 33862
rect 32772 33798 32824 33804
rect 32784 33046 32812 33798
rect 32956 33516 33008 33522
rect 32956 33458 33008 33464
rect 32772 33040 32824 33046
rect 32772 32982 32824 32988
rect 32784 32910 32812 32982
rect 32772 32904 32824 32910
rect 32772 32846 32824 32852
rect 32588 32836 32640 32842
rect 32588 32778 32640 32784
rect 32312 31816 32364 31822
rect 32312 31758 32364 31764
rect 31576 31748 31628 31754
rect 31576 31690 31628 31696
rect 30564 31680 30616 31686
rect 30564 31622 30616 31628
rect 30576 31142 30604 31622
rect 31588 31346 31616 31690
rect 32324 31414 32352 31758
rect 32036 31408 32088 31414
rect 32036 31350 32088 31356
rect 32312 31408 32364 31414
rect 32312 31350 32364 31356
rect 31576 31340 31628 31346
rect 31576 31282 31628 31288
rect 30564 31136 30616 31142
rect 30564 31078 30616 31084
rect 30576 30734 30604 31078
rect 30472 30728 30524 30734
rect 30472 30670 30524 30676
rect 30564 30728 30616 30734
rect 30564 30670 30616 30676
rect 31588 30666 31616 31282
rect 32048 30802 32076 31350
rect 32036 30796 32088 30802
rect 32036 30738 32088 30744
rect 31576 30660 31628 30666
rect 31576 30602 31628 30608
rect 29644 30048 29696 30054
rect 29644 29990 29696 29996
rect 29656 29714 29684 29990
rect 29644 29708 29696 29714
rect 29644 29650 29696 29656
rect 30012 29640 30064 29646
rect 30012 29582 30064 29588
rect 30024 28422 30052 29582
rect 30472 29572 30524 29578
rect 30472 29514 30524 29520
rect 30484 29306 30512 29514
rect 30472 29300 30524 29306
rect 30472 29242 30524 29248
rect 30484 28558 30512 29242
rect 31588 29238 31616 30602
rect 31576 29232 31628 29238
rect 31576 29174 31628 29180
rect 32048 29170 32076 30738
rect 32220 30592 32272 30598
rect 32220 30534 32272 30540
rect 32232 30394 32260 30534
rect 32220 30388 32272 30394
rect 32220 30330 32272 30336
rect 32600 30326 32628 32778
rect 32968 32502 32996 33458
rect 33060 33318 33088 34002
rect 33140 33924 33192 33930
rect 33140 33866 33192 33872
rect 33048 33312 33100 33318
rect 33048 33254 33100 33260
rect 33152 33114 33180 33866
rect 33140 33108 33192 33114
rect 33140 33050 33192 33056
rect 33046 32600 33102 32609
rect 33046 32535 33102 32544
rect 32956 32496 33008 32502
rect 32956 32438 33008 32444
rect 32864 32428 32916 32434
rect 32864 32370 32916 32376
rect 32876 31686 32904 32370
rect 32968 31822 32996 32438
rect 33060 32298 33088 32535
rect 33336 32337 33364 35974
rect 35594 35932 35902 35941
rect 35594 35930 35600 35932
rect 35656 35930 35680 35932
rect 35736 35930 35760 35932
rect 35816 35930 35840 35932
rect 35896 35930 35902 35932
rect 35656 35878 35658 35930
rect 35838 35878 35840 35930
rect 35594 35876 35600 35878
rect 35656 35876 35680 35878
rect 35736 35876 35760 35878
rect 35816 35876 35840 35878
rect 35896 35876 35902 35878
rect 35594 35867 35902 35876
rect 34934 35388 35242 35397
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35323 35242 35332
rect 35594 34844 35902 34853
rect 35594 34842 35600 34844
rect 35656 34842 35680 34844
rect 35736 34842 35760 34844
rect 35816 34842 35840 34844
rect 35896 34842 35902 34844
rect 35656 34790 35658 34842
rect 35838 34790 35840 34842
rect 35594 34788 35600 34790
rect 35656 34788 35680 34790
rect 35736 34788 35760 34790
rect 35816 34788 35840 34790
rect 35896 34788 35902 34790
rect 35594 34779 35902 34788
rect 34428 34536 34480 34542
rect 34428 34478 34480 34484
rect 33784 34128 33836 34134
rect 33784 34070 33836 34076
rect 33416 33992 33468 33998
rect 33416 33934 33468 33940
rect 33428 33658 33456 33934
rect 33796 33930 33824 34070
rect 34440 34066 34468 34478
rect 34934 34300 35242 34309
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34235 35242 34244
rect 34428 34060 34480 34066
rect 34428 34002 34480 34008
rect 33784 33924 33836 33930
rect 33784 33866 33836 33872
rect 33416 33652 33468 33658
rect 33416 33594 33468 33600
rect 33692 33448 33744 33454
rect 33796 33436 33824 33866
rect 37096 33856 37148 33862
rect 37096 33798 37148 33804
rect 35594 33756 35902 33765
rect 35594 33754 35600 33756
rect 35656 33754 35680 33756
rect 35736 33754 35760 33756
rect 35816 33754 35840 33756
rect 35896 33754 35902 33756
rect 35656 33702 35658 33754
rect 35838 33702 35840 33754
rect 35594 33700 35600 33702
rect 35656 33700 35680 33702
rect 35736 33700 35760 33702
rect 35816 33700 35840 33702
rect 35896 33700 35902 33702
rect 35594 33691 35902 33700
rect 33744 33408 33824 33436
rect 33692 33390 33744 33396
rect 33796 33318 33824 33408
rect 36636 33380 36688 33386
rect 36636 33322 36688 33328
rect 33416 33312 33468 33318
rect 33416 33254 33468 33260
rect 33784 33312 33836 33318
rect 33784 33254 33836 33260
rect 34060 33312 34112 33318
rect 34060 33254 34112 33260
rect 33322 32328 33378 32337
rect 33048 32292 33100 32298
rect 33322 32263 33378 32272
rect 33048 32234 33100 32240
rect 33324 32224 33376 32230
rect 33324 32166 33376 32172
rect 32956 31816 33008 31822
rect 32956 31758 33008 31764
rect 33232 31816 33284 31822
rect 33232 31758 33284 31764
rect 32864 31680 32916 31686
rect 32864 31622 32916 31628
rect 32968 31142 32996 31758
rect 33244 31346 33272 31758
rect 33336 31754 33364 32166
rect 33428 31822 33456 33254
rect 33796 32910 33824 33254
rect 33968 33108 34020 33114
rect 33968 33050 34020 33056
rect 33508 32904 33560 32910
rect 33508 32846 33560 32852
rect 33600 32904 33652 32910
rect 33600 32846 33652 32852
rect 33784 32904 33836 32910
rect 33784 32846 33836 32852
rect 33520 32609 33548 32846
rect 33506 32600 33562 32609
rect 33506 32535 33562 32544
rect 33612 32484 33640 32846
rect 33692 32768 33744 32774
rect 33692 32710 33744 32716
rect 33520 32456 33640 32484
rect 33520 31958 33548 32456
rect 33598 32328 33654 32337
rect 33598 32263 33654 32272
rect 33612 32230 33640 32263
rect 33600 32224 33652 32230
rect 33600 32166 33652 32172
rect 33508 31952 33560 31958
rect 33508 31894 33560 31900
rect 33600 31952 33652 31958
rect 33600 31894 33652 31900
rect 33416 31816 33468 31822
rect 33416 31758 33468 31764
rect 33324 31748 33376 31754
rect 33324 31690 33376 31696
rect 33508 31680 33560 31686
rect 33508 31622 33560 31628
rect 33232 31340 33284 31346
rect 33232 31282 33284 31288
rect 32956 31136 33008 31142
rect 32956 31078 33008 31084
rect 33520 30802 33548 31622
rect 33612 31346 33640 31894
rect 33704 31686 33732 32710
rect 33784 32496 33836 32502
rect 33784 32438 33836 32444
rect 33796 32026 33824 32438
rect 33980 32314 34008 33050
rect 33888 32286 34008 32314
rect 33888 32230 33916 32286
rect 33876 32224 33928 32230
rect 33876 32166 33928 32172
rect 33784 32020 33836 32026
rect 33784 31962 33836 31968
rect 33876 31816 33928 31822
rect 33876 31758 33928 31764
rect 33968 31816 34020 31822
rect 33968 31758 34020 31764
rect 33692 31680 33744 31686
rect 33692 31622 33744 31628
rect 33600 31340 33652 31346
rect 33600 31282 33652 31288
rect 33508 30796 33560 30802
rect 33508 30738 33560 30744
rect 32772 30728 32824 30734
rect 32772 30670 32824 30676
rect 32588 30320 32640 30326
rect 32588 30262 32640 30268
rect 32128 29844 32180 29850
rect 32128 29786 32180 29792
rect 32036 29164 32088 29170
rect 32036 29106 32088 29112
rect 30656 28960 30708 28966
rect 30656 28902 30708 28908
rect 31852 28960 31904 28966
rect 31852 28902 31904 28908
rect 30668 28762 30696 28902
rect 31864 28762 31892 28902
rect 30656 28756 30708 28762
rect 30656 28698 30708 28704
rect 31852 28756 31904 28762
rect 31852 28698 31904 28704
rect 30472 28552 30524 28558
rect 30472 28494 30524 28500
rect 32140 28490 32168 29786
rect 32496 29776 32548 29782
rect 32496 29718 32548 29724
rect 32508 29578 32536 29718
rect 32496 29572 32548 29578
rect 32496 29514 32548 29520
rect 32508 29238 32536 29514
rect 32784 29510 32812 30670
rect 33232 30592 33284 30598
rect 33232 30534 33284 30540
rect 32956 29844 33008 29850
rect 32956 29786 33008 29792
rect 32968 29578 32996 29786
rect 33244 29782 33272 30534
rect 33612 30394 33640 31282
rect 33888 30938 33916 31758
rect 33980 31346 34008 31758
rect 33968 31340 34020 31346
rect 33968 31282 34020 31288
rect 33876 30932 33928 30938
rect 33876 30874 33928 30880
rect 33888 30598 33916 30874
rect 33980 30666 34008 31282
rect 34072 31226 34100 33254
rect 34934 33212 35242 33221
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33147 35242 33156
rect 34244 32904 34296 32910
rect 34244 32846 34296 32852
rect 34520 32904 34572 32910
rect 34520 32846 34572 32852
rect 34256 32570 34284 32846
rect 34244 32564 34296 32570
rect 34244 32506 34296 32512
rect 34152 32496 34204 32502
rect 34152 32438 34204 32444
rect 34164 31754 34192 32438
rect 34336 32428 34388 32434
rect 34336 32370 34388 32376
rect 34428 32428 34480 32434
rect 34428 32370 34480 32376
rect 34244 32224 34296 32230
rect 34244 32166 34296 32172
rect 34256 31958 34284 32166
rect 34244 31952 34296 31958
rect 34244 31894 34296 31900
rect 34164 31726 34284 31754
rect 34072 31198 34192 31226
rect 34060 31136 34112 31142
rect 34060 31078 34112 31084
rect 34072 30938 34100 31078
rect 34060 30932 34112 30938
rect 34060 30874 34112 30880
rect 34164 30870 34192 31198
rect 34152 30864 34204 30870
rect 34152 30806 34204 30812
rect 33968 30660 34020 30666
rect 34256 30648 34284 31726
rect 34348 31346 34376 32370
rect 34440 31668 34468 32370
rect 34532 32366 34560 32846
rect 35992 32836 36044 32842
rect 35992 32778 36044 32784
rect 36084 32836 36136 32842
rect 36084 32778 36136 32784
rect 35594 32668 35902 32677
rect 35594 32666 35600 32668
rect 35656 32666 35680 32668
rect 35736 32666 35760 32668
rect 35816 32666 35840 32668
rect 35896 32666 35902 32668
rect 35656 32614 35658 32666
rect 35838 32614 35840 32666
rect 35594 32612 35600 32614
rect 35656 32612 35680 32614
rect 35736 32612 35760 32614
rect 35816 32612 35840 32614
rect 35896 32612 35902 32614
rect 35594 32603 35902 32612
rect 36004 32570 36032 32778
rect 36096 32570 36124 32778
rect 36268 32768 36320 32774
rect 36268 32710 36320 32716
rect 35992 32564 36044 32570
rect 35992 32506 36044 32512
rect 36084 32564 36136 32570
rect 36084 32506 36136 32512
rect 35440 32496 35492 32502
rect 35440 32438 35492 32444
rect 34888 32428 34940 32434
rect 34888 32370 34940 32376
rect 34520 32360 34572 32366
rect 34900 32337 34928 32370
rect 34886 32328 34942 32337
rect 34520 32302 34572 32308
rect 34808 32286 34886 32314
rect 34808 31890 34836 32286
rect 34886 32263 34942 32272
rect 35452 32230 35480 32438
rect 36004 32298 36032 32506
rect 36280 32434 36308 32710
rect 36648 32570 36676 33322
rect 36820 32972 36872 32978
rect 36820 32914 36872 32920
rect 36728 32768 36780 32774
rect 36728 32710 36780 32716
rect 36636 32564 36688 32570
rect 36636 32506 36688 32512
rect 36268 32428 36320 32434
rect 36268 32370 36320 32376
rect 36740 32298 36768 32710
rect 35992 32292 36044 32298
rect 35992 32234 36044 32240
rect 36728 32292 36780 32298
rect 36728 32234 36780 32240
rect 35440 32224 35492 32230
rect 35440 32166 35492 32172
rect 34934 32124 35242 32133
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32059 35242 32068
rect 36740 31958 36768 32234
rect 36728 31952 36780 31958
rect 36728 31894 36780 31900
rect 34796 31884 34848 31890
rect 34796 31826 34848 31832
rect 34704 31816 34756 31822
rect 34704 31758 34756 31764
rect 34612 31748 34664 31754
rect 34612 31690 34664 31696
rect 34520 31680 34572 31686
rect 34440 31640 34520 31668
rect 34336 31340 34388 31346
rect 34336 31282 34388 31288
rect 34440 31278 34468 31640
rect 34520 31622 34572 31628
rect 34428 31272 34480 31278
rect 34428 31214 34480 31220
rect 34624 31142 34652 31690
rect 34716 31346 34744 31758
rect 35594 31580 35902 31589
rect 35594 31578 35600 31580
rect 35656 31578 35680 31580
rect 35736 31578 35760 31580
rect 35816 31578 35840 31580
rect 35896 31578 35902 31580
rect 35656 31526 35658 31578
rect 35838 31526 35840 31578
rect 35594 31524 35600 31526
rect 35656 31524 35680 31526
rect 35736 31524 35760 31526
rect 35816 31524 35840 31526
rect 35896 31524 35902 31526
rect 35594 31515 35902 31524
rect 36740 31482 36768 31894
rect 36832 31754 36860 32914
rect 37108 32910 37136 33798
rect 37464 33584 37516 33590
rect 37464 33526 37516 33532
rect 37280 33448 37332 33454
rect 37280 33390 37332 33396
rect 37292 33130 37320 33390
rect 37372 33312 37424 33318
rect 37372 33254 37424 33260
rect 37200 33102 37320 33130
rect 37200 33046 37228 33102
rect 37188 33040 37240 33046
rect 37188 32982 37240 32988
rect 37096 32904 37148 32910
rect 37096 32846 37148 32852
rect 37384 32026 37412 33254
rect 37476 33114 37504 33526
rect 38660 33516 38712 33522
rect 38660 33458 38712 33464
rect 37464 33108 37516 33114
rect 37464 33050 37516 33056
rect 37832 32836 37884 32842
rect 37832 32778 37884 32784
rect 37556 32768 37608 32774
rect 37556 32710 37608 32716
rect 37568 32502 37596 32710
rect 37556 32496 37608 32502
rect 37556 32438 37608 32444
rect 37844 32434 37872 32778
rect 38568 32768 38620 32774
rect 38672 32722 38700 33458
rect 39028 33312 39080 33318
rect 39028 33254 39080 33260
rect 39040 32842 39068 33254
rect 39028 32836 39080 32842
rect 39028 32778 39080 32784
rect 38620 32716 38700 32722
rect 38568 32710 38700 32716
rect 38580 32694 38700 32710
rect 37832 32428 37884 32434
rect 37832 32370 37884 32376
rect 37372 32020 37424 32026
rect 37372 31962 37424 31968
rect 37556 32020 37608 32026
rect 37556 31962 37608 31968
rect 36832 31726 36952 31754
rect 36728 31476 36780 31482
rect 36728 31418 36780 31424
rect 36636 31408 36688 31414
rect 36636 31350 36688 31356
rect 34704 31340 34756 31346
rect 34704 31282 34756 31288
rect 34716 31226 34744 31282
rect 36360 31272 36412 31278
rect 34716 31198 34836 31226
rect 36360 31214 36412 31220
rect 34612 31136 34664 31142
rect 34612 31078 34664 31084
rect 34704 31136 34756 31142
rect 34704 31078 34756 31084
rect 34624 30802 34652 31078
rect 34612 30796 34664 30802
rect 34612 30738 34664 30744
rect 34716 30734 34744 31078
rect 34808 30938 34836 31198
rect 34934 31036 35242 31045
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30971 35242 30980
rect 36372 30938 36400 31214
rect 34796 30932 34848 30938
rect 34796 30874 34848 30880
rect 36360 30932 36412 30938
rect 36360 30874 36412 30880
rect 36648 30734 36676 31350
rect 36820 31136 36872 31142
rect 36820 31078 36872 31084
rect 34704 30728 34756 30734
rect 34704 30670 34756 30676
rect 36636 30728 36688 30734
rect 36636 30670 36688 30676
rect 33968 30602 34020 30608
rect 34164 30620 34284 30648
rect 35348 30660 35400 30666
rect 33784 30592 33836 30598
rect 33782 30560 33784 30569
rect 33876 30592 33928 30598
rect 33836 30560 33838 30569
rect 33876 30534 33928 30540
rect 33782 30495 33838 30504
rect 33980 30410 34008 30602
rect 33600 30388 33652 30394
rect 33600 30330 33652 30336
rect 33888 30382 34008 30410
rect 33612 30054 33640 30330
rect 33888 30326 33916 30382
rect 33876 30320 33928 30326
rect 33876 30262 33928 30268
rect 34164 30258 34192 30620
rect 35348 30602 35400 30608
rect 34610 30560 34666 30569
rect 34610 30495 34666 30504
rect 34152 30252 34204 30258
rect 34152 30194 34204 30200
rect 33784 30184 33836 30190
rect 33784 30126 33836 30132
rect 33600 30048 33652 30054
rect 33600 29990 33652 29996
rect 33232 29776 33284 29782
rect 33232 29718 33284 29724
rect 32864 29572 32916 29578
rect 32864 29514 32916 29520
rect 32956 29572 33008 29578
rect 32956 29514 33008 29520
rect 32772 29504 32824 29510
rect 32772 29446 32824 29452
rect 32496 29232 32548 29238
rect 32496 29174 32548 29180
rect 32404 29096 32456 29102
rect 32404 29038 32456 29044
rect 32416 28762 32444 29038
rect 32404 28756 32456 28762
rect 32404 28698 32456 28704
rect 32508 28558 32536 29174
rect 32496 28552 32548 28558
rect 32496 28494 32548 28500
rect 32784 28490 32812 29446
rect 32876 28966 32904 29514
rect 32864 28960 32916 28966
rect 32864 28902 32916 28908
rect 33140 28960 33192 28966
rect 33140 28902 33192 28908
rect 32876 28558 32904 28902
rect 33152 28558 33180 28902
rect 32864 28552 32916 28558
rect 32864 28494 32916 28500
rect 33140 28552 33192 28558
rect 33140 28494 33192 28500
rect 30564 28484 30616 28490
rect 30564 28426 30616 28432
rect 32128 28484 32180 28490
rect 32128 28426 32180 28432
rect 32772 28484 32824 28490
rect 32772 28426 32824 28432
rect 30012 28416 30064 28422
rect 30012 28358 30064 28364
rect 30024 28218 30052 28358
rect 30012 28212 30064 28218
rect 30012 28154 30064 28160
rect 30576 27470 30604 28426
rect 30564 27464 30616 27470
rect 30564 27406 30616 27412
rect 30932 27464 30984 27470
rect 30932 27406 30984 27412
rect 32772 27464 32824 27470
rect 32772 27406 32824 27412
rect 29552 27396 29604 27402
rect 29552 27338 29604 27344
rect 29368 24608 29420 24614
rect 29368 24550 29420 24556
rect 29182 24440 29238 24449
rect 29182 24375 29238 24384
rect 29380 24274 29408 24550
rect 29368 24268 29420 24274
rect 29368 24210 29420 24216
rect 29092 24200 29144 24206
rect 29092 24142 29144 24148
rect 28828 23684 28948 23712
rect 28828 23526 28856 23684
rect 28908 23588 28960 23594
rect 28908 23530 28960 23536
rect 28816 23520 28868 23526
rect 28816 23462 28868 23468
rect 28816 23316 28868 23322
rect 28816 23258 28868 23264
rect 28828 23186 28856 23258
rect 28816 23180 28868 23186
rect 28816 23122 28868 23128
rect 28828 22642 28856 23122
rect 28816 22636 28868 22642
rect 28816 22578 28868 22584
rect 28724 21888 28776 21894
rect 28724 21830 28776 21836
rect 28632 21616 28684 21622
rect 28632 21558 28684 21564
rect 28540 21344 28592 21350
rect 28540 21286 28592 21292
rect 28552 20534 28580 21286
rect 28644 20874 28672 21558
rect 28632 20868 28684 20874
rect 28632 20810 28684 20816
rect 28540 20528 28592 20534
rect 28540 20470 28592 20476
rect 28644 20330 28672 20810
rect 28736 20466 28764 21830
rect 28816 20868 28868 20874
rect 28816 20810 28868 20816
rect 28724 20460 28776 20466
rect 28724 20402 28776 20408
rect 28828 20398 28856 20810
rect 28920 20641 28948 23530
rect 29000 23520 29052 23526
rect 29000 23462 29052 23468
rect 29012 22234 29040 23462
rect 29000 22228 29052 22234
rect 29000 22170 29052 22176
rect 29092 22092 29144 22098
rect 29092 22034 29144 22040
rect 28906 20632 28962 20641
rect 28906 20567 28962 20576
rect 28816 20392 28868 20398
rect 28816 20334 28868 20340
rect 28632 20324 28684 20330
rect 28632 20266 28684 20272
rect 28724 19984 28776 19990
rect 28724 19926 28776 19932
rect 28736 19786 28764 19926
rect 28816 19848 28868 19854
rect 28816 19790 28868 19796
rect 28724 19780 28776 19786
rect 28724 19722 28776 19728
rect 28540 19712 28592 19718
rect 28540 19654 28592 19660
rect 28552 19514 28580 19654
rect 28540 19508 28592 19514
rect 28540 19450 28592 19456
rect 28736 19378 28764 19722
rect 28828 19514 28856 19790
rect 28920 19718 28948 20567
rect 29104 20466 29132 22034
rect 29276 21616 29328 21622
rect 29276 21558 29328 21564
rect 29288 20534 29316 21558
rect 29276 20528 29328 20534
rect 29276 20470 29328 20476
rect 29092 20460 29144 20466
rect 29092 20402 29144 20408
rect 29368 20460 29420 20466
rect 29368 20402 29420 20408
rect 28908 19712 28960 19718
rect 28908 19654 28960 19660
rect 28920 19514 28948 19654
rect 28816 19508 28868 19514
rect 28816 19450 28868 19456
rect 28908 19508 28960 19514
rect 28908 19450 28960 19456
rect 28920 19394 28948 19450
rect 28724 19372 28776 19378
rect 28920 19366 29040 19394
rect 28724 19314 28776 19320
rect 28632 19304 28684 19310
rect 28632 19246 28684 19252
rect 28644 18834 28672 19246
rect 28632 18828 28684 18834
rect 28632 18770 28684 18776
rect 28736 15638 28764 19314
rect 28908 18692 28960 18698
rect 28908 18634 28960 18640
rect 28920 18426 28948 18634
rect 28908 18420 28960 18426
rect 28908 18362 28960 18368
rect 28920 16697 28948 18362
rect 29012 17338 29040 19366
rect 29000 17332 29052 17338
rect 29000 17274 29052 17280
rect 28906 16688 28962 16697
rect 28906 16623 28962 16632
rect 28920 16590 28948 16623
rect 29012 16590 29040 17274
rect 28908 16584 28960 16590
rect 28908 16526 28960 16532
rect 29000 16584 29052 16590
rect 29000 16526 29052 16532
rect 28724 15632 28776 15638
rect 28724 15574 28776 15580
rect 28632 14476 28684 14482
rect 28632 14418 28684 14424
rect 28644 13938 28672 14418
rect 28632 13932 28684 13938
rect 28632 13874 28684 13880
rect 28908 13864 28960 13870
rect 28908 13806 28960 13812
rect 28920 13530 28948 13806
rect 28908 13524 28960 13530
rect 28908 13466 28960 13472
rect 29104 13394 29132 20402
rect 29380 20262 29408 20402
rect 29368 20256 29420 20262
rect 29368 20198 29420 20204
rect 29184 20052 29236 20058
rect 29184 19994 29236 20000
rect 29196 16590 29224 19994
rect 29564 19786 29592 27338
rect 30196 26580 30248 26586
rect 30196 26522 30248 26528
rect 30208 26450 30236 26522
rect 29920 26444 29972 26450
rect 29920 26386 29972 26392
rect 30196 26444 30248 26450
rect 30196 26386 30248 26392
rect 29932 21554 29960 26386
rect 30208 26042 30236 26386
rect 30576 26314 30604 27406
rect 30944 27130 30972 27406
rect 32220 27396 32272 27402
rect 32220 27338 32272 27344
rect 30932 27124 30984 27130
rect 30932 27066 30984 27072
rect 32036 26988 32088 26994
rect 32036 26930 32088 26936
rect 30564 26308 30616 26314
rect 30564 26250 30616 26256
rect 30196 26036 30248 26042
rect 30196 25978 30248 25984
rect 30196 25424 30248 25430
rect 30196 25366 30248 25372
rect 30208 24954 30236 25366
rect 30576 25362 30604 26250
rect 30932 26240 30984 26246
rect 30932 26182 30984 26188
rect 30564 25356 30616 25362
rect 30564 25298 30616 25304
rect 30196 24948 30248 24954
rect 30196 24890 30248 24896
rect 30944 24206 30972 26182
rect 31760 25696 31812 25702
rect 31760 25638 31812 25644
rect 31772 25158 31800 25638
rect 31852 25492 31904 25498
rect 31852 25434 31904 25440
rect 31760 25152 31812 25158
rect 31760 25094 31812 25100
rect 31864 24954 31892 25434
rect 32048 25158 32076 26930
rect 32128 25900 32180 25906
rect 32128 25842 32180 25848
rect 32036 25152 32088 25158
rect 32036 25094 32088 25100
rect 31852 24948 31904 24954
rect 31852 24890 31904 24896
rect 32048 24886 32076 25094
rect 31484 24880 31536 24886
rect 31484 24822 31536 24828
rect 32036 24880 32088 24886
rect 32036 24822 32088 24828
rect 31392 24608 31444 24614
rect 31392 24550 31444 24556
rect 31404 24274 31432 24550
rect 31392 24268 31444 24274
rect 31392 24210 31444 24216
rect 30380 24200 30432 24206
rect 30380 24142 30432 24148
rect 30932 24200 30984 24206
rect 30932 24142 30984 24148
rect 31024 24200 31076 24206
rect 31024 24142 31076 24148
rect 30012 24064 30064 24070
rect 30012 24006 30064 24012
rect 30024 23594 30052 24006
rect 30012 23588 30064 23594
rect 30012 23530 30064 23536
rect 30392 23322 30420 24142
rect 30656 24064 30708 24070
rect 30656 24006 30708 24012
rect 30840 24064 30892 24070
rect 30840 24006 30892 24012
rect 30380 23316 30432 23322
rect 30380 23258 30432 23264
rect 30012 22500 30064 22506
rect 30012 22442 30064 22448
rect 29920 21548 29972 21554
rect 29920 21490 29972 21496
rect 29932 21026 29960 21490
rect 30024 21418 30052 22442
rect 30288 22228 30340 22234
rect 30288 22170 30340 22176
rect 30012 21412 30064 21418
rect 30012 21354 30064 21360
rect 29748 20998 29960 21026
rect 30024 21010 30052 21354
rect 30104 21344 30156 21350
rect 30104 21286 30156 21292
rect 30116 21146 30144 21286
rect 30300 21146 30328 22170
rect 30104 21140 30156 21146
rect 30104 21082 30156 21088
rect 30288 21140 30340 21146
rect 30288 21082 30340 21088
rect 30012 21004 30064 21010
rect 29748 20942 29776 20998
rect 30012 20946 30064 20952
rect 29644 20936 29696 20942
rect 29644 20878 29696 20884
rect 29736 20936 29788 20942
rect 29736 20878 29788 20884
rect 29828 20936 29880 20942
rect 29828 20878 29880 20884
rect 29656 20398 29684 20878
rect 29644 20392 29696 20398
rect 29644 20334 29696 20340
rect 29656 19922 29684 20334
rect 29644 19916 29696 19922
rect 29644 19858 29696 19864
rect 29552 19780 29604 19786
rect 29552 19722 29604 19728
rect 29748 19378 29776 20878
rect 29840 20602 29868 20878
rect 29920 20800 29972 20806
rect 29920 20742 29972 20748
rect 29828 20596 29880 20602
rect 29828 20538 29880 20544
rect 29932 20534 29960 20742
rect 29920 20528 29972 20534
rect 29920 20470 29972 20476
rect 30668 19854 30696 24006
rect 30656 19848 30708 19854
rect 30656 19790 30708 19796
rect 30852 19786 30880 24006
rect 31036 23186 31064 24142
rect 31496 24070 31524 24822
rect 31852 24812 31904 24818
rect 31852 24754 31904 24760
rect 31666 24712 31722 24721
rect 31666 24647 31722 24656
rect 31484 24064 31536 24070
rect 31484 24006 31536 24012
rect 31680 23866 31708 24647
rect 31760 24608 31812 24614
rect 31760 24550 31812 24556
rect 31772 24410 31800 24550
rect 31864 24410 31892 24754
rect 32140 24410 32168 25842
rect 32232 25226 32260 27338
rect 32496 27328 32548 27334
rect 32496 27270 32548 27276
rect 32508 26994 32536 27270
rect 32784 27130 32812 27406
rect 32772 27124 32824 27130
rect 32772 27066 32824 27072
rect 32404 26988 32456 26994
rect 32404 26930 32456 26936
rect 32496 26988 32548 26994
rect 32496 26930 32548 26936
rect 32864 26988 32916 26994
rect 32864 26930 32916 26936
rect 32956 26988 33008 26994
rect 33008 26948 33180 26976
rect 32956 26930 33008 26936
rect 32416 26586 32444 26930
rect 32876 26874 32904 26930
rect 32876 26846 32996 26874
rect 32864 26784 32916 26790
rect 32864 26726 32916 26732
rect 32404 26580 32456 26586
rect 32404 26522 32456 26528
rect 32876 26518 32904 26726
rect 32864 26512 32916 26518
rect 32864 26454 32916 26460
rect 32496 26376 32548 26382
rect 32548 26336 32628 26364
rect 32496 26318 32548 26324
rect 32404 26308 32456 26314
rect 32404 26250 32456 26256
rect 32416 25838 32444 26250
rect 32600 25906 32628 26336
rect 32588 25900 32640 25906
rect 32588 25842 32640 25848
rect 32404 25832 32456 25838
rect 32404 25774 32456 25780
rect 32220 25220 32272 25226
rect 32220 25162 32272 25168
rect 31760 24404 31812 24410
rect 31760 24346 31812 24352
rect 31852 24404 31904 24410
rect 31852 24346 31904 24352
rect 32128 24404 32180 24410
rect 32128 24346 32180 24352
rect 32232 24138 32260 25162
rect 32416 24800 32444 25774
rect 32496 24812 32548 24818
rect 32416 24772 32496 24800
rect 32496 24754 32548 24760
rect 32312 24676 32364 24682
rect 32312 24618 32364 24624
rect 32220 24132 32272 24138
rect 32220 24074 32272 24080
rect 32232 23866 32260 24074
rect 31668 23860 31720 23866
rect 31668 23802 31720 23808
rect 31760 23860 31812 23866
rect 31760 23802 31812 23808
rect 32220 23860 32272 23866
rect 32220 23802 32272 23808
rect 31024 23180 31076 23186
rect 31024 23122 31076 23128
rect 31772 23066 31800 23802
rect 32128 23724 32180 23730
rect 32128 23666 32180 23672
rect 32220 23724 32272 23730
rect 32220 23666 32272 23672
rect 31588 23050 31800 23066
rect 31576 23044 31800 23050
rect 31628 23038 31800 23044
rect 31576 22986 31628 22992
rect 31576 22568 31628 22574
rect 31576 22510 31628 22516
rect 31208 22024 31260 22030
rect 31208 21966 31260 21972
rect 31024 21888 31076 21894
rect 31024 21830 31076 21836
rect 31036 21690 31064 21830
rect 31024 21684 31076 21690
rect 31024 21626 31076 21632
rect 31220 21486 31248 21966
rect 31588 21554 31616 22510
rect 31680 21894 31708 23038
rect 32140 22710 32168 23666
rect 32232 23526 32260 23666
rect 32220 23520 32272 23526
rect 32220 23462 32272 23468
rect 32128 22704 32180 22710
rect 32128 22646 32180 22652
rect 32128 22432 32180 22438
rect 32128 22374 32180 22380
rect 32140 22098 32168 22374
rect 32128 22092 32180 22098
rect 32128 22034 32180 22040
rect 31944 21956 31996 21962
rect 31944 21898 31996 21904
rect 31668 21888 31720 21894
rect 31668 21830 31720 21836
rect 31576 21548 31628 21554
rect 31576 21490 31628 21496
rect 31208 21480 31260 21486
rect 31208 21422 31260 21428
rect 31220 20942 31248 21422
rect 31576 21344 31628 21350
rect 31576 21286 31628 21292
rect 31588 21010 31616 21286
rect 31576 21004 31628 21010
rect 31576 20946 31628 20952
rect 31208 20936 31260 20942
rect 31208 20878 31260 20884
rect 31116 20868 31168 20874
rect 31116 20810 31168 20816
rect 30932 20596 30984 20602
rect 30932 20538 30984 20544
rect 30944 20398 30972 20538
rect 31128 20398 31156 20810
rect 30932 20392 30984 20398
rect 30932 20334 30984 20340
rect 31116 20392 31168 20398
rect 31116 20334 31168 20340
rect 31220 19990 31248 20878
rect 31956 20874 31984 21898
rect 32232 21894 32260 23462
rect 32324 23225 32352 24618
rect 32508 23526 32536 24754
rect 32600 24750 32628 25842
rect 32876 25430 32904 26454
rect 32968 25974 32996 26846
rect 33152 26382 33180 26948
rect 33048 26376 33100 26382
rect 33048 26318 33100 26324
rect 33140 26376 33192 26382
rect 33140 26318 33192 26324
rect 32956 25968 33008 25974
rect 32956 25910 33008 25916
rect 32864 25424 32916 25430
rect 32864 25366 32916 25372
rect 32680 24812 32732 24818
rect 32680 24754 32732 24760
rect 32588 24744 32640 24750
rect 32588 24686 32640 24692
rect 32588 24404 32640 24410
rect 32588 24346 32640 24352
rect 32600 23798 32628 24346
rect 32692 24138 32720 24754
rect 32772 24608 32824 24614
rect 32772 24550 32824 24556
rect 32680 24132 32732 24138
rect 32680 24074 32732 24080
rect 32588 23792 32640 23798
rect 32588 23734 32640 23740
rect 32496 23520 32548 23526
rect 32496 23462 32548 23468
rect 32680 23520 32732 23526
rect 32680 23462 32732 23468
rect 32310 23216 32366 23225
rect 32310 23151 32366 23160
rect 32586 23216 32642 23225
rect 32586 23151 32642 23160
rect 32600 23118 32628 23151
rect 32692 23118 32720 23462
rect 32588 23112 32640 23118
rect 32588 23054 32640 23060
rect 32680 23112 32732 23118
rect 32680 23054 32732 23060
rect 32312 22976 32364 22982
rect 32312 22918 32364 22924
rect 32220 21888 32272 21894
rect 32220 21830 32272 21836
rect 32232 21554 32260 21830
rect 32324 21690 32352 22918
rect 32404 22636 32456 22642
rect 32404 22578 32456 22584
rect 32680 22636 32732 22642
rect 32680 22578 32732 22584
rect 32312 21684 32364 21690
rect 32416 21672 32444 22578
rect 32692 22234 32720 22578
rect 32784 22506 32812 24550
rect 32876 23186 32904 25366
rect 32968 23798 32996 25910
rect 33060 25226 33088 26318
rect 33244 26246 33272 29718
rect 33796 29646 33824 30126
rect 33968 30048 34020 30054
rect 33968 29990 34020 29996
rect 33980 29646 34008 29990
rect 33784 29640 33836 29646
rect 33784 29582 33836 29588
rect 33968 29640 34020 29646
rect 33968 29582 34020 29588
rect 33796 28762 33824 29582
rect 33980 29306 34008 29582
rect 34164 29578 34192 30194
rect 34624 30054 34652 30495
rect 35360 30394 35388 30602
rect 35594 30492 35902 30501
rect 35594 30490 35600 30492
rect 35656 30490 35680 30492
rect 35736 30490 35760 30492
rect 35816 30490 35840 30492
rect 35896 30490 35902 30492
rect 35656 30438 35658 30490
rect 35838 30438 35840 30490
rect 35594 30436 35600 30438
rect 35656 30436 35680 30438
rect 35736 30436 35760 30438
rect 35816 30436 35840 30438
rect 35896 30436 35902 30438
rect 35594 30427 35902 30436
rect 35348 30388 35400 30394
rect 35348 30330 35400 30336
rect 36648 30326 36676 30670
rect 36832 30598 36860 31078
rect 36924 30734 36952 31726
rect 36912 30728 36964 30734
rect 36912 30670 36964 30676
rect 36820 30592 36872 30598
rect 36820 30534 36872 30540
rect 36636 30320 36688 30326
rect 36636 30262 36688 30268
rect 36648 30122 36676 30262
rect 36924 30190 36952 30670
rect 37280 30660 37332 30666
rect 37280 30602 37332 30608
rect 36912 30184 36964 30190
rect 36912 30126 36964 30132
rect 36636 30116 36688 30122
rect 36636 30058 36688 30064
rect 34612 30048 34664 30054
rect 34612 29990 34664 29996
rect 36544 30048 36596 30054
rect 36544 29990 36596 29996
rect 34934 29948 35242 29957
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29883 35242 29892
rect 34152 29572 34204 29578
rect 34152 29514 34204 29520
rect 34980 29504 35032 29510
rect 34980 29446 35032 29452
rect 33968 29300 34020 29306
rect 33968 29242 34020 29248
rect 34992 29102 35020 29446
rect 35594 29404 35902 29413
rect 35594 29402 35600 29404
rect 35656 29402 35680 29404
rect 35736 29402 35760 29404
rect 35816 29402 35840 29404
rect 35896 29402 35902 29404
rect 35656 29350 35658 29402
rect 35838 29350 35840 29402
rect 35594 29348 35600 29350
rect 35656 29348 35680 29350
rect 35736 29348 35760 29350
rect 35816 29348 35840 29350
rect 35896 29348 35902 29350
rect 35594 29339 35902 29348
rect 35992 29164 36044 29170
rect 35992 29106 36044 29112
rect 34980 29096 35032 29102
rect 34980 29038 35032 29044
rect 34934 28860 35242 28869
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28795 35242 28804
rect 33784 28756 33836 28762
rect 33784 28698 33836 28704
rect 36004 28626 36032 29106
rect 35992 28620 36044 28626
rect 35992 28562 36044 28568
rect 36268 28484 36320 28490
rect 36268 28426 36320 28432
rect 35594 28316 35902 28325
rect 35594 28314 35600 28316
rect 35656 28314 35680 28316
rect 35736 28314 35760 28316
rect 35816 28314 35840 28316
rect 35896 28314 35902 28316
rect 35656 28262 35658 28314
rect 35838 28262 35840 28314
rect 35594 28260 35600 28262
rect 35656 28260 35680 28262
rect 35736 28260 35760 28262
rect 35816 28260 35840 28262
rect 35896 28260 35902 28262
rect 35594 28251 35902 28260
rect 36280 28218 36308 28426
rect 36268 28212 36320 28218
rect 36268 28154 36320 28160
rect 36556 28150 36584 29990
rect 36924 29170 36952 30126
rect 37292 29850 37320 30602
rect 37464 30048 37516 30054
rect 37464 29990 37516 29996
rect 37280 29844 37332 29850
rect 37280 29786 37332 29792
rect 37476 29578 37504 29990
rect 37568 29850 37596 31962
rect 38384 31884 38436 31890
rect 38384 31826 38436 31832
rect 37832 31816 37884 31822
rect 37832 31758 37884 31764
rect 37844 30938 37872 31758
rect 37924 31748 37976 31754
rect 37924 31690 37976 31696
rect 37936 31482 37964 31690
rect 37924 31476 37976 31482
rect 37924 31418 37976 31424
rect 37832 30932 37884 30938
rect 37832 30874 37884 30880
rect 37556 29844 37608 29850
rect 37556 29786 37608 29792
rect 37844 29782 37872 30874
rect 37832 29776 37884 29782
rect 37832 29718 37884 29724
rect 38200 29708 38252 29714
rect 38200 29650 38252 29656
rect 37464 29572 37516 29578
rect 37464 29514 37516 29520
rect 37648 29504 37700 29510
rect 37648 29446 37700 29452
rect 37660 29238 37688 29446
rect 38016 29300 38068 29306
rect 38016 29242 38068 29248
rect 37648 29232 37700 29238
rect 37648 29174 37700 29180
rect 36912 29164 36964 29170
rect 36912 29106 36964 29112
rect 38028 28762 38056 29242
rect 38212 28762 38240 29650
rect 38016 28756 38068 28762
rect 38016 28698 38068 28704
rect 38200 28756 38252 28762
rect 38200 28698 38252 28704
rect 38028 28490 38056 28698
rect 38396 28490 38424 31826
rect 38672 31414 38700 32694
rect 38752 31952 38804 31958
rect 38752 31894 38804 31900
rect 38764 31414 38792 31894
rect 38660 31408 38712 31414
rect 38660 31350 38712 31356
rect 38752 31408 38804 31414
rect 38752 31350 38804 31356
rect 38672 31278 38700 31350
rect 38660 31272 38712 31278
rect 38660 31214 38712 31220
rect 38568 30660 38620 30666
rect 38672 30648 38700 31214
rect 38752 31136 38804 31142
rect 38752 31078 38804 31084
rect 38764 30666 38792 31078
rect 38620 30620 38700 30648
rect 38568 30602 38620 30608
rect 38568 30252 38620 30258
rect 38568 30194 38620 30200
rect 38580 30122 38608 30194
rect 38568 30116 38620 30122
rect 38568 30058 38620 30064
rect 38016 28484 38068 28490
rect 38016 28426 38068 28432
rect 38384 28484 38436 28490
rect 38384 28426 38436 28432
rect 37740 28416 37792 28422
rect 37740 28358 37792 28364
rect 36544 28144 36596 28150
rect 36544 28086 36596 28092
rect 37752 28014 37780 28358
rect 37832 28144 37884 28150
rect 37832 28086 37884 28092
rect 37844 28014 37872 28086
rect 37740 28008 37792 28014
rect 37740 27950 37792 27956
rect 37832 28008 37884 28014
rect 37832 27950 37884 27956
rect 34934 27772 35242 27781
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27707 35242 27716
rect 37648 27464 37700 27470
rect 37648 27406 37700 27412
rect 34704 27396 34756 27402
rect 34704 27338 34756 27344
rect 36268 27396 36320 27402
rect 36268 27338 36320 27344
rect 33324 27328 33376 27334
rect 33324 27270 33376 27276
rect 34520 27328 34572 27334
rect 34520 27270 34572 27276
rect 33336 26994 33364 27270
rect 34532 27130 34560 27270
rect 34520 27124 34572 27130
rect 34520 27066 34572 27072
rect 33324 26988 33376 26994
rect 33324 26930 33376 26936
rect 33692 26988 33744 26994
rect 33692 26930 33744 26936
rect 33336 26450 33364 26930
rect 33704 26518 33732 26930
rect 34612 26920 34664 26926
rect 34612 26862 34664 26868
rect 34520 26852 34572 26858
rect 34520 26794 34572 26800
rect 33692 26512 33744 26518
rect 33692 26454 33744 26460
rect 34532 26450 34560 26794
rect 33324 26444 33376 26450
rect 33324 26386 33376 26392
rect 34520 26444 34572 26450
rect 34520 26386 34572 26392
rect 34428 26376 34480 26382
rect 34428 26318 34480 26324
rect 33232 26240 33284 26246
rect 33232 26182 33284 26188
rect 33324 25696 33376 25702
rect 33324 25638 33376 25644
rect 33336 25294 33364 25638
rect 34336 25492 34388 25498
rect 34336 25434 34388 25440
rect 33232 25288 33284 25294
rect 33232 25230 33284 25236
rect 33324 25288 33376 25294
rect 33324 25230 33376 25236
rect 33048 25220 33100 25226
rect 33048 25162 33100 25168
rect 33060 24886 33088 25162
rect 33244 25158 33272 25230
rect 33232 25152 33284 25158
rect 33232 25094 33284 25100
rect 33048 24880 33100 24886
rect 33048 24822 33100 24828
rect 33140 24880 33192 24886
rect 33140 24822 33192 24828
rect 33244 24834 33272 25094
rect 33060 24274 33088 24822
rect 33152 24410 33180 24822
rect 33244 24806 33364 24834
rect 33232 24744 33284 24750
rect 33232 24686 33284 24692
rect 33140 24404 33192 24410
rect 33140 24346 33192 24352
rect 33048 24268 33100 24274
rect 33048 24210 33100 24216
rect 33140 24200 33192 24206
rect 33140 24142 33192 24148
rect 33048 24132 33100 24138
rect 33048 24074 33100 24080
rect 32956 23792 33008 23798
rect 32956 23734 33008 23740
rect 32864 23180 32916 23186
rect 32864 23122 32916 23128
rect 32772 22500 32824 22506
rect 32772 22442 32824 22448
rect 32680 22228 32732 22234
rect 32680 22170 32732 22176
rect 32496 21684 32548 21690
rect 32416 21644 32496 21672
rect 32312 21626 32364 21632
rect 32496 21626 32548 21632
rect 32784 21554 32812 22442
rect 32876 22438 32904 23122
rect 33060 23118 33088 24074
rect 33152 23866 33180 24142
rect 33140 23860 33192 23866
rect 33140 23802 33192 23808
rect 33140 23724 33192 23730
rect 33140 23666 33192 23672
rect 33048 23112 33100 23118
rect 33048 23054 33100 23060
rect 33152 22438 33180 23666
rect 33244 22574 33272 24686
rect 33336 23225 33364 24806
rect 33416 24812 33468 24818
rect 33416 24754 33468 24760
rect 33428 23730 33456 24754
rect 34058 24440 34114 24449
rect 34058 24375 34060 24384
rect 34112 24375 34114 24384
rect 34060 24346 34112 24352
rect 34348 24313 34376 25434
rect 34440 24750 34468 26318
rect 34428 24744 34480 24750
rect 34428 24686 34480 24692
rect 34520 24608 34572 24614
rect 34520 24550 34572 24556
rect 34532 24410 34560 24550
rect 34520 24404 34572 24410
rect 34520 24346 34572 24352
rect 33966 24304 34022 24313
rect 33966 24239 34022 24248
rect 34334 24304 34390 24313
rect 34334 24239 34390 24248
rect 33980 24206 34008 24239
rect 33968 24200 34020 24206
rect 33968 24142 34020 24148
rect 33980 24070 34008 24142
rect 33968 24064 34020 24070
rect 33968 24006 34020 24012
rect 33692 23792 33744 23798
rect 33692 23734 33744 23740
rect 33416 23724 33468 23730
rect 33416 23666 33468 23672
rect 33598 23624 33654 23633
rect 33598 23559 33654 23568
rect 33612 23526 33640 23559
rect 33600 23520 33652 23526
rect 33600 23462 33652 23468
rect 33322 23216 33378 23225
rect 33704 23186 33732 23734
rect 33322 23151 33378 23160
rect 33692 23180 33744 23186
rect 33692 23122 33744 23128
rect 33980 22982 34008 24006
rect 34348 23798 34376 24239
rect 34520 24200 34572 24206
rect 34520 24142 34572 24148
rect 34336 23792 34388 23798
rect 34336 23734 34388 23740
rect 33968 22976 34020 22982
rect 33968 22918 34020 22924
rect 33232 22568 33284 22574
rect 33232 22510 33284 22516
rect 34428 22500 34480 22506
rect 34428 22442 34480 22448
rect 32864 22432 32916 22438
rect 32864 22374 32916 22380
rect 33140 22432 33192 22438
rect 33140 22374 33192 22380
rect 33600 22432 33652 22438
rect 33600 22374 33652 22380
rect 32876 21690 32904 22374
rect 33140 22160 33192 22166
rect 33140 22102 33192 22108
rect 32864 21684 32916 21690
rect 32864 21626 32916 21632
rect 32220 21548 32272 21554
rect 32220 21490 32272 21496
rect 32772 21548 32824 21554
rect 32772 21490 32824 21496
rect 32876 21350 32904 21626
rect 33152 21418 33180 22102
rect 33612 22030 33640 22374
rect 34440 22234 34468 22442
rect 34428 22228 34480 22234
rect 34428 22170 34480 22176
rect 33600 22024 33652 22030
rect 33600 21966 33652 21972
rect 33612 21622 33640 21966
rect 34532 21690 34560 24142
rect 34624 22778 34652 26862
rect 34716 26586 34744 27338
rect 35594 27228 35902 27237
rect 35594 27226 35600 27228
rect 35656 27226 35680 27228
rect 35736 27226 35760 27228
rect 35816 27226 35840 27228
rect 35896 27226 35902 27228
rect 35656 27174 35658 27226
rect 35838 27174 35840 27226
rect 35594 27172 35600 27174
rect 35656 27172 35680 27174
rect 35736 27172 35760 27174
rect 35816 27172 35840 27174
rect 35896 27172 35902 27174
rect 35594 27163 35902 27172
rect 35992 27124 36044 27130
rect 35992 27066 36044 27072
rect 34888 26988 34940 26994
rect 34888 26930 34940 26936
rect 34900 26858 34928 26930
rect 34888 26852 34940 26858
rect 34888 26794 34940 26800
rect 34796 26784 34848 26790
rect 34796 26726 34848 26732
rect 34704 26580 34756 26586
rect 34704 26522 34756 26528
rect 34808 26450 34836 26726
rect 34934 26684 35242 26693
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26619 35242 26628
rect 35164 26580 35216 26586
rect 35164 26522 35216 26528
rect 35808 26580 35860 26586
rect 35808 26522 35860 26528
rect 34704 26444 34756 26450
rect 34704 26386 34756 26392
rect 34796 26444 34848 26450
rect 34796 26386 34848 26392
rect 34612 22772 34664 22778
rect 34612 22714 34664 22720
rect 34624 22094 34652 22714
rect 34716 22642 34744 26386
rect 35072 26376 35124 26382
rect 35070 26344 35072 26353
rect 35124 26344 35126 26353
rect 35070 26279 35126 26288
rect 35176 25906 35204 26522
rect 35624 26376 35676 26382
rect 35544 26336 35624 26364
rect 35544 26246 35572 26336
rect 35820 26364 35848 26522
rect 35900 26512 35952 26518
rect 35898 26480 35900 26489
rect 35952 26480 35954 26489
rect 35898 26415 35954 26424
rect 35900 26376 35952 26382
rect 35820 26336 35900 26364
rect 35624 26318 35676 26324
rect 35900 26318 35952 26324
rect 35256 26240 35308 26246
rect 35256 26182 35308 26188
rect 35532 26240 35584 26246
rect 35532 26182 35584 26188
rect 35164 25900 35216 25906
rect 35164 25842 35216 25848
rect 35268 25838 35296 26182
rect 35594 26140 35902 26149
rect 35594 26138 35600 26140
rect 35656 26138 35680 26140
rect 35736 26138 35760 26140
rect 35816 26138 35840 26140
rect 35896 26138 35902 26140
rect 35656 26086 35658 26138
rect 35838 26086 35840 26138
rect 35594 26084 35600 26086
rect 35656 26084 35680 26086
rect 35736 26084 35760 26086
rect 35816 26084 35840 26086
rect 35896 26084 35902 26086
rect 35594 26075 35902 26084
rect 35532 26036 35584 26042
rect 35532 25978 35584 25984
rect 35544 25838 35572 25978
rect 35624 25968 35676 25974
rect 35624 25910 35676 25916
rect 35256 25832 35308 25838
rect 35256 25774 35308 25780
rect 35532 25832 35584 25838
rect 35532 25774 35584 25780
rect 35636 25702 35664 25910
rect 35808 25900 35860 25906
rect 35808 25842 35860 25848
rect 35532 25696 35584 25702
rect 35532 25638 35584 25644
rect 35624 25696 35676 25702
rect 35624 25638 35676 25644
rect 34934 25596 35242 25605
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25531 35242 25540
rect 34980 25356 35032 25362
rect 34980 25298 35032 25304
rect 34992 24818 35020 25298
rect 35072 25288 35124 25294
rect 35072 25230 35124 25236
rect 35084 24818 35112 25230
rect 35544 25140 35572 25638
rect 35452 25112 35572 25140
rect 35820 25140 35848 25842
rect 36004 25294 36032 27066
rect 36280 27062 36308 27338
rect 36728 27328 36780 27334
rect 36728 27270 36780 27276
rect 36544 27124 36596 27130
rect 36544 27066 36596 27072
rect 36268 27056 36320 27062
rect 36268 26998 36320 27004
rect 36084 26784 36136 26790
rect 36084 26726 36136 26732
rect 36096 25906 36124 26726
rect 36450 26480 36506 26489
rect 36450 26415 36506 26424
rect 36464 26382 36492 26415
rect 36360 26376 36412 26382
rect 36358 26344 36360 26353
rect 36452 26376 36504 26382
rect 36412 26344 36414 26353
rect 36268 26308 36320 26314
rect 36452 26318 36504 26324
rect 36358 26279 36414 26288
rect 36268 26250 36320 26256
rect 36176 26240 36228 26246
rect 36176 26182 36228 26188
rect 36084 25900 36136 25906
rect 36084 25842 36136 25848
rect 35992 25288 36044 25294
rect 35992 25230 36044 25236
rect 36084 25220 36136 25226
rect 36084 25162 36136 25168
rect 35820 25112 36032 25140
rect 36096 25129 36124 25162
rect 35452 24886 35480 25112
rect 35594 25052 35902 25061
rect 35594 25050 35600 25052
rect 35656 25050 35680 25052
rect 35736 25050 35760 25052
rect 35816 25050 35840 25052
rect 35896 25050 35902 25052
rect 35656 24998 35658 25050
rect 35838 24998 35840 25050
rect 35594 24996 35600 24998
rect 35656 24996 35680 24998
rect 35736 24996 35760 24998
rect 35816 24996 35840 24998
rect 35896 24996 35902 24998
rect 35594 24987 35902 24996
rect 35440 24880 35492 24886
rect 35440 24822 35492 24828
rect 34980 24812 35032 24818
rect 34808 24772 34980 24800
rect 34808 24274 34836 24772
rect 34980 24754 35032 24760
rect 35072 24812 35124 24818
rect 35072 24754 35124 24760
rect 35716 24812 35768 24818
rect 35716 24754 35768 24760
rect 34934 24508 35242 24517
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24443 35242 24452
rect 34980 24336 35032 24342
rect 34980 24278 35032 24284
rect 35256 24336 35308 24342
rect 35256 24278 35308 24284
rect 35622 24304 35678 24313
rect 34796 24268 34848 24274
rect 34796 24210 34848 24216
rect 34992 23866 35020 24278
rect 35162 24168 35218 24177
rect 35162 24103 35218 24112
rect 34980 23860 35032 23866
rect 34980 23802 35032 23808
rect 35176 23730 35204 24103
rect 35268 23730 35296 24278
rect 35348 24268 35400 24274
rect 35622 24239 35678 24248
rect 35348 24210 35400 24216
rect 34888 23724 34940 23730
rect 34888 23666 34940 23672
rect 35164 23724 35216 23730
rect 35164 23666 35216 23672
rect 35256 23724 35308 23730
rect 35256 23666 35308 23672
rect 34796 23656 34848 23662
rect 34796 23598 34848 23604
rect 34808 23322 34836 23598
rect 34900 23526 34928 23666
rect 34888 23520 34940 23526
rect 34888 23462 34940 23468
rect 34934 23420 35242 23429
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23355 35242 23364
rect 34796 23316 34848 23322
rect 34796 23258 34848 23264
rect 34808 22710 34836 23258
rect 35360 23186 35388 24210
rect 35636 24206 35664 24239
rect 35624 24200 35676 24206
rect 35624 24142 35676 24148
rect 35728 24138 35756 24754
rect 36004 24410 36032 25112
rect 36082 25120 36138 25129
rect 36082 25055 36138 25064
rect 36084 24744 36136 24750
rect 36188 24732 36216 26182
rect 36280 25498 36308 26250
rect 36268 25492 36320 25498
rect 36268 25434 36320 25440
rect 36280 24818 36308 25434
rect 36268 24812 36320 24818
rect 36268 24754 36320 24760
rect 36136 24704 36216 24732
rect 36084 24686 36136 24692
rect 36096 24410 36124 24686
rect 36372 24562 36400 26279
rect 36556 25226 36584 27066
rect 36636 26920 36688 26926
rect 36636 26862 36688 26868
rect 36648 26586 36676 26862
rect 36636 26580 36688 26586
rect 36636 26522 36688 26528
rect 36740 26518 36768 27270
rect 37660 26994 37688 27406
rect 37844 27130 37872 27950
rect 37832 27124 37884 27130
rect 37832 27066 37884 27072
rect 37648 26988 37700 26994
rect 37648 26930 37700 26936
rect 36820 26920 36872 26926
rect 36820 26862 36872 26868
rect 36728 26512 36780 26518
rect 36728 26454 36780 26460
rect 36728 25832 36780 25838
rect 36728 25774 36780 25780
rect 36544 25220 36596 25226
rect 36544 25162 36596 25168
rect 36372 24534 36492 24562
rect 35992 24404 36044 24410
rect 35992 24346 36044 24352
rect 36084 24404 36136 24410
rect 36084 24346 36136 24352
rect 36360 24336 36412 24342
rect 36360 24278 36412 24284
rect 35900 24268 35952 24274
rect 35952 24228 36308 24256
rect 35900 24210 35952 24216
rect 36084 24166 36136 24172
rect 35716 24132 35768 24138
rect 35716 24074 35768 24080
rect 35900 24132 35952 24138
rect 35952 24092 36032 24120
rect 36136 24126 36216 24154
rect 36084 24108 36136 24114
rect 35900 24074 35952 24080
rect 36004 24041 36032 24092
rect 35990 24032 36046 24041
rect 35594 23964 35902 23973
rect 35990 23967 36046 23976
rect 35594 23962 35600 23964
rect 35656 23962 35680 23964
rect 35736 23962 35760 23964
rect 35816 23962 35840 23964
rect 35896 23962 35902 23964
rect 35656 23910 35658 23962
rect 35838 23910 35840 23962
rect 35594 23908 35600 23910
rect 35656 23908 35680 23910
rect 35736 23908 35760 23910
rect 35816 23908 35840 23910
rect 35896 23908 35902 23910
rect 35594 23899 35902 23908
rect 35440 23860 35492 23866
rect 35440 23802 35492 23808
rect 35452 23769 35480 23802
rect 35438 23760 35494 23769
rect 35438 23695 35440 23704
rect 35492 23695 35494 23704
rect 35440 23666 35492 23672
rect 36188 23662 36216 24126
rect 35808 23656 35860 23662
rect 35808 23598 35860 23604
rect 36176 23656 36228 23662
rect 36176 23598 36228 23604
rect 35348 23180 35400 23186
rect 35400 23140 35480 23168
rect 35348 23122 35400 23128
rect 35346 23080 35402 23089
rect 35346 23015 35402 23024
rect 34796 22704 34848 22710
rect 34796 22646 34848 22652
rect 35360 22642 35388 23015
rect 34704 22636 34756 22642
rect 34704 22578 34756 22584
rect 35348 22636 35400 22642
rect 35348 22578 35400 22584
rect 35348 22432 35400 22438
rect 35348 22374 35400 22380
rect 34934 22332 35242 22341
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22267 35242 22276
rect 34624 22066 34836 22094
rect 34612 22024 34664 22030
rect 34612 21966 34664 21972
rect 34520 21684 34572 21690
rect 34520 21626 34572 21632
rect 33600 21616 33652 21622
rect 33600 21558 33652 21564
rect 34060 21548 34112 21554
rect 34060 21490 34112 21496
rect 34152 21548 34204 21554
rect 34152 21490 34204 21496
rect 34428 21548 34480 21554
rect 34428 21490 34480 21496
rect 34520 21548 34572 21554
rect 34520 21490 34572 21496
rect 33140 21412 33192 21418
rect 33140 21354 33192 21360
rect 32864 21344 32916 21350
rect 32864 21286 32916 21292
rect 31944 20868 31996 20874
rect 31944 20810 31996 20816
rect 31300 20800 31352 20806
rect 31300 20742 31352 20748
rect 31312 20534 31340 20742
rect 31300 20528 31352 20534
rect 31300 20470 31352 20476
rect 31758 20496 31814 20505
rect 31758 20431 31814 20440
rect 31392 20392 31444 20398
rect 31392 20334 31444 20340
rect 31208 19984 31260 19990
rect 31208 19926 31260 19932
rect 31404 19854 31432 20334
rect 31576 19984 31628 19990
rect 31628 19944 31708 19972
rect 31576 19926 31628 19932
rect 31392 19848 31444 19854
rect 31576 19848 31628 19854
rect 31392 19790 31444 19796
rect 31496 19808 31576 19836
rect 30840 19780 30892 19786
rect 30840 19722 30892 19728
rect 29828 19712 29880 19718
rect 29828 19654 29880 19660
rect 30380 19712 30432 19718
rect 30380 19654 30432 19660
rect 29736 19372 29788 19378
rect 29736 19314 29788 19320
rect 29840 19281 29868 19654
rect 30288 19440 30340 19446
rect 30288 19382 30340 19388
rect 30196 19372 30248 19378
rect 30196 19314 30248 19320
rect 29826 19272 29882 19281
rect 29748 19230 29826 19258
rect 29368 18624 29420 18630
rect 29368 18566 29420 18572
rect 29380 18358 29408 18566
rect 29368 18352 29420 18358
rect 29368 18294 29420 18300
rect 29460 18148 29512 18154
rect 29460 18090 29512 18096
rect 29368 17128 29420 17134
rect 29368 17070 29420 17076
rect 29380 16590 29408 17070
rect 29472 16998 29500 18090
rect 29460 16992 29512 16998
rect 29460 16934 29512 16940
rect 29644 16992 29696 16998
rect 29644 16934 29696 16940
rect 29184 16584 29236 16590
rect 29184 16526 29236 16532
rect 29368 16584 29420 16590
rect 29472 16561 29500 16934
rect 29552 16584 29604 16590
rect 29368 16526 29420 16532
rect 29458 16552 29514 16561
rect 29196 16250 29224 16526
rect 29184 16244 29236 16250
rect 29184 16186 29236 16192
rect 29276 16176 29328 16182
rect 29380 16164 29408 16526
rect 29552 16526 29604 16532
rect 29458 16487 29514 16496
rect 29564 16454 29592 16526
rect 29552 16448 29604 16454
rect 29552 16390 29604 16396
rect 29328 16136 29408 16164
rect 29276 16118 29328 16124
rect 29564 15484 29592 16390
rect 29656 16182 29684 16934
rect 29644 16176 29696 16182
rect 29644 16118 29696 16124
rect 29748 15910 29776 19230
rect 29826 19207 29882 19216
rect 30208 18290 30236 19314
rect 30300 18766 30328 19382
rect 30392 18970 30420 19654
rect 31496 19378 31524 19808
rect 31576 19790 31628 19796
rect 31680 19378 31708 19944
rect 31772 19854 31800 20431
rect 33600 20392 33652 20398
rect 33600 20334 33652 20340
rect 32036 19916 32088 19922
rect 32036 19858 32088 19864
rect 31760 19848 31812 19854
rect 31760 19790 31812 19796
rect 31484 19372 31536 19378
rect 31484 19314 31536 19320
rect 31668 19372 31720 19378
rect 32048 19334 32076 19858
rect 32220 19712 32272 19718
rect 32220 19654 32272 19660
rect 31668 19314 31720 19320
rect 30564 19304 30616 19310
rect 30564 19246 30616 19252
rect 30576 18970 30604 19246
rect 31024 19168 31076 19174
rect 31024 19110 31076 19116
rect 30380 18964 30432 18970
rect 30380 18906 30432 18912
rect 30564 18964 30616 18970
rect 30564 18906 30616 18912
rect 30564 18828 30616 18834
rect 30564 18770 30616 18776
rect 30288 18760 30340 18766
rect 30288 18702 30340 18708
rect 30576 18290 30604 18770
rect 30748 18760 30800 18766
rect 30748 18702 30800 18708
rect 30760 18290 30788 18702
rect 30840 18692 30892 18698
rect 30840 18634 30892 18640
rect 30196 18284 30248 18290
rect 30196 18226 30248 18232
rect 30564 18284 30616 18290
rect 30564 18226 30616 18232
rect 30748 18284 30800 18290
rect 30748 18226 30800 18232
rect 30104 18216 30156 18222
rect 30104 18158 30156 18164
rect 29918 17232 29974 17241
rect 29828 17196 29880 17202
rect 29918 17167 29920 17176
rect 29828 17138 29880 17144
rect 29972 17167 29974 17176
rect 29920 17138 29972 17144
rect 29840 16794 29868 17138
rect 29828 16788 29880 16794
rect 29828 16730 29880 16736
rect 29828 16584 29880 16590
rect 29828 16526 29880 16532
rect 29736 15904 29788 15910
rect 29736 15846 29788 15852
rect 29644 15496 29696 15502
rect 29564 15456 29644 15484
rect 29644 15438 29696 15444
rect 29092 13388 29144 13394
rect 29092 13330 29144 13336
rect 29656 13258 29684 15438
rect 29840 15434 29868 16526
rect 29828 15428 29880 15434
rect 29828 15370 29880 15376
rect 29932 14498 29960 17138
rect 30116 16454 30144 18158
rect 30380 17740 30432 17746
rect 30380 17682 30432 17688
rect 30288 17672 30340 17678
rect 30288 17614 30340 17620
rect 30300 16998 30328 17614
rect 30288 16992 30340 16998
rect 30288 16934 30340 16940
rect 30196 16516 30248 16522
rect 30196 16458 30248 16464
rect 30104 16448 30156 16454
rect 30104 16390 30156 16396
rect 30208 15570 30236 16458
rect 30392 16250 30420 17682
rect 30472 17536 30524 17542
rect 30472 17478 30524 17484
rect 30484 16590 30512 17478
rect 30576 16726 30604 18226
rect 30760 17542 30788 18226
rect 30748 17536 30800 17542
rect 30748 17478 30800 17484
rect 30656 17196 30708 17202
rect 30656 17138 30708 17144
rect 30668 16794 30696 17138
rect 30748 17128 30800 17134
rect 30748 17070 30800 17076
rect 30760 16969 30788 17070
rect 30746 16960 30802 16969
rect 30746 16895 30802 16904
rect 30656 16788 30708 16794
rect 30656 16730 30708 16736
rect 30564 16720 30616 16726
rect 30564 16662 30616 16668
rect 30472 16584 30524 16590
rect 30472 16526 30524 16532
rect 30380 16244 30432 16250
rect 30380 16186 30432 16192
rect 30196 15564 30248 15570
rect 30196 15506 30248 15512
rect 30484 15502 30512 16526
rect 30656 16448 30708 16454
rect 30656 16390 30708 16396
rect 30668 16182 30696 16390
rect 30656 16176 30708 16182
rect 30656 16118 30708 16124
rect 30288 15496 30340 15502
rect 30288 15438 30340 15444
rect 30472 15496 30524 15502
rect 30472 15438 30524 15444
rect 30196 14952 30248 14958
rect 30196 14894 30248 14900
rect 29748 14470 29960 14498
rect 30012 14544 30064 14550
rect 30012 14486 30064 14492
rect 29748 13462 29776 14470
rect 29828 14408 29880 14414
rect 29828 14350 29880 14356
rect 29920 14408 29972 14414
rect 30024 14362 30052 14486
rect 30208 14482 30236 14894
rect 30300 14770 30328 15438
rect 30472 15360 30524 15366
rect 30668 15314 30696 16118
rect 30748 15564 30800 15570
rect 30748 15506 30800 15512
rect 30472 15302 30524 15308
rect 30484 15094 30512 15302
rect 30576 15286 30696 15314
rect 30576 15094 30604 15286
rect 30472 15088 30524 15094
rect 30472 15030 30524 15036
rect 30564 15088 30616 15094
rect 30564 15030 30616 15036
rect 30300 14742 30420 14770
rect 30288 14612 30340 14618
rect 30288 14554 30340 14560
rect 30196 14476 30248 14482
rect 30196 14418 30248 14424
rect 29972 14356 30052 14362
rect 29920 14350 30052 14356
rect 29840 13462 29868 14350
rect 29932 14334 30052 14350
rect 30300 14346 30328 14554
rect 30392 14362 30420 14742
rect 30392 14346 30512 14362
rect 30288 14340 30340 14346
rect 30392 14340 30524 14346
rect 30392 14334 30472 14340
rect 30288 14282 30340 14288
rect 30472 14282 30524 14288
rect 30576 14278 30604 15030
rect 30760 14550 30788 15506
rect 30852 14634 30880 18634
rect 31036 17610 31064 19110
rect 31392 18692 31444 18698
rect 31392 18634 31444 18640
rect 31116 18624 31168 18630
rect 31116 18566 31168 18572
rect 31128 18222 31156 18566
rect 31116 18216 31168 18222
rect 31116 18158 31168 18164
rect 31116 18080 31168 18086
rect 31116 18022 31168 18028
rect 31024 17604 31076 17610
rect 31024 17546 31076 17552
rect 31022 17368 31078 17377
rect 31022 17303 31078 17312
rect 31036 17202 31064 17303
rect 31128 17202 31156 18022
rect 31404 17626 31432 18634
rect 31496 18154 31524 19314
rect 31680 18834 31708 19314
rect 31864 19306 32076 19334
rect 31668 18828 31720 18834
rect 31668 18770 31720 18776
rect 31484 18148 31536 18154
rect 31484 18090 31536 18096
rect 31680 17898 31708 18770
rect 31864 18329 31892 19306
rect 32128 18692 32180 18698
rect 32128 18634 32180 18640
rect 32140 18426 32168 18634
rect 32128 18420 32180 18426
rect 32128 18362 32180 18368
rect 31850 18320 31906 18329
rect 31850 18255 31906 18264
rect 31588 17870 31708 17898
rect 31588 17746 31616 17870
rect 31576 17740 31628 17746
rect 31576 17682 31628 17688
rect 31404 17610 31524 17626
rect 31404 17604 31536 17610
rect 31404 17598 31484 17604
rect 31484 17546 31536 17552
rect 31024 17196 31076 17202
rect 31024 17138 31076 17144
rect 31116 17196 31168 17202
rect 31116 17138 31168 17144
rect 31208 17196 31260 17202
rect 31208 17138 31260 17144
rect 31392 17196 31444 17202
rect 31392 17138 31444 17144
rect 31220 17066 31248 17138
rect 31208 17060 31260 17066
rect 31208 17002 31260 17008
rect 30932 16788 30984 16794
rect 30932 16730 30984 16736
rect 31024 16788 31076 16794
rect 31024 16730 31076 16736
rect 30944 14958 30972 16730
rect 31036 16697 31064 16730
rect 31022 16688 31078 16697
rect 31022 16623 31078 16632
rect 31220 16574 31248 17002
rect 31404 16726 31432 17138
rect 31392 16720 31444 16726
rect 31390 16688 31392 16697
rect 31444 16688 31446 16697
rect 31390 16623 31446 16632
rect 31022 16552 31078 16561
rect 31022 16487 31078 16496
rect 31128 16546 31248 16574
rect 31036 15910 31064 16487
rect 31128 16250 31156 16546
rect 31496 16522 31524 17546
rect 31668 17536 31720 17542
rect 31668 17478 31720 17484
rect 31680 17202 31708 17478
rect 31668 17196 31720 17202
rect 31668 17138 31720 17144
rect 31864 16998 31892 18255
rect 32232 17338 32260 19654
rect 33612 19378 33640 20334
rect 34072 20058 34100 21490
rect 34164 21146 34192 21490
rect 34336 21412 34388 21418
rect 34336 21354 34388 21360
rect 34152 21140 34204 21146
rect 34152 21082 34204 21088
rect 34348 21010 34376 21354
rect 34440 21146 34468 21490
rect 34428 21140 34480 21146
rect 34428 21082 34480 21088
rect 34336 21004 34388 21010
rect 34336 20946 34388 20952
rect 34532 20806 34560 21490
rect 34520 20800 34572 20806
rect 34520 20742 34572 20748
rect 34060 20052 34112 20058
rect 34060 19994 34112 20000
rect 34624 19854 34652 21966
rect 34704 21956 34756 21962
rect 34704 21898 34756 21904
rect 34716 21010 34744 21898
rect 34704 21004 34756 21010
rect 34704 20946 34756 20952
rect 34702 20904 34758 20913
rect 34702 20839 34758 20848
rect 34716 20806 34744 20839
rect 34704 20800 34756 20806
rect 34704 20742 34756 20748
rect 34716 20641 34744 20742
rect 34702 20632 34758 20641
rect 34808 20602 34836 22066
rect 35360 22030 35388 22374
rect 35348 22024 35400 22030
rect 35348 21966 35400 21972
rect 35072 21888 35124 21894
rect 35072 21830 35124 21836
rect 35164 21888 35216 21894
rect 35164 21830 35216 21836
rect 35348 21888 35400 21894
rect 35348 21830 35400 21836
rect 35084 21350 35112 21830
rect 35176 21554 35204 21830
rect 35164 21548 35216 21554
rect 35164 21490 35216 21496
rect 35072 21344 35124 21350
rect 35072 21286 35124 21292
rect 34934 21244 35242 21253
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21179 35242 21188
rect 35360 21146 35388 21830
rect 35452 21486 35480 23140
rect 35622 23080 35678 23089
rect 35622 23015 35624 23024
rect 35676 23015 35678 23024
rect 35820 23032 35848 23598
rect 36188 23225 36216 23598
rect 36174 23216 36230 23225
rect 36174 23151 36230 23160
rect 36280 23118 36308 24228
rect 36268 23112 36320 23118
rect 36174 23080 36230 23089
rect 35820 23004 36032 23032
rect 36268 23054 36320 23060
rect 36174 23015 36230 23024
rect 35624 22986 35676 22992
rect 35594 22876 35902 22885
rect 35594 22874 35600 22876
rect 35656 22874 35680 22876
rect 35736 22874 35760 22876
rect 35816 22874 35840 22876
rect 35896 22874 35902 22876
rect 35656 22822 35658 22874
rect 35838 22822 35840 22874
rect 35594 22820 35600 22822
rect 35656 22820 35680 22822
rect 35736 22820 35760 22822
rect 35816 22820 35840 22822
rect 35896 22820 35902 22822
rect 35594 22811 35902 22820
rect 36004 22778 36032 23004
rect 35992 22772 36044 22778
rect 35992 22714 36044 22720
rect 35808 22704 35860 22710
rect 35808 22646 35860 22652
rect 35622 22400 35678 22409
rect 35622 22335 35678 22344
rect 35636 22234 35664 22335
rect 35624 22228 35676 22234
rect 35624 22170 35676 22176
rect 35716 22228 35768 22234
rect 35716 22170 35768 22176
rect 35728 22030 35756 22170
rect 35820 22030 35848 22646
rect 35900 22568 35952 22574
rect 35898 22536 35900 22545
rect 35952 22536 35954 22545
rect 35898 22471 35954 22480
rect 36004 22234 36032 22714
rect 36084 22636 36136 22642
rect 36084 22578 36136 22584
rect 35992 22228 36044 22234
rect 35992 22170 36044 22176
rect 35716 22024 35768 22030
rect 35716 21966 35768 21972
rect 35808 22024 35860 22030
rect 35808 21966 35860 21972
rect 35594 21788 35902 21797
rect 35594 21786 35600 21788
rect 35656 21786 35680 21788
rect 35736 21786 35760 21788
rect 35816 21786 35840 21788
rect 35896 21786 35902 21788
rect 35656 21734 35658 21786
rect 35838 21734 35840 21786
rect 35594 21732 35600 21734
rect 35656 21732 35680 21734
rect 35736 21732 35760 21734
rect 35816 21732 35840 21734
rect 35896 21732 35902 21734
rect 35594 21723 35902 21732
rect 35440 21480 35492 21486
rect 35440 21422 35492 21428
rect 35900 21480 35952 21486
rect 35900 21422 35952 21428
rect 35164 21140 35216 21146
rect 35164 21082 35216 21088
rect 35348 21140 35400 21146
rect 35348 21082 35400 21088
rect 35176 20942 35204 21082
rect 35164 20936 35216 20942
rect 35164 20878 35216 20884
rect 35808 20936 35860 20942
rect 35912 20890 35940 21422
rect 36004 21332 36032 22170
rect 36096 21486 36124 22578
rect 36188 21622 36216 23015
rect 36372 22574 36400 24278
rect 36464 23118 36492 24534
rect 36634 24440 36690 24449
rect 36634 24375 36690 24384
rect 36544 24200 36596 24206
rect 36544 24142 36596 24148
rect 36556 23526 36584 24142
rect 36648 23798 36676 24375
rect 36740 24206 36768 25774
rect 36832 25362 36860 26862
rect 37188 26376 37240 26382
rect 37188 26318 37240 26324
rect 36912 25968 36964 25974
rect 36912 25910 36964 25916
rect 36820 25356 36872 25362
rect 36820 25298 36872 25304
rect 36820 25220 36872 25226
rect 36820 25162 36872 25168
rect 36832 24721 36860 25162
rect 36818 24712 36874 24721
rect 36818 24647 36874 24656
rect 36818 24304 36874 24313
rect 36818 24239 36820 24248
rect 36872 24239 36874 24248
rect 36820 24210 36872 24216
rect 36924 24206 36952 25910
rect 37200 25906 37228 26318
rect 37648 26036 37700 26042
rect 37648 25978 37700 25984
rect 37188 25900 37240 25906
rect 37188 25842 37240 25848
rect 37096 25356 37148 25362
rect 37096 25298 37148 25304
rect 37004 25288 37056 25294
rect 37002 25256 37004 25265
rect 37056 25256 37058 25265
rect 37002 25191 37058 25200
rect 37016 25158 37044 25191
rect 37004 25152 37056 25158
rect 37004 25094 37056 25100
rect 36728 24200 36780 24206
rect 36912 24200 36964 24206
rect 36728 24142 36780 24148
rect 36818 24168 36874 24177
rect 36912 24142 36964 24148
rect 37016 24138 37044 25094
rect 37108 24206 37136 25298
rect 37200 25294 37228 25842
rect 37464 25424 37516 25430
rect 37464 25366 37516 25372
rect 37188 25288 37240 25294
rect 37188 25230 37240 25236
rect 37476 24614 37504 25366
rect 37660 25226 37688 25978
rect 37740 25696 37792 25702
rect 37740 25638 37792 25644
rect 37752 25362 37780 25638
rect 37740 25356 37792 25362
rect 37740 25298 37792 25304
rect 37648 25220 37700 25226
rect 37648 25162 37700 25168
rect 37556 25152 37608 25158
rect 37556 25094 37608 25100
rect 37568 24818 37596 25094
rect 37556 24812 37608 24818
rect 37556 24754 37608 24760
rect 37464 24608 37516 24614
rect 37464 24550 37516 24556
rect 37738 24440 37794 24449
rect 37738 24375 37794 24384
rect 37096 24200 37148 24206
rect 37096 24142 37148 24148
rect 36818 24103 36874 24112
rect 37004 24132 37056 24138
rect 36832 23905 36860 24103
rect 37004 24074 37056 24080
rect 36818 23896 36874 23905
rect 36818 23831 36874 23840
rect 36832 23798 36860 23831
rect 36636 23792 36688 23798
rect 36636 23734 36688 23740
rect 36820 23792 36872 23798
rect 36820 23734 36872 23740
rect 36912 23656 36964 23662
rect 36912 23598 36964 23604
rect 36544 23520 36596 23526
rect 36544 23462 36596 23468
rect 36452 23112 36504 23118
rect 36452 23054 36504 23060
rect 36452 22636 36504 22642
rect 36556 22624 36584 23462
rect 36636 23112 36688 23118
rect 36636 23054 36688 23060
rect 36648 22642 36676 23054
rect 36820 22976 36872 22982
rect 36820 22918 36872 22924
rect 36504 22596 36584 22624
rect 36636 22636 36688 22642
rect 36452 22578 36504 22584
rect 36636 22578 36688 22584
rect 36360 22568 36412 22574
rect 36360 22510 36412 22516
rect 36372 22409 36400 22510
rect 36358 22400 36414 22409
rect 36358 22335 36414 22344
rect 36268 22228 36320 22234
rect 36268 22170 36320 22176
rect 36176 21616 36228 21622
rect 36176 21558 36228 21564
rect 36084 21480 36136 21486
rect 36084 21422 36136 21428
rect 36084 21344 36136 21350
rect 36004 21304 36084 21332
rect 36084 21286 36136 21292
rect 35860 20884 36032 20890
rect 35808 20878 36032 20884
rect 34702 20567 34758 20576
rect 34796 20596 34848 20602
rect 34796 20538 34848 20544
rect 34796 20460 34848 20466
rect 34796 20402 34848 20408
rect 34704 20392 34756 20398
rect 34704 20334 34756 20340
rect 34716 20058 34744 20334
rect 34808 20058 34836 20402
rect 35176 20398 35204 20878
rect 35820 20862 36032 20878
rect 35594 20700 35902 20709
rect 35594 20698 35600 20700
rect 35656 20698 35680 20700
rect 35736 20698 35760 20700
rect 35816 20698 35840 20700
rect 35896 20698 35902 20700
rect 35656 20646 35658 20698
rect 35838 20646 35840 20698
rect 35594 20644 35600 20646
rect 35656 20644 35680 20646
rect 35736 20644 35760 20646
rect 35816 20644 35840 20646
rect 35896 20644 35902 20646
rect 35594 20635 35902 20644
rect 35716 20460 35768 20466
rect 35716 20402 35768 20408
rect 35164 20392 35216 20398
rect 35164 20334 35216 20340
rect 35348 20392 35400 20398
rect 35348 20334 35400 20340
rect 34934 20156 35242 20165
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20091 35242 20100
rect 34704 20052 34756 20058
rect 34704 19994 34756 20000
rect 34796 20052 34848 20058
rect 34796 19994 34848 20000
rect 34808 19922 34928 19938
rect 34796 19916 34928 19922
rect 34848 19910 34928 19916
rect 34796 19858 34848 19864
rect 34520 19848 34572 19854
rect 34518 19816 34520 19825
rect 34612 19848 34664 19854
rect 34572 19816 34574 19825
rect 34244 19780 34296 19786
rect 34612 19790 34664 19796
rect 34704 19848 34756 19854
rect 34704 19790 34756 19796
rect 34518 19751 34574 19760
rect 34244 19722 34296 19728
rect 34256 19514 34284 19722
rect 34532 19530 34560 19751
rect 34612 19712 34664 19718
rect 34612 19654 34664 19660
rect 34244 19508 34296 19514
rect 34244 19450 34296 19456
rect 34348 19502 34560 19530
rect 33600 19372 33652 19378
rect 33600 19314 33652 19320
rect 32496 19168 32548 19174
rect 32496 19110 32548 19116
rect 32508 18290 32536 19110
rect 34348 18902 34376 19502
rect 34428 19372 34480 19378
rect 34428 19314 34480 19320
rect 34336 18896 34388 18902
rect 34336 18838 34388 18844
rect 34440 18850 34468 19314
rect 34520 19304 34572 19310
rect 34520 19246 34572 19252
rect 34532 18970 34560 19246
rect 34520 18964 34572 18970
rect 34520 18906 34572 18912
rect 34060 18828 34112 18834
rect 34440 18822 34560 18850
rect 34624 18834 34652 19654
rect 34716 19310 34744 19790
rect 34704 19304 34756 19310
rect 34704 19246 34756 19252
rect 34060 18770 34112 18776
rect 34072 18290 34100 18770
rect 32496 18284 32548 18290
rect 32496 18226 32548 18232
rect 34060 18284 34112 18290
rect 34060 18226 34112 18232
rect 33508 18216 33560 18222
rect 33508 18158 33560 18164
rect 32312 18148 32364 18154
rect 32312 18090 32364 18096
rect 32324 17542 32352 18090
rect 32496 18080 32548 18086
rect 32496 18022 32548 18028
rect 32312 17536 32364 17542
rect 32312 17478 32364 17484
rect 32220 17332 32272 17338
rect 32220 17274 32272 17280
rect 32128 17264 32180 17270
rect 32128 17206 32180 17212
rect 31760 16992 31812 16998
rect 31852 16992 31904 16998
rect 31760 16934 31812 16940
rect 31850 16960 31852 16969
rect 31904 16960 31906 16969
rect 31484 16516 31536 16522
rect 31484 16458 31536 16464
rect 31208 16448 31260 16454
rect 31208 16390 31260 16396
rect 31116 16244 31168 16250
rect 31116 16186 31168 16192
rect 31220 16114 31248 16390
rect 31772 16114 31800 16934
rect 31850 16895 31906 16904
rect 31208 16108 31260 16114
rect 31208 16050 31260 16056
rect 31760 16108 31812 16114
rect 31760 16050 31812 16056
rect 31024 15904 31076 15910
rect 31024 15846 31076 15852
rect 31036 15638 31064 15846
rect 31024 15632 31076 15638
rect 31024 15574 31076 15580
rect 32140 15570 32168 17206
rect 32128 15564 32180 15570
rect 32128 15506 32180 15512
rect 32140 15162 32168 15506
rect 32128 15156 32180 15162
rect 32128 15098 32180 15104
rect 30932 14952 30984 14958
rect 30932 14894 30984 14900
rect 30852 14606 31064 14634
rect 30748 14544 30800 14550
rect 30748 14486 30800 14492
rect 30932 14544 30984 14550
rect 30932 14486 30984 14492
rect 30944 14414 30972 14486
rect 30932 14408 30984 14414
rect 30932 14350 30984 14356
rect 30012 14272 30064 14278
rect 30012 14214 30064 14220
rect 30380 14272 30432 14278
rect 30380 14214 30432 14220
rect 30564 14272 30616 14278
rect 30564 14214 30616 14220
rect 30024 14090 30052 14214
rect 29932 14074 30052 14090
rect 29920 14068 30052 14074
rect 29972 14062 30052 14068
rect 29920 14010 29972 14016
rect 29736 13456 29788 13462
rect 29736 13398 29788 13404
rect 29828 13456 29880 13462
rect 29828 13398 29880 13404
rect 29736 13320 29788 13326
rect 29736 13262 29788 13268
rect 29644 13252 29696 13258
rect 29644 13194 29696 13200
rect 29000 12844 29052 12850
rect 29000 12786 29052 12792
rect 29368 12844 29420 12850
rect 29368 12786 29420 12792
rect 29644 12844 29696 12850
rect 29644 12786 29696 12792
rect 29012 12442 29040 12786
rect 29184 12776 29236 12782
rect 29184 12718 29236 12724
rect 29000 12436 29052 12442
rect 29000 12378 29052 12384
rect 28724 12232 28776 12238
rect 28908 12232 28960 12238
rect 28724 12174 28776 12180
rect 28828 12192 28908 12220
rect 28736 11558 28764 12174
rect 28828 11762 28856 12192
rect 28908 12174 28960 12180
rect 28816 11756 28868 11762
rect 28816 11698 28868 11704
rect 28724 11552 28776 11558
rect 28724 11494 28776 11500
rect 28540 11280 28592 11286
rect 28540 11222 28592 11228
rect 28448 10804 28500 10810
rect 28448 10746 28500 10752
rect 28552 10674 28580 11222
rect 27988 10668 28040 10674
rect 27988 10610 28040 10616
rect 28356 10668 28408 10674
rect 28356 10610 28408 10616
rect 28540 10668 28592 10674
rect 28540 10610 28592 10616
rect 27712 10260 27764 10266
rect 27712 10202 27764 10208
rect 27620 10192 27672 10198
rect 27620 10134 27672 10140
rect 27724 10062 27752 10202
rect 27344 10056 27396 10062
rect 27344 9998 27396 10004
rect 27712 10056 27764 10062
rect 27712 9998 27764 10004
rect 27356 8838 27384 9998
rect 27724 9722 27752 9998
rect 27712 9716 27764 9722
rect 27712 9658 27764 9664
rect 27620 8968 27672 8974
rect 27620 8910 27672 8916
rect 27344 8832 27396 8838
rect 27344 8774 27396 8780
rect 27632 8430 27660 8910
rect 27068 8424 27120 8430
rect 27068 8366 27120 8372
rect 27620 8424 27672 8430
rect 27620 8366 27672 8372
rect 26976 8288 27028 8294
rect 26976 8230 27028 8236
rect 26792 7948 26844 7954
rect 26792 7890 26844 7896
rect 26240 7336 26292 7342
rect 26240 7278 26292 7284
rect 26608 7336 26660 7342
rect 26608 7278 26660 7284
rect 26252 7002 26280 7278
rect 26804 7274 26832 7890
rect 26988 7886 27016 8230
rect 27080 7886 27108 8366
rect 27344 7948 27396 7954
rect 27344 7890 27396 7896
rect 26976 7880 27028 7886
rect 26976 7822 27028 7828
rect 27068 7880 27120 7886
rect 27068 7822 27120 7828
rect 27252 7540 27304 7546
rect 27252 7482 27304 7488
rect 26792 7268 26844 7274
rect 26792 7210 26844 7216
rect 26240 6996 26292 7002
rect 26240 6938 26292 6944
rect 26252 5370 26280 6938
rect 27264 6798 27292 7482
rect 27356 6798 27384 7890
rect 27620 7404 27672 7410
rect 27620 7346 27672 7352
rect 27252 6792 27304 6798
rect 27252 6734 27304 6740
rect 27344 6792 27396 6798
rect 27344 6734 27396 6740
rect 27436 6792 27488 6798
rect 27632 6780 27660 7346
rect 27488 6752 27660 6780
rect 27436 6734 27488 6740
rect 27436 6316 27488 6322
rect 27436 6258 27488 6264
rect 27448 5914 27476 6258
rect 27436 5908 27488 5914
rect 27436 5850 27488 5856
rect 27620 5636 27672 5642
rect 27620 5578 27672 5584
rect 27632 5370 27660 5578
rect 26240 5364 26292 5370
rect 26240 5306 26292 5312
rect 27620 5364 27672 5370
rect 27620 5306 27672 5312
rect 27724 4826 27752 9658
rect 28000 9382 28028 10610
rect 28724 10532 28776 10538
rect 28724 10474 28776 10480
rect 28736 9994 28764 10474
rect 28724 9988 28776 9994
rect 28724 9930 28776 9936
rect 28736 9586 28764 9930
rect 28724 9580 28776 9586
rect 28724 9522 28776 9528
rect 27988 9376 28040 9382
rect 27988 9318 28040 9324
rect 28080 9172 28132 9178
rect 28080 9114 28132 9120
rect 27804 9104 27856 9110
rect 27804 9046 27856 9052
rect 27816 8906 27844 9046
rect 27804 8900 27856 8906
rect 27804 8842 27856 8848
rect 27816 8022 27844 8842
rect 28092 8362 28120 9114
rect 28540 9036 28592 9042
rect 28540 8978 28592 8984
rect 28552 8430 28580 8978
rect 28632 8968 28684 8974
rect 28632 8910 28684 8916
rect 28540 8424 28592 8430
rect 28540 8366 28592 8372
rect 28080 8356 28132 8362
rect 28080 8298 28132 8304
rect 27804 8016 27856 8022
rect 27804 7958 27856 7964
rect 27816 6254 27844 7958
rect 28092 7886 28120 8298
rect 28448 8288 28500 8294
rect 28448 8230 28500 8236
rect 28460 8022 28488 8230
rect 28448 8016 28500 8022
rect 28448 7958 28500 7964
rect 28552 7954 28580 8366
rect 28644 8294 28672 8910
rect 28632 8288 28684 8294
rect 28632 8230 28684 8236
rect 28644 8090 28672 8230
rect 28632 8084 28684 8090
rect 28632 8026 28684 8032
rect 28540 7948 28592 7954
rect 28540 7890 28592 7896
rect 28080 7880 28132 7886
rect 28080 7822 28132 7828
rect 28552 7410 28580 7890
rect 28540 7404 28592 7410
rect 28540 7346 28592 7352
rect 28172 7200 28224 7206
rect 28172 7142 28224 7148
rect 27804 6248 27856 6254
rect 27804 6190 27856 6196
rect 27816 5556 27844 6190
rect 27896 6112 27948 6118
rect 27896 6054 27948 6060
rect 27908 5710 27936 6054
rect 27896 5704 27948 5710
rect 27896 5646 27948 5652
rect 27896 5568 27948 5574
rect 27816 5528 27896 5556
rect 27896 5510 27948 5516
rect 28080 5568 28132 5574
rect 28080 5510 28132 5516
rect 27804 5364 27856 5370
rect 27804 5306 27856 5312
rect 26148 4820 26200 4826
rect 26148 4762 26200 4768
rect 27712 4820 27764 4826
rect 27712 4762 27764 4768
rect 27724 4622 27752 4762
rect 27712 4616 27764 4622
rect 27712 4558 27764 4564
rect 27816 4554 27844 5306
rect 26056 4548 26108 4554
rect 26056 4490 26108 4496
rect 27804 4548 27856 4554
rect 27804 4490 27856 4496
rect 26068 4214 26096 4490
rect 27816 4214 27844 4490
rect 26056 4208 26108 4214
rect 26056 4150 26108 4156
rect 27804 4208 27856 4214
rect 27804 4150 27856 4156
rect 25320 4140 25372 4146
rect 25320 4082 25372 4088
rect 25332 3738 25360 4082
rect 25964 3936 26016 3942
rect 25964 3878 26016 3884
rect 25320 3732 25372 3738
rect 25320 3674 25372 3680
rect 25780 3732 25832 3738
rect 25780 3674 25832 3680
rect 23940 3596 23992 3602
rect 23940 3538 23992 3544
rect 24768 3596 24820 3602
rect 24768 3538 24820 3544
rect 23756 3188 23808 3194
rect 23756 3130 23808 3136
rect 23952 3058 23980 3538
rect 25792 3534 25820 3674
rect 25976 3534 26004 3878
rect 25688 3528 25740 3534
rect 25688 3470 25740 3476
rect 25780 3528 25832 3534
rect 25780 3470 25832 3476
rect 25964 3528 26016 3534
rect 25964 3470 26016 3476
rect 25700 3194 25728 3470
rect 25688 3188 25740 3194
rect 25688 3130 25740 3136
rect 26068 3126 26096 4150
rect 26516 4140 26568 4146
rect 26516 4082 26568 4088
rect 26528 3738 26556 4082
rect 26516 3732 26568 3738
rect 26516 3674 26568 3680
rect 27816 3466 27844 4150
rect 27908 3738 27936 5510
rect 28092 5302 28120 5510
rect 28184 5370 28212 7142
rect 28552 7002 28580 7346
rect 28540 6996 28592 7002
rect 28540 6938 28592 6944
rect 28644 6254 28672 8026
rect 28736 7886 28764 9522
rect 28828 9518 28856 11698
rect 29196 11558 29224 12718
rect 29276 11688 29328 11694
rect 29274 11656 29276 11665
rect 29328 11656 29330 11665
rect 29380 11642 29408 12786
rect 29552 12708 29604 12714
rect 29552 12650 29604 12656
rect 29460 12096 29512 12102
rect 29460 12038 29512 12044
rect 29330 11614 29408 11642
rect 29274 11591 29330 11600
rect 29184 11552 29236 11558
rect 29184 11494 29236 11500
rect 28908 11348 28960 11354
rect 28908 11290 28960 11296
rect 28920 10674 28948 11290
rect 29090 11248 29146 11257
rect 29090 11183 29146 11192
rect 29276 11212 29328 11218
rect 29104 11150 29132 11183
rect 29276 11154 29328 11160
rect 29000 11144 29052 11150
rect 29000 11086 29052 11092
rect 29092 11144 29144 11150
rect 29092 11086 29144 11092
rect 29012 10985 29040 11086
rect 28998 10976 29054 10985
rect 28998 10911 29054 10920
rect 28908 10668 28960 10674
rect 28908 10610 28960 10616
rect 29184 10668 29236 10674
rect 29184 10610 29236 10616
rect 29092 10600 29144 10606
rect 29092 10542 29144 10548
rect 29104 9994 29132 10542
rect 29000 9988 29052 9994
rect 29000 9930 29052 9936
rect 29092 9988 29144 9994
rect 29092 9930 29144 9936
rect 29012 9654 29040 9930
rect 29000 9648 29052 9654
rect 29000 9590 29052 9596
rect 28816 9512 28868 9518
rect 28816 9454 28868 9460
rect 28816 9376 28868 9382
rect 28816 9318 28868 9324
rect 28828 9178 28856 9318
rect 28816 9172 28868 9178
rect 28816 9114 28868 9120
rect 29012 8634 29040 9590
rect 29092 9580 29144 9586
rect 29196 9568 29224 10610
rect 29288 9722 29316 11154
rect 29380 10266 29408 11614
rect 29472 10674 29500 12038
rect 29564 11898 29592 12650
rect 29656 11937 29684 12786
rect 29748 12442 29776 13262
rect 29736 12436 29788 12442
rect 29736 12378 29788 12384
rect 29642 11928 29698 11937
rect 29552 11892 29604 11898
rect 29642 11863 29698 11872
rect 29552 11834 29604 11840
rect 29552 11756 29604 11762
rect 29552 11698 29604 11704
rect 29564 11082 29592 11698
rect 29656 11626 29684 11863
rect 29734 11792 29790 11801
rect 29734 11727 29736 11736
rect 29788 11727 29790 11736
rect 29736 11698 29788 11704
rect 29644 11620 29696 11626
rect 29644 11562 29696 11568
rect 29840 11354 29868 13398
rect 30024 13394 30052 14062
rect 30392 14006 30420 14214
rect 30380 14000 30432 14006
rect 30380 13942 30432 13948
rect 30472 13728 30524 13734
rect 30472 13670 30524 13676
rect 30012 13388 30064 13394
rect 30012 13330 30064 13336
rect 30024 12986 30052 13330
rect 30484 13326 30512 13670
rect 30944 13326 30972 14350
rect 31036 14006 31064 14606
rect 31668 14544 31720 14550
rect 31668 14486 31720 14492
rect 31024 14000 31076 14006
rect 31024 13942 31076 13948
rect 31036 13870 31064 13942
rect 31680 13938 31708 14486
rect 31668 13932 31720 13938
rect 31668 13874 31720 13880
rect 31024 13864 31076 13870
rect 31024 13806 31076 13812
rect 32324 13326 32352 17478
rect 32402 17368 32458 17377
rect 32508 17338 32536 18022
rect 32402 17303 32404 17312
rect 32456 17303 32458 17312
rect 32496 17332 32548 17338
rect 32404 17274 32456 17280
rect 32496 17274 32548 17280
rect 33520 17202 33548 18158
rect 33784 17536 33836 17542
rect 33784 17478 33836 17484
rect 33796 17270 33824 17478
rect 33784 17264 33836 17270
rect 33784 17206 33836 17212
rect 33508 17196 33560 17202
rect 33508 17138 33560 17144
rect 33520 16658 33548 17138
rect 34072 16726 34100 18226
rect 34532 17678 34560 18822
rect 34612 18828 34664 18834
rect 34612 18770 34664 18776
rect 34716 18766 34744 19246
rect 34900 19174 34928 19910
rect 35360 19854 35388 20334
rect 35440 19984 35492 19990
rect 35440 19926 35492 19932
rect 35348 19848 35400 19854
rect 35348 19790 35400 19796
rect 35348 19440 35400 19446
rect 35348 19382 35400 19388
rect 34888 19168 34940 19174
rect 34794 19136 34850 19145
rect 34888 19110 34940 19116
rect 34794 19071 34850 19080
rect 34808 18766 34836 19071
rect 34934 19068 35242 19077
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 19003 35242 19012
rect 34704 18760 34756 18766
rect 34704 18702 34756 18708
rect 34796 18760 34848 18766
rect 34796 18702 34848 18708
rect 34934 17980 35242 17989
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17915 35242 17924
rect 34704 17876 34756 17882
rect 34704 17818 34756 17824
rect 34520 17672 34572 17678
rect 34520 17614 34572 17620
rect 34244 17264 34296 17270
rect 34244 17206 34296 17212
rect 34256 16794 34284 17206
rect 34520 17128 34572 17134
rect 34520 17070 34572 17076
rect 34244 16788 34296 16794
rect 34244 16730 34296 16736
rect 34060 16720 34112 16726
rect 34060 16662 34112 16668
rect 33508 16652 33560 16658
rect 33508 16594 33560 16600
rect 32772 16516 32824 16522
rect 32772 16458 32824 16464
rect 32784 16250 32812 16458
rect 32772 16244 32824 16250
rect 32772 16186 32824 16192
rect 33520 16182 33548 16594
rect 33508 16176 33560 16182
rect 33508 16118 33560 16124
rect 33520 15570 33548 16118
rect 34072 15910 34100 16662
rect 34060 15904 34112 15910
rect 34060 15846 34112 15852
rect 34532 15706 34560 17070
rect 34520 15700 34572 15706
rect 34520 15642 34572 15648
rect 33508 15564 33560 15570
rect 33508 15506 33560 15512
rect 32588 15496 32640 15502
rect 32588 15438 32640 15444
rect 32600 14482 32628 15438
rect 32772 15428 32824 15434
rect 32772 15370 32824 15376
rect 32588 14476 32640 14482
rect 32588 14418 32640 14424
rect 32784 14006 32812 15370
rect 34244 15088 34296 15094
rect 34244 15030 34296 15036
rect 32864 14340 32916 14346
rect 32864 14282 32916 14288
rect 32876 14074 32904 14282
rect 32864 14068 32916 14074
rect 32864 14010 32916 14016
rect 34256 14006 34284 15030
rect 34336 14884 34388 14890
rect 34336 14826 34388 14832
rect 34348 14618 34376 14826
rect 34336 14612 34388 14618
rect 34336 14554 34388 14560
rect 34348 14074 34376 14554
rect 34336 14068 34388 14074
rect 34336 14010 34388 14016
rect 32772 14000 32824 14006
rect 32772 13942 32824 13948
rect 34244 14000 34296 14006
rect 34244 13942 34296 13948
rect 32588 13932 32640 13938
rect 32588 13874 32640 13880
rect 30472 13320 30524 13326
rect 30472 13262 30524 13268
rect 30932 13320 30984 13326
rect 30932 13262 30984 13268
rect 31116 13320 31168 13326
rect 31116 13262 31168 13268
rect 32312 13320 32364 13326
rect 32312 13262 32364 13268
rect 30380 13184 30432 13190
rect 30380 13126 30432 13132
rect 30012 12980 30064 12986
rect 30012 12922 30064 12928
rect 30288 12776 30340 12782
rect 30288 12718 30340 12724
rect 29920 12164 29972 12170
rect 29920 12106 29972 12112
rect 29828 11348 29880 11354
rect 29828 11290 29880 11296
rect 29932 11286 29960 12106
rect 30300 12102 30328 12718
rect 30392 12238 30420 13126
rect 31128 12986 31156 13262
rect 32600 13258 32628 13874
rect 32784 13802 32812 13942
rect 34532 13938 34560 15642
rect 34716 14822 34744 17818
rect 34888 17672 34940 17678
rect 34888 17614 34940 17620
rect 35072 17672 35124 17678
rect 35072 17614 35124 17620
rect 35256 17672 35308 17678
rect 35256 17614 35308 17620
rect 34900 17066 34928 17614
rect 35084 17320 35112 17614
rect 35268 17542 35296 17614
rect 35256 17536 35308 17542
rect 35256 17478 35308 17484
rect 35164 17332 35216 17338
rect 35084 17292 35164 17320
rect 35164 17274 35216 17280
rect 35268 17134 35296 17478
rect 35256 17128 35308 17134
rect 35256 17070 35308 17076
rect 34888 17060 34940 17066
rect 34808 17020 34888 17048
rect 34808 16658 34836 17020
rect 34888 17002 34940 17008
rect 34934 16892 35242 16901
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16827 35242 16836
rect 34796 16652 34848 16658
rect 34796 16594 34848 16600
rect 35256 16652 35308 16658
rect 35256 16594 35308 16600
rect 35164 16584 35216 16590
rect 35164 16526 35216 16532
rect 35176 16454 35204 16526
rect 34888 16448 34940 16454
rect 34888 16390 34940 16396
rect 35164 16448 35216 16454
rect 35164 16390 35216 16396
rect 34900 16046 34928 16390
rect 35268 16250 35296 16594
rect 35360 16522 35388 19382
rect 35452 19310 35480 19926
rect 35728 19854 35756 20402
rect 35716 19848 35768 19854
rect 35622 19816 35678 19825
rect 35716 19790 35768 19796
rect 35622 19751 35624 19760
rect 35676 19751 35678 19760
rect 35624 19722 35676 19728
rect 35594 19612 35902 19621
rect 35594 19610 35600 19612
rect 35656 19610 35680 19612
rect 35736 19610 35760 19612
rect 35816 19610 35840 19612
rect 35896 19610 35902 19612
rect 35656 19558 35658 19610
rect 35838 19558 35840 19610
rect 35594 19556 35600 19558
rect 35656 19556 35680 19558
rect 35736 19556 35760 19558
rect 35816 19556 35840 19558
rect 35896 19556 35902 19558
rect 35594 19547 35902 19556
rect 35440 19304 35492 19310
rect 35440 19246 35492 19252
rect 36004 19258 36032 20862
rect 36096 19854 36124 21286
rect 36280 21010 36308 22170
rect 36372 21162 36400 22335
rect 36464 22234 36492 22578
rect 36452 22228 36504 22234
rect 36452 22170 36504 22176
rect 36372 21134 36492 21162
rect 36268 21004 36320 21010
rect 36268 20946 36320 20952
rect 36360 21004 36412 21010
rect 36360 20946 36412 20952
rect 36372 20913 36400 20946
rect 36358 20904 36414 20913
rect 36358 20839 36414 20848
rect 36464 20602 36492 21134
rect 36452 20596 36504 20602
rect 36452 20538 36504 20544
rect 36268 20460 36320 20466
rect 36268 20402 36320 20408
rect 36280 19938 36308 20402
rect 36464 20058 36492 20538
rect 36648 20058 36676 22578
rect 36832 22574 36860 22918
rect 36820 22568 36872 22574
rect 36726 22536 36782 22545
rect 36820 22510 36872 22516
rect 36726 22471 36782 22480
rect 36740 21690 36768 22471
rect 36728 21684 36780 21690
rect 36728 21626 36780 21632
rect 36740 21146 36768 21626
rect 36728 21140 36780 21146
rect 36728 21082 36780 21088
rect 36818 20904 36874 20913
rect 36818 20839 36820 20848
rect 36872 20839 36874 20848
rect 36820 20810 36872 20816
rect 36452 20052 36504 20058
rect 36452 19994 36504 20000
rect 36636 20052 36688 20058
rect 36636 19994 36688 20000
rect 36188 19910 36308 19938
rect 36084 19848 36136 19854
rect 36084 19790 36136 19796
rect 36084 19712 36136 19718
rect 36084 19654 36136 19660
rect 36096 19378 36124 19654
rect 36084 19372 36136 19378
rect 36084 19314 36136 19320
rect 35532 19236 35584 19242
rect 36004 19230 36124 19258
rect 35532 19178 35584 19184
rect 35544 18970 35572 19178
rect 35532 18964 35584 18970
rect 35532 18906 35584 18912
rect 35594 18524 35902 18533
rect 35594 18522 35600 18524
rect 35656 18522 35680 18524
rect 35736 18522 35760 18524
rect 35816 18522 35840 18524
rect 35896 18522 35902 18524
rect 35656 18470 35658 18522
rect 35838 18470 35840 18522
rect 35594 18468 35600 18470
rect 35656 18468 35680 18470
rect 35736 18468 35760 18470
rect 35816 18468 35840 18470
rect 35896 18468 35902 18470
rect 35594 18459 35902 18468
rect 35992 18216 36044 18222
rect 35992 18158 36044 18164
rect 36004 17882 36032 18158
rect 35992 17876 36044 17882
rect 35992 17818 36044 17824
rect 35992 17604 36044 17610
rect 35992 17546 36044 17552
rect 35594 17436 35902 17445
rect 35594 17434 35600 17436
rect 35656 17434 35680 17436
rect 35736 17434 35760 17436
rect 35816 17434 35840 17436
rect 35896 17434 35902 17436
rect 35656 17382 35658 17434
rect 35838 17382 35840 17434
rect 35594 17380 35600 17382
rect 35656 17380 35680 17382
rect 35736 17380 35760 17382
rect 35816 17380 35840 17382
rect 35896 17380 35902 17382
rect 35594 17371 35902 17380
rect 35716 17196 35768 17202
rect 35716 17138 35768 17144
rect 35900 17196 35952 17202
rect 35900 17138 35952 17144
rect 35532 17128 35584 17134
rect 35532 17070 35584 17076
rect 35440 16584 35492 16590
rect 35438 16552 35440 16561
rect 35544 16572 35572 17070
rect 35728 16590 35756 17138
rect 35912 16998 35940 17138
rect 35900 16992 35952 16998
rect 35900 16934 35952 16940
rect 35808 16788 35860 16794
rect 35808 16730 35860 16736
rect 35820 16697 35848 16730
rect 35806 16688 35862 16697
rect 36004 16658 36032 17546
rect 36096 17338 36124 19230
rect 36188 17814 36216 19910
rect 36924 19854 36952 23598
rect 37464 23180 37516 23186
rect 37464 23122 37516 23128
rect 37476 22098 37504 23122
rect 37556 22636 37608 22642
rect 37556 22578 37608 22584
rect 37464 22092 37516 22098
rect 37464 22034 37516 22040
rect 37280 21956 37332 21962
rect 37280 21898 37332 21904
rect 37292 21622 37320 21898
rect 37280 21616 37332 21622
rect 37280 21558 37332 21564
rect 37188 20256 37240 20262
rect 37188 20198 37240 20204
rect 36912 19848 36964 19854
rect 36912 19790 36964 19796
rect 36268 19780 36320 19786
rect 36268 19722 36320 19728
rect 36452 19780 36504 19786
rect 36452 19722 36504 19728
rect 36280 19514 36308 19722
rect 36268 19508 36320 19514
rect 36268 19450 36320 19456
rect 36176 17808 36228 17814
rect 36176 17750 36228 17756
rect 36176 17672 36228 17678
rect 36176 17614 36228 17620
rect 36084 17332 36136 17338
rect 36084 17274 36136 17280
rect 36084 17196 36136 17202
rect 36084 17138 36136 17144
rect 36096 16697 36124 17138
rect 36188 17066 36216 17614
rect 36176 17060 36228 17066
rect 36176 17002 36228 17008
rect 36082 16688 36138 16697
rect 35806 16623 35862 16632
rect 35992 16652 36044 16658
rect 36082 16623 36138 16632
rect 35992 16594 36044 16600
rect 35492 16552 35572 16572
rect 35494 16544 35572 16552
rect 35716 16584 35768 16590
rect 35348 16516 35400 16522
rect 35768 16532 36032 16538
rect 35716 16526 36032 16532
rect 35728 16522 36032 16526
rect 35728 16516 36044 16522
rect 35728 16510 35992 16516
rect 35438 16487 35494 16496
rect 35348 16458 35400 16464
rect 35256 16244 35308 16250
rect 35256 16186 35308 16192
rect 35360 16182 35388 16458
rect 35348 16176 35400 16182
rect 35348 16118 35400 16124
rect 34888 16040 34940 16046
rect 34888 15982 34940 15988
rect 34934 15804 35242 15813
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15739 35242 15748
rect 34704 14816 34756 14822
rect 34704 14758 34756 14764
rect 34934 14716 35242 14725
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14651 35242 14660
rect 34704 14476 34756 14482
rect 34704 14418 34756 14424
rect 35256 14476 35308 14482
rect 35256 14418 35308 14424
rect 34520 13932 34572 13938
rect 34520 13874 34572 13880
rect 33508 13864 33560 13870
rect 33508 13806 33560 13812
rect 33692 13864 33744 13870
rect 33692 13806 33744 13812
rect 32772 13796 32824 13802
rect 32772 13738 32824 13744
rect 32784 13530 32812 13738
rect 32772 13524 32824 13530
rect 32772 13466 32824 13472
rect 33324 13320 33376 13326
rect 33324 13262 33376 13268
rect 32588 13252 32640 13258
rect 32588 13194 32640 13200
rect 31668 13184 31720 13190
rect 31668 13126 31720 13132
rect 31116 12980 31168 12986
rect 31116 12922 31168 12928
rect 30472 12640 30524 12646
rect 30472 12582 30524 12588
rect 30484 12238 30512 12582
rect 31680 12442 31708 13126
rect 32220 12980 32272 12986
rect 32220 12922 32272 12928
rect 33048 12980 33100 12986
rect 33048 12922 33100 12928
rect 31668 12436 31720 12442
rect 31668 12378 31720 12384
rect 30380 12232 30432 12238
rect 30380 12174 30432 12180
rect 30472 12232 30524 12238
rect 30472 12174 30524 12180
rect 30564 12232 30616 12238
rect 30564 12174 30616 12180
rect 31484 12232 31536 12238
rect 31484 12174 31536 12180
rect 31760 12232 31812 12238
rect 32232 12209 32260 12922
rect 32588 12844 32640 12850
rect 32588 12786 32640 12792
rect 32600 12442 32628 12786
rect 33060 12714 33088 12922
rect 33140 12776 33192 12782
rect 33140 12718 33192 12724
rect 33048 12708 33100 12714
rect 33048 12650 33100 12656
rect 32588 12436 32640 12442
rect 32588 12378 32640 12384
rect 32600 12345 32628 12378
rect 32680 12368 32732 12374
rect 32586 12336 32642 12345
rect 32680 12310 32732 12316
rect 32586 12271 32642 12280
rect 31760 12174 31812 12180
rect 32218 12200 32274 12209
rect 30288 12096 30340 12102
rect 30288 12038 30340 12044
rect 30392 11830 30420 12174
rect 30380 11824 30432 11830
rect 30380 11766 30432 11772
rect 30196 11756 30248 11762
rect 30196 11698 30248 11704
rect 29920 11280 29972 11286
rect 29920 11222 29972 11228
rect 29552 11076 29604 11082
rect 29552 11018 29604 11024
rect 29564 10810 29592 11018
rect 30208 10810 30236 11698
rect 30392 11286 30420 11766
rect 30472 11552 30524 11558
rect 30472 11494 30524 11500
rect 30380 11280 30432 11286
rect 30380 11222 30432 11228
rect 30484 11150 30512 11494
rect 30576 11354 30604 12174
rect 31024 12164 31076 12170
rect 31024 12106 31076 12112
rect 31036 11830 31064 12106
rect 31024 11824 31076 11830
rect 31024 11766 31076 11772
rect 31116 11824 31168 11830
rect 31116 11766 31168 11772
rect 30748 11688 30800 11694
rect 30748 11630 30800 11636
rect 30564 11348 30616 11354
rect 30564 11290 30616 11296
rect 30472 11144 30524 11150
rect 30472 11086 30524 11092
rect 29552 10804 29604 10810
rect 29552 10746 29604 10752
rect 30196 10804 30248 10810
rect 30196 10746 30248 10752
rect 30760 10742 30788 11630
rect 30932 11552 30984 11558
rect 30932 11494 30984 11500
rect 30944 11257 30972 11494
rect 30930 11248 30986 11257
rect 30930 11183 30986 11192
rect 30748 10736 30800 10742
rect 30748 10678 30800 10684
rect 29460 10668 29512 10674
rect 29460 10610 29512 10616
rect 30380 10668 30432 10674
rect 30380 10610 30432 10616
rect 29460 10464 29512 10470
rect 29460 10406 29512 10412
rect 29472 10266 29500 10406
rect 29368 10260 29420 10266
rect 29368 10202 29420 10208
rect 29460 10260 29512 10266
rect 29460 10202 29512 10208
rect 30392 10130 30420 10610
rect 30472 10464 30524 10470
rect 30472 10406 30524 10412
rect 30484 10266 30512 10406
rect 30944 10266 30972 11183
rect 31036 10985 31064 11766
rect 31128 11218 31156 11766
rect 31496 11626 31524 12174
rect 31484 11620 31536 11626
rect 31484 11562 31536 11568
rect 31116 11212 31168 11218
rect 31116 11154 31168 11160
rect 31022 10976 31078 10985
rect 31022 10911 31078 10920
rect 31036 10742 31064 10911
rect 31772 10810 31800 12174
rect 32218 12135 32274 12144
rect 31760 10804 31812 10810
rect 31760 10746 31812 10752
rect 31024 10736 31076 10742
rect 31024 10678 31076 10684
rect 31024 10600 31076 10606
rect 31208 10600 31260 10606
rect 31076 10548 31156 10554
rect 31024 10542 31156 10548
rect 31208 10542 31260 10548
rect 31036 10526 31156 10542
rect 30472 10260 30524 10266
rect 30472 10202 30524 10208
rect 30932 10260 30984 10266
rect 30932 10202 30984 10208
rect 30484 10130 30512 10202
rect 31128 10146 31156 10526
rect 31220 10266 31248 10542
rect 31760 10532 31812 10538
rect 31760 10474 31812 10480
rect 31208 10260 31260 10266
rect 31208 10202 31260 10208
rect 31300 10192 31352 10198
rect 31128 10140 31300 10146
rect 31128 10134 31352 10140
rect 30380 10124 30432 10130
rect 30380 10066 30432 10072
rect 30472 10124 30524 10130
rect 31128 10118 31340 10134
rect 31484 10124 31536 10130
rect 30472 10066 30524 10072
rect 31484 10066 31536 10072
rect 30392 9722 30420 10066
rect 31208 10056 31260 10062
rect 31208 9998 31260 10004
rect 29276 9716 29328 9722
rect 29276 9658 29328 9664
rect 30380 9716 30432 9722
rect 30380 9658 30432 9664
rect 29144 9540 29224 9568
rect 29092 9522 29144 9528
rect 29104 9178 29132 9522
rect 31220 9382 31248 9998
rect 31496 9518 31524 10066
rect 31484 9512 31536 9518
rect 31484 9454 31536 9460
rect 31208 9376 31260 9382
rect 31208 9318 31260 9324
rect 29092 9172 29144 9178
rect 29092 9114 29144 9120
rect 29000 8628 29052 8634
rect 29000 8570 29052 8576
rect 29104 8090 29132 9114
rect 31496 8634 31524 9454
rect 31772 9058 31800 10474
rect 32232 10266 32260 12135
rect 32588 12096 32640 12102
rect 32588 12038 32640 12044
rect 32496 11892 32548 11898
rect 32496 11834 32548 11840
rect 32312 11756 32364 11762
rect 32364 11716 32444 11744
rect 32312 11698 32364 11704
rect 32312 11212 32364 11218
rect 32312 11154 32364 11160
rect 32324 10577 32352 11154
rect 32416 10713 32444 11716
rect 32508 11150 32536 11834
rect 32600 11762 32628 12038
rect 32588 11756 32640 11762
rect 32588 11698 32640 11704
rect 32692 11626 32720 12310
rect 33060 12238 33088 12650
rect 33152 12442 33180 12718
rect 33232 12640 33284 12646
rect 33232 12582 33284 12588
rect 33140 12436 33192 12442
rect 33140 12378 33192 12384
rect 33048 12232 33100 12238
rect 32968 12192 33048 12220
rect 32772 11756 32824 11762
rect 32772 11698 32824 11704
rect 32864 11756 32916 11762
rect 32864 11698 32916 11704
rect 32680 11620 32732 11626
rect 32680 11562 32732 11568
rect 32496 11144 32548 11150
rect 32496 11086 32548 11092
rect 32692 10810 32720 11562
rect 32784 10810 32812 11698
rect 32876 11286 32904 11698
rect 32864 11280 32916 11286
rect 32864 11222 32916 11228
rect 32680 10804 32732 10810
rect 32680 10746 32732 10752
rect 32772 10804 32824 10810
rect 32772 10746 32824 10752
rect 32402 10704 32458 10713
rect 32402 10639 32458 10648
rect 32588 10668 32640 10674
rect 32310 10568 32366 10577
rect 32310 10503 32366 10512
rect 32324 10470 32352 10503
rect 32312 10464 32364 10470
rect 32312 10406 32364 10412
rect 32220 10260 32272 10266
rect 32220 10202 32272 10208
rect 32128 10192 32180 10198
rect 31850 10160 31906 10169
rect 32128 10134 32180 10140
rect 32310 10160 32366 10169
rect 31850 10095 31906 10104
rect 31864 9450 31892 10095
rect 31944 10056 31996 10062
rect 31944 9998 31996 10004
rect 31956 9450 31984 9998
rect 32036 9920 32088 9926
rect 32036 9862 32088 9868
rect 32048 9654 32076 9862
rect 32036 9648 32088 9654
rect 32036 9590 32088 9596
rect 32140 9586 32168 10134
rect 32310 10095 32312 10104
rect 32364 10095 32366 10104
rect 32312 10066 32364 10072
rect 32312 9988 32364 9994
rect 32312 9930 32364 9936
rect 32128 9580 32180 9586
rect 32128 9522 32180 9528
rect 31852 9444 31904 9450
rect 31852 9386 31904 9392
rect 31944 9444 31996 9450
rect 31944 9386 31996 9392
rect 31956 9178 31984 9386
rect 31944 9172 31996 9178
rect 31944 9114 31996 9120
rect 32140 9110 32168 9522
rect 32324 9382 32352 9930
rect 32416 9382 32444 10639
rect 32588 10610 32640 10616
rect 32772 10668 32824 10674
rect 32772 10610 32824 10616
rect 32494 10160 32550 10169
rect 32494 10095 32550 10104
rect 32312 9376 32364 9382
rect 32312 9318 32364 9324
rect 32404 9376 32456 9382
rect 32404 9318 32456 9324
rect 32220 9172 32272 9178
rect 32220 9114 32272 9120
rect 32128 9104 32180 9110
rect 31772 9030 31892 9058
rect 32128 9046 32180 9052
rect 31760 8968 31812 8974
rect 31760 8910 31812 8916
rect 31484 8628 31536 8634
rect 31484 8570 31536 8576
rect 31300 8492 31352 8498
rect 31300 8434 31352 8440
rect 29092 8084 29144 8090
rect 29092 8026 29144 8032
rect 31312 7954 31340 8434
rect 31772 8294 31800 8910
rect 31760 8288 31812 8294
rect 31760 8230 31812 8236
rect 31772 8022 31800 8230
rect 31760 8016 31812 8022
rect 31760 7958 31812 7964
rect 30840 7948 30892 7954
rect 30840 7890 30892 7896
rect 31300 7948 31352 7954
rect 31300 7890 31352 7896
rect 28724 7880 28776 7886
rect 28724 7822 28776 7828
rect 29552 7880 29604 7886
rect 29552 7822 29604 7828
rect 29564 7478 29592 7822
rect 29828 7812 29880 7818
rect 29828 7754 29880 7760
rect 30380 7812 30432 7818
rect 30380 7754 30432 7760
rect 29552 7472 29604 7478
rect 29552 7414 29604 7420
rect 29840 7274 29868 7754
rect 30392 7546 30420 7754
rect 30380 7540 30432 7546
rect 30432 7500 30512 7528
rect 30380 7482 30432 7488
rect 29828 7268 29880 7274
rect 29828 7210 29880 7216
rect 29276 7200 29328 7206
rect 29276 7142 29328 7148
rect 28632 6248 28684 6254
rect 28684 6208 28764 6236
rect 28632 6190 28684 6196
rect 28736 5574 28764 6208
rect 29184 6112 29236 6118
rect 29184 6054 29236 6060
rect 29196 5710 29224 6054
rect 29288 5914 29316 7142
rect 30380 6656 30432 6662
rect 30380 6598 30432 6604
rect 30392 6458 30420 6598
rect 30380 6452 30432 6458
rect 30380 6394 30432 6400
rect 29460 6316 29512 6322
rect 29460 6258 29512 6264
rect 29276 5908 29328 5914
rect 29276 5850 29328 5856
rect 29184 5704 29236 5710
rect 29184 5646 29236 5652
rect 28724 5568 28776 5574
rect 28724 5510 28776 5516
rect 28172 5364 28224 5370
rect 28172 5306 28224 5312
rect 28080 5296 28132 5302
rect 28080 5238 28132 5244
rect 28080 5024 28132 5030
rect 28080 4966 28132 4972
rect 28092 4554 28120 4966
rect 28080 4548 28132 4554
rect 28080 4490 28132 4496
rect 27988 3936 28040 3942
rect 28092 3890 28120 4490
rect 28736 4078 28764 5510
rect 29472 5370 29500 6258
rect 30484 5642 30512 7500
rect 30852 7290 30880 7890
rect 31300 7744 31352 7750
rect 31300 7686 31352 7692
rect 31312 7410 31340 7686
rect 31300 7404 31352 7410
rect 31300 7346 31352 7352
rect 30668 7274 30880 7290
rect 30656 7268 30880 7274
rect 30708 7262 30880 7268
rect 30656 7210 30708 7216
rect 30668 6866 30696 7210
rect 30656 6860 30708 6866
rect 30656 6802 30708 6808
rect 30380 5636 30432 5642
rect 30380 5578 30432 5584
rect 30472 5636 30524 5642
rect 30472 5578 30524 5584
rect 30392 5370 30420 5578
rect 29460 5364 29512 5370
rect 29460 5306 29512 5312
rect 30380 5364 30432 5370
rect 30380 5306 30432 5312
rect 28724 4072 28776 4078
rect 28724 4014 28776 4020
rect 28040 3884 28120 3890
rect 27988 3878 28120 3884
rect 28000 3862 28120 3878
rect 27896 3732 27948 3738
rect 27896 3674 27948 3680
rect 28092 3602 28120 3862
rect 28080 3596 28132 3602
rect 28080 3538 28132 3544
rect 30380 3596 30432 3602
rect 30380 3538 30432 3544
rect 27804 3460 27856 3466
rect 27804 3402 27856 3408
rect 28092 3194 28120 3538
rect 29368 3528 29420 3534
rect 29368 3470 29420 3476
rect 30288 3528 30340 3534
rect 30288 3470 30340 3476
rect 28816 3460 28868 3466
rect 28816 3402 28868 3408
rect 28356 3392 28408 3398
rect 28356 3334 28408 3340
rect 28080 3188 28132 3194
rect 28080 3130 28132 3136
rect 28368 3126 28396 3334
rect 28828 3126 28856 3402
rect 26056 3120 26108 3126
rect 26056 3062 26108 3068
rect 28356 3120 28408 3126
rect 28356 3062 28408 3068
rect 28816 3120 28868 3126
rect 28816 3062 28868 3068
rect 23940 3052 23992 3058
rect 23940 2994 23992 3000
rect 29000 2984 29052 2990
rect 29000 2926 29052 2932
rect 23388 2916 23440 2922
rect 23388 2858 23440 2864
rect 23296 2508 23348 2514
rect 23296 2450 23348 2456
rect 23400 2446 23428 2858
rect 29012 2650 29040 2926
rect 29380 2650 29408 3470
rect 30300 2650 30328 3470
rect 30392 3126 30420 3538
rect 30564 3460 30616 3466
rect 30564 3402 30616 3408
rect 30380 3120 30432 3126
rect 30380 3062 30432 3068
rect 30576 2774 30604 3402
rect 30668 2854 30696 6802
rect 31312 6798 31340 7346
rect 31668 7200 31720 7206
rect 31668 7142 31720 7148
rect 31300 6792 31352 6798
rect 31300 6734 31352 6740
rect 31392 6248 31444 6254
rect 31392 6190 31444 6196
rect 31404 5166 31432 6190
rect 31680 5302 31708 7142
rect 31772 6254 31800 7958
rect 31864 7546 31892 9030
rect 32140 8090 32168 9046
rect 32232 8430 32260 9114
rect 32508 9058 32536 10095
rect 32600 10062 32628 10610
rect 32680 10124 32732 10130
rect 32680 10066 32732 10072
rect 32588 10056 32640 10062
rect 32588 9998 32640 10004
rect 32600 9722 32628 9998
rect 32588 9716 32640 9722
rect 32588 9658 32640 9664
rect 32692 9602 32720 10066
rect 32784 9926 32812 10610
rect 32968 10266 32996 12192
rect 33048 12174 33100 12180
rect 33046 11928 33102 11937
rect 33244 11898 33272 12582
rect 33336 12238 33364 13262
rect 33520 12986 33548 13806
rect 33508 12980 33560 12986
rect 33508 12922 33560 12928
rect 33416 12912 33468 12918
rect 33416 12854 33468 12860
rect 33324 12232 33376 12238
rect 33324 12174 33376 12180
rect 33322 11928 33378 11937
rect 33046 11863 33102 11872
rect 33232 11892 33284 11898
rect 33060 11762 33088 11863
rect 33322 11863 33324 11872
rect 33232 11834 33284 11840
rect 33376 11863 33378 11872
rect 33324 11834 33376 11840
rect 33048 11756 33100 11762
rect 33048 11698 33100 11704
rect 33324 11756 33376 11762
rect 33324 11698 33376 11704
rect 33336 11354 33364 11698
rect 33428 11558 33456 12854
rect 33508 12844 33560 12850
rect 33508 12786 33560 12792
rect 33416 11552 33468 11558
rect 33416 11494 33468 11500
rect 33324 11348 33376 11354
rect 33324 11290 33376 11296
rect 33336 11150 33364 11290
rect 33520 11218 33548 12786
rect 33704 12714 33732 13806
rect 33968 13252 34020 13258
rect 33968 13194 34020 13200
rect 33692 12708 33744 12714
rect 33692 12650 33744 12656
rect 33784 12436 33836 12442
rect 33784 12378 33836 12384
rect 33690 12336 33746 12345
rect 33690 12271 33746 12280
rect 33704 12238 33732 12271
rect 33796 12238 33824 12378
rect 33980 12238 34008 13194
rect 34242 12336 34298 12345
rect 34242 12271 34244 12280
rect 34296 12271 34298 12280
rect 34244 12242 34296 12248
rect 33692 12232 33744 12238
rect 33784 12232 33836 12238
rect 33692 12174 33744 12180
rect 33782 12200 33784 12209
rect 33968 12232 34020 12238
rect 33836 12200 33838 12209
rect 33600 11756 33652 11762
rect 33600 11698 33652 11704
rect 33508 11212 33560 11218
rect 33508 11154 33560 11160
rect 33324 11144 33376 11150
rect 33324 11086 33376 11092
rect 33048 10668 33100 10674
rect 33048 10610 33100 10616
rect 32956 10260 33008 10266
rect 32956 10202 33008 10208
rect 32772 9920 32824 9926
rect 32824 9868 32996 9874
rect 32772 9862 32996 9868
rect 32784 9846 32996 9862
rect 32968 9722 32996 9846
rect 33060 9738 33088 10610
rect 33612 10169 33640 11698
rect 33598 10160 33654 10169
rect 33598 10095 33654 10104
rect 33704 9994 33732 12174
rect 33968 12174 34020 12180
rect 34428 12232 34480 12238
rect 34428 12174 34480 12180
rect 33782 12135 33838 12144
rect 33784 11756 33836 11762
rect 33784 11698 33836 11704
rect 33796 10062 33824 11698
rect 34336 11552 34388 11558
rect 34336 11494 34388 11500
rect 34348 11082 34376 11494
rect 34440 11098 34468 12174
rect 34612 11756 34664 11762
rect 34612 11698 34664 11704
rect 34624 11665 34652 11698
rect 34610 11656 34666 11665
rect 34610 11591 34666 11600
rect 34336 11076 34388 11082
rect 34440 11070 34560 11098
rect 34336 11018 34388 11024
rect 34532 11014 34560 11070
rect 34428 11008 34480 11014
rect 34428 10950 34480 10956
rect 34520 11008 34572 11014
rect 34520 10950 34572 10956
rect 34440 10674 34468 10950
rect 34428 10668 34480 10674
rect 34428 10610 34480 10616
rect 34624 10470 34652 11591
rect 34716 10690 34744 14418
rect 35268 14278 35296 14418
rect 35360 14346 35388 16118
rect 35452 16046 35480 16487
rect 35992 16458 36044 16464
rect 35594 16348 35902 16357
rect 35594 16346 35600 16348
rect 35656 16346 35680 16348
rect 35736 16346 35760 16348
rect 35816 16346 35840 16348
rect 35896 16346 35902 16348
rect 35656 16294 35658 16346
rect 35838 16294 35840 16346
rect 35594 16292 35600 16294
rect 35656 16292 35680 16294
rect 35736 16292 35760 16294
rect 35816 16292 35840 16294
rect 35896 16292 35902 16294
rect 35594 16283 35902 16292
rect 35808 16244 35860 16250
rect 35808 16186 35860 16192
rect 35440 16040 35492 16046
rect 35440 15982 35492 15988
rect 35820 15910 35848 16186
rect 36004 15978 36032 16458
rect 36084 16448 36136 16454
rect 36084 16390 36136 16396
rect 36096 16114 36124 16390
rect 36188 16250 36216 17002
rect 36176 16244 36228 16250
rect 36176 16186 36228 16192
rect 36084 16108 36136 16114
rect 36084 16050 36136 16056
rect 35992 15972 36044 15978
rect 35992 15914 36044 15920
rect 35716 15904 35768 15910
rect 35716 15846 35768 15852
rect 35808 15904 35860 15910
rect 35808 15846 35860 15852
rect 35728 15570 35756 15846
rect 35716 15564 35768 15570
rect 35716 15506 35768 15512
rect 35594 15260 35902 15269
rect 35594 15258 35600 15260
rect 35656 15258 35680 15260
rect 35736 15258 35760 15260
rect 35816 15258 35840 15260
rect 35896 15258 35902 15260
rect 35656 15206 35658 15258
rect 35838 15206 35840 15258
rect 35594 15204 35600 15206
rect 35656 15204 35680 15206
rect 35736 15204 35760 15206
rect 35816 15204 35840 15206
rect 35896 15204 35902 15206
rect 35594 15195 35902 15204
rect 35440 15020 35492 15026
rect 35440 14962 35492 14968
rect 35348 14340 35400 14346
rect 35348 14282 35400 14288
rect 35256 14272 35308 14278
rect 35256 14214 35308 14220
rect 35268 13938 35296 14214
rect 35256 13932 35308 13938
rect 35256 13874 35308 13880
rect 34934 13628 35242 13637
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13563 35242 13572
rect 35452 13530 35480 14962
rect 36280 14618 36308 19450
rect 36360 19372 36412 19378
rect 36360 19314 36412 19320
rect 35992 14612 36044 14618
rect 35992 14554 36044 14560
rect 36268 14612 36320 14618
rect 36268 14554 36320 14560
rect 35594 14172 35902 14181
rect 35594 14170 35600 14172
rect 35656 14170 35680 14172
rect 35736 14170 35760 14172
rect 35816 14170 35840 14172
rect 35896 14170 35902 14172
rect 35656 14118 35658 14170
rect 35838 14118 35840 14170
rect 35594 14116 35600 14118
rect 35656 14116 35680 14118
rect 35736 14116 35760 14118
rect 35816 14116 35840 14118
rect 35896 14116 35902 14118
rect 35594 14107 35902 14116
rect 36004 14006 36032 14554
rect 36176 14408 36228 14414
rect 36176 14350 36228 14356
rect 36188 14074 36216 14350
rect 36176 14068 36228 14074
rect 36176 14010 36228 14016
rect 35992 14000 36044 14006
rect 35992 13942 36044 13948
rect 36268 13932 36320 13938
rect 36268 13874 36320 13880
rect 36084 13796 36136 13802
rect 36084 13738 36136 13744
rect 35440 13524 35492 13530
rect 35440 13466 35492 13472
rect 36096 13326 36124 13738
rect 36280 13530 36308 13874
rect 36372 13870 36400 19314
rect 36464 17542 36492 19722
rect 36728 19712 36780 19718
rect 36728 19654 36780 19660
rect 36544 17672 36596 17678
rect 36544 17614 36596 17620
rect 36452 17536 36504 17542
rect 36452 17478 36504 17484
rect 36556 17202 36584 17614
rect 36544 17196 36596 17202
rect 36544 17138 36596 17144
rect 36544 17060 36596 17066
rect 36544 17002 36596 17008
rect 36556 16522 36584 17002
rect 36636 16992 36688 16998
rect 36636 16934 36688 16940
rect 36648 16590 36676 16934
rect 36740 16726 36768 19654
rect 36820 18624 36872 18630
rect 36818 18592 36820 18601
rect 36872 18592 36874 18601
rect 36818 18527 36874 18536
rect 36820 17672 36872 17678
rect 36820 17614 36872 17620
rect 36832 17338 36860 17614
rect 36820 17332 36872 17338
rect 36820 17274 36872 17280
rect 36728 16720 36780 16726
rect 36820 16720 36872 16726
rect 36728 16662 36780 16668
rect 36818 16688 36820 16697
rect 36872 16688 36874 16697
rect 36818 16623 36874 16632
rect 36636 16584 36688 16590
rect 36636 16526 36688 16532
rect 36544 16516 36596 16522
rect 36544 16458 36596 16464
rect 36544 16108 36596 16114
rect 36544 16050 36596 16056
rect 36556 15706 36584 16050
rect 36544 15700 36596 15706
rect 36544 15642 36596 15648
rect 36452 14816 36504 14822
rect 36452 14758 36504 14764
rect 36464 14414 36492 14758
rect 36452 14408 36504 14414
rect 36452 14350 36504 14356
rect 36544 13932 36596 13938
rect 36544 13874 36596 13880
rect 36360 13864 36412 13870
rect 36360 13806 36412 13812
rect 36556 13802 36584 13874
rect 36648 13841 36676 16526
rect 36728 16448 36780 16454
rect 36728 16390 36780 16396
rect 36740 15434 36768 16390
rect 36832 16114 36860 16623
rect 36820 16108 36872 16114
rect 36820 16050 36872 16056
rect 36820 15904 36872 15910
rect 36820 15846 36872 15852
rect 36728 15428 36780 15434
rect 36728 15370 36780 15376
rect 36634 13832 36690 13841
rect 36544 13796 36596 13802
rect 36634 13767 36690 13776
rect 36544 13738 36596 13744
rect 36452 13728 36504 13734
rect 36452 13670 36504 13676
rect 36464 13530 36492 13670
rect 36268 13524 36320 13530
rect 36268 13466 36320 13472
rect 36452 13524 36504 13530
rect 36452 13466 36504 13472
rect 36544 13524 36596 13530
rect 36544 13466 36596 13472
rect 36556 13410 36584 13466
rect 36464 13382 36584 13410
rect 36636 13388 36688 13394
rect 36464 13326 36492 13382
rect 36636 13330 36688 13336
rect 36084 13320 36136 13326
rect 36084 13262 36136 13268
rect 36452 13320 36504 13326
rect 36452 13262 36504 13268
rect 36544 13320 36596 13326
rect 36544 13262 36596 13268
rect 36556 13190 36584 13262
rect 36544 13184 36596 13190
rect 36544 13126 36596 13132
rect 35594 13084 35902 13093
rect 35594 13082 35600 13084
rect 35656 13082 35680 13084
rect 35736 13082 35760 13084
rect 35816 13082 35840 13084
rect 35896 13082 35902 13084
rect 35656 13030 35658 13082
rect 35838 13030 35840 13082
rect 35594 13028 35600 13030
rect 35656 13028 35680 13030
rect 35736 13028 35760 13030
rect 35816 13028 35840 13030
rect 35896 13028 35902 13030
rect 35594 13019 35902 13028
rect 36648 12986 36676 13330
rect 36636 12980 36688 12986
rect 36636 12922 36688 12928
rect 36268 12844 36320 12850
rect 36268 12786 36320 12792
rect 34934 12540 35242 12549
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12475 35242 12484
rect 35716 12436 35768 12442
rect 35716 12378 35768 12384
rect 35728 12238 35756 12378
rect 34888 12232 34940 12238
rect 34888 12174 34940 12180
rect 35164 12232 35216 12238
rect 35440 12232 35492 12238
rect 35164 12174 35216 12180
rect 35346 12200 35402 12209
rect 34900 11898 34928 12174
rect 35176 11914 35204 12174
rect 35440 12174 35492 12180
rect 35716 12232 35768 12238
rect 35716 12174 35768 12180
rect 35992 12232 36044 12238
rect 36044 12192 36124 12220
rect 35992 12174 36044 12180
rect 35346 12135 35402 12144
rect 35360 12102 35388 12135
rect 35348 12096 35400 12102
rect 35348 12038 35400 12044
rect 35176 11898 35296 11914
rect 34888 11892 34940 11898
rect 34888 11834 34940 11840
rect 35072 11892 35124 11898
rect 35176 11892 35308 11898
rect 35176 11886 35256 11892
rect 35072 11834 35124 11840
rect 35256 11834 35308 11840
rect 35084 11665 35112 11834
rect 35256 11756 35308 11762
rect 35256 11698 35308 11704
rect 35070 11656 35126 11665
rect 35070 11591 35126 11600
rect 35268 11540 35296 11698
rect 35348 11688 35400 11694
rect 35348 11630 35400 11636
rect 35360 11558 35388 11630
rect 34808 11512 35296 11540
rect 35348 11552 35400 11558
rect 34808 11234 34836 11512
rect 35348 11494 35400 11500
rect 34934 11452 35242 11461
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11387 35242 11396
rect 35452 11286 35480 12174
rect 35992 12096 36044 12102
rect 35992 12038 36044 12044
rect 35594 11996 35902 12005
rect 35594 11994 35600 11996
rect 35656 11994 35680 11996
rect 35736 11994 35760 11996
rect 35816 11994 35840 11996
rect 35896 11994 35902 11996
rect 35656 11942 35658 11994
rect 35838 11942 35840 11994
rect 35594 11940 35600 11942
rect 35656 11940 35680 11942
rect 35736 11940 35760 11942
rect 35816 11940 35840 11942
rect 35896 11940 35902 11942
rect 35594 11931 35902 11940
rect 36004 11830 36032 12038
rect 36096 11830 36124 12192
rect 36280 12170 36308 12786
rect 36268 12164 36320 12170
rect 36188 12124 36268 12152
rect 35992 11824 36044 11830
rect 35992 11766 36044 11772
rect 36084 11824 36136 11830
rect 36084 11766 36136 11772
rect 36188 11608 36216 12124
rect 36268 12106 36320 12112
rect 36452 12096 36504 12102
rect 36452 12038 36504 12044
rect 36268 11756 36320 11762
rect 36320 11716 36400 11744
rect 36268 11698 36320 11704
rect 36268 11620 36320 11626
rect 36188 11580 36268 11608
rect 35440 11280 35492 11286
rect 35070 11248 35126 11257
rect 34808 11206 34928 11234
rect 34900 11150 34928 11206
rect 35440 11222 35492 11228
rect 35070 11183 35126 11192
rect 34796 11144 34848 11150
rect 34796 11086 34848 11092
rect 34888 11144 34940 11150
rect 34888 11086 34940 11092
rect 34808 10810 34836 11086
rect 34796 10804 34848 10810
rect 34796 10746 34848 10752
rect 34900 10742 34928 11086
rect 35084 10742 35112 11183
rect 35440 11144 35492 11150
rect 35346 11112 35402 11121
rect 35440 11086 35492 11092
rect 35346 11047 35348 11056
rect 35400 11047 35402 11056
rect 35348 11018 35400 11024
rect 35452 10792 35480 11086
rect 35594 10908 35902 10917
rect 35594 10906 35600 10908
rect 35656 10906 35680 10908
rect 35736 10906 35760 10908
rect 35816 10906 35840 10908
rect 35896 10906 35902 10908
rect 35656 10854 35658 10906
rect 35838 10854 35840 10906
rect 35594 10852 35600 10854
rect 35656 10852 35680 10854
rect 35736 10852 35760 10854
rect 35816 10852 35840 10854
rect 35896 10852 35902 10854
rect 35594 10843 35902 10852
rect 36188 10810 36216 11580
rect 36268 11562 36320 11568
rect 36176 10804 36228 10810
rect 35452 10764 35756 10792
rect 34888 10736 34940 10742
rect 34716 10662 34836 10690
rect 35072 10736 35124 10742
rect 34888 10678 34940 10684
rect 35070 10704 35072 10713
rect 35124 10704 35126 10713
rect 34704 10532 34756 10538
rect 34704 10474 34756 10480
rect 34612 10464 34664 10470
rect 34612 10406 34664 10412
rect 33784 10056 33836 10062
rect 33784 9998 33836 10004
rect 33692 9988 33744 9994
rect 33692 9930 33744 9936
rect 32956 9716 33008 9722
rect 32956 9658 33008 9664
rect 33060 9710 33456 9738
rect 32600 9586 32720 9602
rect 32968 9586 32996 9658
rect 32588 9580 32720 9586
rect 32640 9574 32720 9580
rect 32956 9580 33008 9586
rect 32588 9522 32640 9528
rect 32956 9522 33008 9528
rect 32600 9450 32628 9522
rect 32588 9444 32640 9450
rect 32588 9386 32640 9392
rect 32508 9030 32628 9058
rect 32312 8968 32364 8974
rect 32312 8910 32364 8916
rect 32496 8968 32548 8974
rect 32496 8910 32548 8916
rect 32324 8566 32352 8910
rect 32312 8560 32364 8566
rect 32312 8502 32364 8508
rect 32508 8498 32536 8910
rect 32600 8634 32628 9030
rect 32968 8838 32996 9522
rect 33060 9110 33088 9710
rect 33232 9580 33284 9586
rect 33232 9522 33284 9528
rect 33244 9178 33272 9522
rect 33428 9518 33456 9710
rect 33796 9586 33824 9998
rect 33784 9580 33836 9586
rect 33784 9522 33836 9528
rect 33416 9512 33468 9518
rect 33416 9454 33468 9460
rect 33416 9376 33468 9382
rect 33796 9330 33824 9522
rect 34716 9450 34744 10474
rect 34808 10198 34836 10662
rect 35070 10639 35126 10648
rect 35348 10668 35400 10674
rect 35348 10610 35400 10616
rect 35624 10668 35676 10674
rect 35624 10610 35676 10616
rect 34934 10364 35242 10373
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10299 35242 10308
rect 35360 10266 35388 10610
rect 35636 10538 35664 10610
rect 35624 10532 35676 10538
rect 35624 10474 35676 10480
rect 35728 10452 35756 10764
rect 36176 10746 36228 10752
rect 36084 10736 36136 10742
rect 36084 10678 36136 10684
rect 35900 10668 35952 10674
rect 35900 10610 35952 10616
rect 35912 10577 35940 10610
rect 35898 10568 35954 10577
rect 35898 10503 35954 10512
rect 36096 10470 36124 10678
rect 35808 10464 35860 10470
rect 35728 10424 35808 10452
rect 35808 10406 35860 10412
rect 35900 10464 35952 10470
rect 35900 10406 35952 10412
rect 36084 10464 36136 10470
rect 36084 10406 36136 10412
rect 35348 10260 35400 10266
rect 35348 10202 35400 10208
rect 35808 10260 35860 10266
rect 35808 10202 35860 10208
rect 34796 10192 34848 10198
rect 34796 10134 34848 10140
rect 35820 9926 35848 10202
rect 35912 10130 35940 10406
rect 36188 10198 36216 10746
rect 36372 10577 36400 11716
rect 36464 11354 36492 12038
rect 36544 11756 36596 11762
rect 36544 11698 36596 11704
rect 36636 11756 36688 11762
rect 36636 11698 36688 11704
rect 36452 11348 36504 11354
rect 36452 11290 36504 11296
rect 36464 10674 36492 11290
rect 36556 11218 36584 11698
rect 36648 11558 36676 11698
rect 36636 11552 36688 11558
rect 36636 11494 36688 11500
rect 36544 11212 36596 11218
rect 36544 11154 36596 11160
rect 36452 10668 36504 10674
rect 36452 10610 36504 10616
rect 36636 10668 36688 10674
rect 36636 10610 36688 10616
rect 36358 10568 36414 10577
rect 36358 10503 36414 10512
rect 36176 10192 36228 10198
rect 36176 10134 36228 10140
rect 36268 10192 36320 10198
rect 36268 10134 36320 10140
rect 35900 10124 35952 10130
rect 35900 10066 35952 10072
rect 36176 9988 36228 9994
rect 36280 9976 36308 10134
rect 36372 10062 36400 10503
rect 36360 10056 36412 10062
rect 36360 9998 36412 10004
rect 36228 9948 36308 9976
rect 36452 9988 36504 9994
rect 36176 9930 36228 9936
rect 36452 9930 36504 9936
rect 35808 9920 35860 9926
rect 35808 9862 35860 9868
rect 36084 9920 36136 9926
rect 36084 9862 36136 9868
rect 35594 9820 35902 9829
rect 35594 9818 35600 9820
rect 35656 9818 35680 9820
rect 35736 9818 35760 9820
rect 35816 9818 35840 9820
rect 35896 9818 35902 9820
rect 35656 9766 35658 9818
rect 35838 9766 35840 9818
rect 35594 9764 35600 9766
rect 35656 9764 35680 9766
rect 35736 9764 35760 9766
rect 35816 9764 35840 9766
rect 35896 9764 35902 9766
rect 35594 9755 35902 9764
rect 34704 9444 34756 9450
rect 34704 9386 34756 9392
rect 33468 9324 33824 9330
rect 33416 9318 33824 9324
rect 33428 9302 33824 9318
rect 34934 9276 35242 9285
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9211 35242 9220
rect 33232 9172 33284 9178
rect 33232 9114 33284 9120
rect 33048 9104 33100 9110
rect 33048 9046 33100 9052
rect 32956 8832 33008 8838
rect 32956 8774 33008 8780
rect 35992 8832 36044 8838
rect 35992 8774 36044 8780
rect 35594 8732 35902 8741
rect 35594 8730 35600 8732
rect 35656 8730 35680 8732
rect 35736 8730 35760 8732
rect 35816 8730 35840 8732
rect 35896 8730 35902 8732
rect 35656 8678 35658 8730
rect 35838 8678 35840 8730
rect 35594 8676 35600 8678
rect 35656 8676 35680 8678
rect 35736 8676 35760 8678
rect 35816 8676 35840 8678
rect 35896 8676 35902 8678
rect 35594 8667 35902 8676
rect 32588 8628 32640 8634
rect 32588 8570 32640 8576
rect 36004 8498 36032 8774
rect 36096 8566 36124 9862
rect 36464 8922 36492 9930
rect 36648 9586 36676 10610
rect 36636 9580 36688 9586
rect 36636 9522 36688 9528
rect 36648 9178 36676 9522
rect 36740 9178 36768 15370
rect 36832 14550 36860 15846
rect 36924 14618 36952 19790
rect 37096 18760 37148 18766
rect 37094 18728 37096 18737
rect 37148 18728 37150 18737
rect 37094 18663 37150 18672
rect 37096 18624 37148 18630
rect 37096 18566 37148 18572
rect 37108 18426 37136 18566
rect 37096 18420 37148 18426
rect 37096 18362 37148 18368
rect 37108 17814 37136 18362
rect 37096 17808 37148 17814
rect 37096 17750 37148 17756
rect 37094 17640 37150 17649
rect 37004 17604 37056 17610
rect 37094 17575 37096 17584
rect 37004 17546 37056 17552
rect 37148 17575 37150 17584
rect 37096 17546 37148 17552
rect 37016 17490 37044 17546
rect 37016 17462 37136 17490
rect 37108 16794 37136 17462
rect 37200 17338 37228 20198
rect 37372 19780 37424 19786
rect 37372 19722 37424 19728
rect 37384 19310 37412 19722
rect 37372 19304 37424 19310
rect 37372 19246 37424 19252
rect 37372 18352 37424 18358
rect 37372 18294 37424 18300
rect 37384 18086 37412 18294
rect 37372 18080 37424 18086
rect 37372 18022 37424 18028
rect 37188 17332 37240 17338
rect 37188 17274 37240 17280
rect 37200 16794 37228 17274
rect 37280 17128 37332 17134
rect 37280 17070 37332 17076
rect 37096 16788 37148 16794
rect 37096 16730 37148 16736
rect 37188 16788 37240 16794
rect 37188 16730 37240 16736
rect 37002 16552 37058 16561
rect 37292 16522 37320 17070
rect 37002 16487 37058 16496
rect 37280 16516 37332 16522
rect 37016 16114 37044 16487
rect 37280 16458 37332 16464
rect 37292 16425 37320 16458
rect 37278 16416 37334 16425
rect 37278 16351 37334 16360
rect 37004 16108 37056 16114
rect 37004 16050 37056 16056
rect 37004 15972 37056 15978
rect 37004 15914 37056 15920
rect 36912 14612 36964 14618
rect 36912 14554 36964 14560
rect 36820 14544 36872 14550
rect 36820 14486 36872 14492
rect 36832 14414 36860 14486
rect 36820 14408 36872 14414
rect 36820 14350 36872 14356
rect 36912 14340 36964 14346
rect 36912 14282 36964 14288
rect 36820 13728 36872 13734
rect 36820 13670 36872 13676
rect 36832 12850 36860 13670
rect 36924 13258 36952 14282
rect 37016 13938 37044 15914
rect 37280 15496 37332 15502
rect 37280 15438 37332 15444
rect 37292 14482 37320 15438
rect 37384 15366 37412 18022
rect 37568 17610 37596 22578
rect 37648 22432 37700 22438
rect 37648 22374 37700 22380
rect 37660 22030 37688 22374
rect 37648 22024 37700 22030
rect 37648 21966 37700 21972
rect 37752 18426 37780 24375
rect 37844 22778 37872 27066
rect 38476 25152 38528 25158
rect 38476 25094 38528 25100
rect 38016 24880 38068 24886
rect 38016 24822 38068 24828
rect 38028 23866 38056 24822
rect 38488 24818 38516 25094
rect 38476 24812 38528 24818
rect 38476 24754 38528 24760
rect 38292 24608 38344 24614
rect 38292 24550 38344 24556
rect 38304 24342 38332 24550
rect 38292 24336 38344 24342
rect 38292 24278 38344 24284
rect 37924 23860 37976 23866
rect 37924 23802 37976 23808
rect 38016 23860 38068 23866
rect 38016 23802 38068 23808
rect 37936 23594 37964 23802
rect 38304 23730 38332 24278
rect 38580 24041 38608 30058
rect 38672 29306 38700 30620
rect 38752 30660 38804 30666
rect 38752 30602 38804 30608
rect 38764 30190 38792 30602
rect 38844 30592 38896 30598
rect 38844 30534 38896 30540
rect 38856 30326 38884 30534
rect 38844 30320 38896 30326
rect 38844 30262 38896 30268
rect 43352 30320 43404 30326
rect 43352 30262 43404 30268
rect 42432 30252 42484 30258
rect 42432 30194 42484 30200
rect 42524 30252 42576 30258
rect 42524 30194 42576 30200
rect 42708 30252 42760 30258
rect 42708 30194 42760 30200
rect 38752 30184 38804 30190
rect 38752 30126 38804 30132
rect 40316 29776 40368 29782
rect 40316 29718 40368 29724
rect 40776 29776 40828 29782
rect 40776 29718 40828 29724
rect 39672 29640 39724 29646
rect 39672 29582 39724 29588
rect 38660 29300 38712 29306
rect 38660 29242 38712 29248
rect 39684 28966 39712 29582
rect 40328 29170 40356 29718
rect 40592 29640 40644 29646
rect 40592 29582 40644 29588
rect 40500 29504 40552 29510
rect 40500 29446 40552 29452
rect 39948 29164 40000 29170
rect 40224 29164 40276 29170
rect 40000 29124 40080 29152
rect 39948 29106 40000 29112
rect 39672 28960 39724 28966
rect 39672 28902 39724 28908
rect 39684 28558 39712 28902
rect 39672 28552 39724 28558
rect 39672 28494 39724 28500
rect 38936 28484 38988 28490
rect 38936 28426 38988 28432
rect 38948 28257 38976 28426
rect 38934 28248 38990 28257
rect 38934 28183 38990 28192
rect 40052 28150 40080 29124
rect 40224 29106 40276 29112
rect 40316 29164 40368 29170
rect 40316 29106 40368 29112
rect 40236 28558 40264 29106
rect 40224 28552 40276 28558
rect 40224 28494 40276 28500
rect 40040 28144 40092 28150
rect 40038 28112 40040 28121
rect 40092 28112 40094 28121
rect 38936 28076 38988 28082
rect 40038 28047 40094 28056
rect 38936 28018 38988 28024
rect 38948 26586 38976 28018
rect 39948 27328 40000 27334
rect 39948 27270 40000 27276
rect 39960 27130 39988 27270
rect 39948 27124 40000 27130
rect 39948 27066 40000 27072
rect 38936 26580 38988 26586
rect 38936 26522 38988 26528
rect 38660 26444 38712 26450
rect 38660 26386 38712 26392
rect 38672 25294 38700 26386
rect 38948 25974 38976 26522
rect 39028 26512 39080 26518
rect 39028 26454 39080 26460
rect 38936 25968 38988 25974
rect 38936 25910 38988 25916
rect 38752 25696 38804 25702
rect 38752 25638 38804 25644
rect 38764 25294 38792 25638
rect 38936 25492 38988 25498
rect 38936 25434 38988 25440
rect 38844 25424 38896 25430
rect 38844 25366 38896 25372
rect 38660 25288 38712 25294
rect 38660 25230 38712 25236
rect 38752 25288 38804 25294
rect 38752 25230 38804 25236
rect 38566 24032 38622 24041
rect 38566 23967 38622 23976
rect 38384 23860 38436 23866
rect 38384 23802 38436 23808
rect 38108 23724 38160 23730
rect 38292 23724 38344 23730
rect 38160 23684 38292 23712
rect 38108 23666 38160 23672
rect 38292 23666 38344 23672
rect 38120 23633 38148 23666
rect 38106 23624 38162 23633
rect 37924 23588 37976 23594
rect 38106 23559 38162 23568
rect 37924 23530 37976 23536
rect 38304 23186 38332 23666
rect 38292 23180 38344 23186
rect 38292 23122 38344 23128
rect 37832 22772 37884 22778
rect 37832 22714 37884 22720
rect 38396 22642 38424 23802
rect 38672 23798 38700 25230
rect 38856 25226 38884 25366
rect 38844 25220 38896 25226
rect 38844 25162 38896 25168
rect 38856 25129 38884 25162
rect 38842 25120 38898 25129
rect 38842 25055 38898 25064
rect 38856 24857 38884 25055
rect 38842 24848 38898 24857
rect 38842 24783 38898 24792
rect 38752 24676 38804 24682
rect 38752 24618 38804 24624
rect 38764 24585 38792 24618
rect 38750 24576 38806 24585
rect 38750 24511 38806 24520
rect 38764 24070 38792 24511
rect 38752 24064 38804 24070
rect 38752 24006 38804 24012
rect 38660 23792 38712 23798
rect 38660 23734 38712 23740
rect 38568 23520 38620 23526
rect 38764 23474 38792 24006
rect 38948 23526 38976 25434
rect 39040 25294 39068 26454
rect 39960 26382 39988 27066
rect 40224 26988 40276 26994
rect 40224 26930 40276 26936
rect 40236 26586 40264 26930
rect 40224 26580 40276 26586
rect 40224 26522 40276 26528
rect 40132 26512 40184 26518
rect 40328 26466 40356 29106
rect 40408 29096 40460 29102
rect 40408 29038 40460 29044
rect 40420 28914 40448 29038
rect 40512 29034 40540 29446
rect 40500 29028 40552 29034
rect 40500 28970 40552 28976
rect 40420 28886 40540 28914
rect 40512 28558 40540 28886
rect 40604 28694 40632 29582
rect 40788 29170 40816 29718
rect 41064 29566 41276 29594
rect 41064 29238 41092 29566
rect 41248 29510 41276 29566
rect 41420 29572 41472 29578
rect 41420 29514 41472 29520
rect 41144 29504 41196 29510
rect 41144 29446 41196 29452
rect 41236 29504 41288 29510
rect 41236 29446 41288 29452
rect 41156 29306 41184 29446
rect 41144 29300 41196 29306
rect 41144 29242 41196 29248
rect 41052 29232 41104 29238
rect 41052 29174 41104 29180
rect 40776 29164 40828 29170
rect 40776 29106 40828 29112
rect 41156 29034 41184 29242
rect 41432 29170 41460 29514
rect 41420 29164 41472 29170
rect 41420 29106 41472 29112
rect 41328 29096 41380 29102
rect 41328 29038 41380 29044
rect 41144 29028 41196 29034
rect 41144 28970 41196 28976
rect 41340 28694 41368 29038
rect 40592 28688 40644 28694
rect 40592 28630 40644 28636
rect 41328 28688 41380 28694
rect 41328 28630 41380 28636
rect 40500 28552 40552 28558
rect 40500 28494 40552 28500
rect 40512 27946 40540 28494
rect 41236 28484 41288 28490
rect 41236 28426 41288 28432
rect 41248 28218 41276 28426
rect 41236 28212 41288 28218
rect 41236 28154 41288 28160
rect 40500 27940 40552 27946
rect 40500 27882 40552 27888
rect 40960 27872 41012 27878
rect 40960 27814 41012 27820
rect 40972 27606 41000 27814
rect 40960 27600 41012 27606
rect 40960 27542 41012 27548
rect 40500 27532 40552 27538
rect 40500 27474 40552 27480
rect 40408 27396 40460 27402
rect 40408 27338 40460 27344
rect 40420 26926 40448 27338
rect 40408 26920 40460 26926
rect 40408 26862 40460 26868
rect 40184 26460 40356 26466
rect 40132 26454 40356 26460
rect 40144 26438 40356 26454
rect 39948 26376 40000 26382
rect 39948 26318 40000 26324
rect 39304 26240 39356 26246
rect 39304 26182 39356 26188
rect 39488 26240 39540 26246
rect 39488 26182 39540 26188
rect 40040 26240 40092 26246
rect 40040 26182 40092 26188
rect 40224 26240 40276 26246
rect 40224 26182 40276 26188
rect 39316 25906 39344 26182
rect 39304 25900 39356 25906
rect 39304 25842 39356 25848
rect 39500 25838 39528 26182
rect 40052 26042 40080 26182
rect 40040 26036 40092 26042
rect 40040 25978 40092 25984
rect 39672 25900 39724 25906
rect 39672 25842 39724 25848
rect 39396 25832 39448 25838
rect 39396 25774 39448 25780
rect 39488 25832 39540 25838
rect 39488 25774 39540 25780
rect 39408 25702 39436 25774
rect 39396 25696 39448 25702
rect 39396 25638 39448 25644
rect 39118 25392 39174 25401
rect 39500 25362 39528 25774
rect 39118 25327 39174 25336
rect 39488 25356 39540 25362
rect 39132 25294 39160 25327
rect 39488 25298 39540 25304
rect 39028 25288 39080 25294
rect 39028 25230 39080 25236
rect 39120 25288 39172 25294
rect 39120 25230 39172 25236
rect 39396 25288 39448 25294
rect 39396 25230 39448 25236
rect 39304 25152 39356 25158
rect 39132 25112 39304 25140
rect 39132 24070 39160 25112
rect 39304 25094 39356 25100
rect 39120 24064 39172 24070
rect 39120 24006 39172 24012
rect 38620 23468 38792 23474
rect 38568 23462 38792 23468
rect 38936 23520 38988 23526
rect 38936 23462 38988 23468
rect 38580 23446 38792 23462
rect 38948 23254 38976 23462
rect 38936 23248 38988 23254
rect 38936 23190 38988 23196
rect 39132 23118 39160 24006
rect 39212 23724 39264 23730
rect 39212 23666 39264 23672
rect 39224 23322 39252 23666
rect 39212 23316 39264 23322
rect 39212 23258 39264 23264
rect 39408 23202 39436 25230
rect 39684 25226 39712 25842
rect 39948 25832 40000 25838
rect 39948 25774 40000 25780
rect 39856 25764 39908 25770
rect 39856 25706 39908 25712
rect 39868 25294 39896 25706
rect 39856 25288 39908 25294
rect 39856 25230 39908 25236
rect 39672 25220 39724 25226
rect 39672 25162 39724 25168
rect 39960 24818 39988 25774
rect 40052 25294 40080 25978
rect 40236 25498 40264 26182
rect 40328 25838 40356 26438
rect 40420 26364 40448 26862
rect 40512 26790 40540 27474
rect 40972 26976 41000 27542
rect 41248 27334 41276 28154
rect 41432 27470 41460 29106
rect 42444 28762 42472 30194
rect 42536 29850 42564 30194
rect 42720 29850 42748 30194
rect 42524 29844 42576 29850
rect 42524 29786 42576 29792
rect 42708 29844 42760 29850
rect 42708 29786 42760 29792
rect 42536 29646 42564 29786
rect 42524 29640 42576 29646
rect 42524 29582 42576 29588
rect 42432 28756 42484 28762
rect 42432 28698 42484 28704
rect 42248 28484 42300 28490
rect 42248 28426 42300 28432
rect 42260 28082 42288 28426
rect 42248 28076 42300 28082
rect 42248 28018 42300 28024
rect 41788 28008 41840 28014
rect 41788 27950 41840 27956
rect 41604 27532 41656 27538
rect 41604 27474 41656 27480
rect 41420 27464 41472 27470
rect 41420 27406 41472 27412
rect 41236 27328 41288 27334
rect 41236 27270 41288 27276
rect 41248 26994 41276 27270
rect 41052 26988 41104 26994
rect 40972 26948 41052 26976
rect 41052 26930 41104 26936
rect 41236 26988 41288 26994
rect 41236 26930 41288 26936
rect 41616 26926 41644 27474
rect 41800 27402 41828 27950
rect 41788 27396 41840 27402
rect 41788 27338 41840 27344
rect 41800 26994 41828 27338
rect 41788 26988 41840 26994
rect 41788 26930 41840 26936
rect 41604 26920 41656 26926
rect 41604 26862 41656 26868
rect 42340 26920 42392 26926
rect 42340 26862 42392 26868
rect 40500 26784 40552 26790
rect 40500 26726 40552 26732
rect 40512 26586 40540 26726
rect 40500 26580 40552 26586
rect 40500 26522 40552 26528
rect 42064 26444 42116 26450
rect 42064 26386 42116 26392
rect 40500 26376 40552 26382
rect 40420 26336 40500 26364
rect 40500 26318 40552 26324
rect 40868 25968 40920 25974
rect 40868 25910 40920 25916
rect 40316 25832 40368 25838
rect 40316 25774 40368 25780
rect 40224 25492 40276 25498
rect 40224 25434 40276 25440
rect 40328 25362 40356 25774
rect 40592 25696 40644 25702
rect 40592 25638 40644 25644
rect 40316 25356 40368 25362
rect 40316 25298 40368 25304
rect 40040 25288 40092 25294
rect 40040 25230 40092 25236
rect 40052 24886 40080 25230
rect 40040 24880 40092 24886
rect 40040 24822 40092 24828
rect 39948 24812 40000 24818
rect 39948 24754 40000 24760
rect 39856 24676 39908 24682
rect 39856 24618 39908 24624
rect 39580 24608 39632 24614
rect 39580 24550 39632 24556
rect 39672 24608 39724 24614
rect 39672 24550 39724 24556
rect 39592 24206 39620 24550
rect 39684 24274 39712 24550
rect 39764 24336 39816 24342
rect 39764 24278 39816 24284
rect 39672 24268 39724 24274
rect 39672 24210 39724 24216
rect 39580 24200 39632 24206
rect 39580 24142 39632 24148
rect 39488 24132 39540 24138
rect 39488 24074 39540 24080
rect 39316 23174 39436 23202
rect 39120 23112 39172 23118
rect 39120 23054 39172 23060
rect 38660 22976 38712 22982
rect 38660 22918 38712 22924
rect 38672 22778 38700 22918
rect 38660 22772 38712 22778
rect 38660 22714 38712 22720
rect 38384 22636 38436 22642
rect 38384 22578 38436 22584
rect 37832 22432 37884 22438
rect 37832 22374 37884 22380
rect 37844 20505 37872 22374
rect 38476 21888 38528 21894
rect 38476 21830 38528 21836
rect 37924 20936 37976 20942
rect 37924 20878 37976 20884
rect 37830 20496 37886 20505
rect 37830 20431 37886 20440
rect 37936 19922 37964 20878
rect 38200 20868 38252 20874
rect 38200 20810 38252 20816
rect 38212 20602 38240 20810
rect 38488 20806 38516 21830
rect 38672 21146 38700 22714
rect 39132 22642 39160 23054
rect 39120 22636 39172 22642
rect 39120 22578 39172 22584
rect 39316 22094 39344 23174
rect 39396 23112 39448 23118
rect 39396 23054 39448 23060
rect 39408 22778 39436 23054
rect 39396 22772 39448 22778
rect 39396 22714 39448 22720
rect 39500 22094 39528 24074
rect 39592 23322 39620 24142
rect 39776 23798 39804 24278
rect 39868 23882 39896 24618
rect 39960 24410 39988 24754
rect 39948 24404 40000 24410
rect 39948 24346 40000 24352
rect 39960 24206 39988 24346
rect 39948 24200 40000 24206
rect 39948 24142 40000 24148
rect 40052 24138 40080 24822
rect 40132 24608 40184 24614
rect 40132 24550 40184 24556
rect 40500 24608 40552 24614
rect 40500 24550 40552 24556
rect 40040 24132 40092 24138
rect 40040 24074 40092 24080
rect 39948 24064 40000 24070
rect 40000 24012 40080 24018
rect 39948 24006 40080 24012
rect 39960 23990 40080 24006
rect 39868 23866 39988 23882
rect 40052 23866 40080 23990
rect 39856 23860 39988 23866
rect 39908 23854 39988 23860
rect 39856 23802 39908 23808
rect 39672 23792 39724 23798
rect 39670 23760 39672 23769
rect 39764 23792 39816 23798
rect 39724 23760 39726 23769
rect 39764 23734 39816 23740
rect 39670 23695 39726 23704
rect 39580 23316 39632 23322
rect 39580 23258 39632 23264
rect 39580 22976 39632 22982
rect 39580 22918 39632 22924
rect 39592 22642 39620 22918
rect 39580 22636 39632 22642
rect 39580 22578 39632 22584
rect 39316 22066 39436 22094
rect 39500 22066 39620 22094
rect 39304 21616 39356 21622
rect 39304 21558 39356 21564
rect 38660 21140 38712 21146
rect 38660 21082 38712 21088
rect 38476 20800 38528 20806
rect 38476 20742 38528 20748
rect 38200 20596 38252 20602
rect 38200 20538 38252 20544
rect 37924 19916 37976 19922
rect 37924 19858 37976 19864
rect 37936 19258 37964 19858
rect 38488 19854 38516 20742
rect 38476 19848 38528 19854
rect 38476 19790 38528 19796
rect 38108 19372 38160 19378
rect 38108 19314 38160 19320
rect 38016 19304 38068 19310
rect 37936 19252 38016 19258
rect 37936 19246 38068 19252
rect 37936 19230 38056 19246
rect 37936 18834 37964 19230
rect 37924 18828 37976 18834
rect 37924 18770 37976 18776
rect 37740 18420 37792 18426
rect 37740 18362 37792 18368
rect 38016 18420 38068 18426
rect 38016 18362 38068 18368
rect 38028 18329 38056 18362
rect 38014 18320 38070 18329
rect 37740 18284 37792 18290
rect 38014 18255 38070 18264
rect 37740 18226 37792 18232
rect 37752 17746 37780 18226
rect 38028 17882 38056 18255
rect 38016 17876 38068 17882
rect 38016 17818 38068 17824
rect 38120 17814 38148 19314
rect 38200 18692 38252 18698
rect 38200 18634 38252 18640
rect 38292 18692 38344 18698
rect 38292 18634 38344 18640
rect 38212 18358 38240 18634
rect 38200 18352 38252 18358
rect 38200 18294 38252 18300
rect 38304 18086 38332 18634
rect 38672 18442 38700 21082
rect 39316 20942 39344 21558
rect 39304 20936 39356 20942
rect 39304 20878 39356 20884
rect 39028 20596 39080 20602
rect 39028 20538 39080 20544
rect 38844 19712 38896 19718
rect 38844 19654 38896 19660
rect 38936 19712 38988 19718
rect 38936 19654 38988 19660
rect 38488 18414 38700 18442
rect 38292 18080 38344 18086
rect 38292 18022 38344 18028
rect 38488 17882 38516 18414
rect 38568 18284 38620 18290
rect 38568 18226 38620 18232
rect 38660 18284 38712 18290
rect 38712 18244 38792 18272
rect 38660 18226 38712 18232
rect 38476 17876 38528 17882
rect 38476 17818 38528 17824
rect 38108 17808 38160 17814
rect 38108 17750 38160 17756
rect 37740 17740 37792 17746
rect 37740 17682 37792 17688
rect 37556 17604 37608 17610
rect 37556 17546 37608 17552
rect 38120 17338 38148 17750
rect 38108 17332 38160 17338
rect 38108 17274 38160 17280
rect 38120 16946 38148 17274
rect 37936 16918 38148 16946
rect 38476 16992 38528 16998
rect 38476 16934 38528 16940
rect 37832 16584 37884 16590
rect 37832 16526 37884 16532
rect 37464 16448 37516 16454
rect 37464 16390 37516 16396
rect 37476 16046 37504 16390
rect 37844 16114 37872 16526
rect 37832 16108 37884 16114
rect 37832 16050 37884 16056
rect 37464 16040 37516 16046
rect 37462 16008 37464 16017
rect 37516 16008 37518 16017
rect 37462 15943 37518 15952
rect 37832 15904 37884 15910
rect 37832 15846 37884 15852
rect 37556 15428 37608 15434
rect 37556 15370 37608 15376
rect 37372 15360 37424 15366
rect 37372 15302 37424 15308
rect 37568 15162 37596 15370
rect 37556 15156 37608 15162
rect 37556 15098 37608 15104
rect 37464 14952 37516 14958
rect 37464 14894 37516 14900
rect 37280 14476 37332 14482
rect 37280 14418 37332 14424
rect 37292 13938 37320 14418
rect 37004 13932 37056 13938
rect 37004 13874 37056 13880
rect 37280 13932 37332 13938
rect 37280 13874 37332 13880
rect 36912 13252 36964 13258
rect 36912 13194 36964 13200
rect 36820 12844 36872 12850
rect 36820 12786 36872 12792
rect 36924 9654 36952 13194
rect 37016 12850 37044 13874
rect 37096 13796 37148 13802
rect 37096 13738 37148 13744
rect 37108 13394 37136 13738
rect 37188 13456 37240 13462
rect 37188 13398 37240 13404
rect 37096 13388 37148 13394
rect 37096 13330 37148 13336
rect 37004 12844 37056 12850
rect 37004 12786 37056 12792
rect 37096 12776 37148 12782
rect 37096 12718 37148 12724
rect 37108 10810 37136 12718
rect 37200 10996 37228 13398
rect 37476 13258 37504 14894
rect 37844 14822 37872 15846
rect 37936 15026 37964 16918
rect 38488 16726 38516 16934
rect 38476 16720 38528 16726
rect 38476 16662 38528 16668
rect 38292 16516 38344 16522
rect 38292 16458 38344 16464
rect 38384 16516 38436 16522
rect 38384 16458 38436 16464
rect 38200 16108 38252 16114
rect 38200 16050 38252 16056
rect 38108 15904 38160 15910
rect 38108 15846 38160 15852
rect 38120 15026 38148 15846
rect 38212 15570 38240 16050
rect 38304 15706 38332 16458
rect 38292 15700 38344 15706
rect 38292 15642 38344 15648
rect 38200 15564 38252 15570
rect 38200 15506 38252 15512
rect 37924 15020 37976 15026
rect 37924 14962 37976 14968
rect 38108 15020 38160 15026
rect 38108 14962 38160 14968
rect 38396 14958 38424 16458
rect 38488 16454 38516 16662
rect 38476 16448 38528 16454
rect 38476 16390 38528 16396
rect 38580 16114 38608 18226
rect 38660 18148 38712 18154
rect 38660 18090 38712 18096
rect 38672 17882 38700 18090
rect 38764 18086 38792 18244
rect 38856 18222 38884 19654
rect 38948 19378 38976 19654
rect 38936 19372 38988 19378
rect 38936 19314 38988 19320
rect 38936 18284 38988 18290
rect 38936 18226 38988 18232
rect 38844 18216 38896 18222
rect 38948 18193 38976 18226
rect 38844 18158 38896 18164
rect 38934 18184 38990 18193
rect 38934 18119 38990 18128
rect 38752 18080 38804 18086
rect 38752 18022 38804 18028
rect 38660 17876 38712 17882
rect 38660 17818 38712 17824
rect 38764 17678 38792 18022
rect 38752 17672 38804 17678
rect 38752 17614 38804 17620
rect 38936 17332 38988 17338
rect 38936 17274 38988 17280
rect 38750 17232 38806 17241
rect 38750 17167 38752 17176
rect 38804 17167 38806 17176
rect 38752 17138 38804 17144
rect 38660 16992 38712 16998
rect 38660 16934 38712 16940
rect 38672 16794 38700 16934
rect 38660 16788 38712 16794
rect 38660 16730 38712 16736
rect 38948 16590 38976 17274
rect 38936 16584 38988 16590
rect 38750 16552 38806 16561
rect 38936 16526 38988 16532
rect 38750 16487 38752 16496
rect 38804 16487 38806 16496
rect 38844 16516 38896 16522
rect 38752 16458 38804 16464
rect 38844 16458 38896 16464
rect 38660 16448 38712 16454
rect 38660 16390 38712 16396
rect 38672 16250 38700 16390
rect 38660 16244 38712 16250
rect 38660 16186 38712 16192
rect 38672 16114 38700 16186
rect 38568 16108 38620 16114
rect 38568 16050 38620 16056
rect 38660 16108 38712 16114
rect 38660 16050 38712 16056
rect 38580 15994 38608 16050
rect 38856 16046 38884 16458
rect 39040 16266 39068 20538
rect 39304 20460 39356 20466
rect 39304 20402 39356 20408
rect 39120 20392 39172 20398
rect 39120 20334 39172 20340
rect 39132 19786 39160 20334
rect 39120 19780 39172 19786
rect 39120 19722 39172 19728
rect 39120 19372 39172 19378
rect 39120 19314 39172 19320
rect 39212 19372 39264 19378
rect 39212 19314 39264 19320
rect 39132 18193 39160 19314
rect 39224 18970 39252 19314
rect 39212 18964 39264 18970
rect 39212 18906 39264 18912
rect 39210 18320 39266 18329
rect 39210 18255 39212 18264
rect 39264 18255 39266 18264
rect 39212 18226 39264 18232
rect 39118 18184 39174 18193
rect 39118 18119 39174 18128
rect 38948 16250 39068 16266
rect 38936 16244 39068 16250
rect 38988 16238 39068 16244
rect 38936 16186 38988 16192
rect 39028 16176 39080 16182
rect 39028 16118 39080 16124
rect 38844 16040 38896 16046
rect 38580 15966 38700 15994
rect 38844 15982 38896 15988
rect 38568 15904 38620 15910
rect 38568 15846 38620 15852
rect 38580 15162 38608 15846
rect 38672 15638 38700 15966
rect 39040 15706 39068 16118
rect 39028 15700 39080 15706
rect 39028 15642 39080 15648
rect 38660 15632 38712 15638
rect 38660 15574 38712 15580
rect 39040 15502 39068 15642
rect 39132 15638 39160 18119
rect 39224 17814 39252 18226
rect 39212 17808 39264 17814
rect 39212 17750 39264 17756
rect 39316 17338 39344 20402
rect 39408 17864 39436 22066
rect 39488 20392 39540 20398
rect 39488 20334 39540 20340
rect 39500 19854 39528 20334
rect 39488 19848 39540 19854
rect 39488 19790 39540 19796
rect 39488 19168 39540 19174
rect 39488 19110 39540 19116
rect 39592 19122 39620 22066
rect 39684 21418 39712 23695
rect 39776 23186 39804 23734
rect 39764 23180 39816 23186
rect 39764 23122 39816 23128
rect 39960 23118 39988 23854
rect 40040 23860 40092 23866
rect 40040 23802 40092 23808
rect 40144 23712 40172 24550
rect 40512 24313 40540 24550
rect 40498 24304 40554 24313
rect 40498 24239 40554 24248
rect 40500 23792 40552 23798
rect 40052 23684 40172 23712
rect 40498 23760 40500 23769
rect 40552 23760 40554 23769
rect 40498 23695 40554 23704
rect 39948 23112 40000 23118
rect 39948 23054 40000 23060
rect 40052 23066 40080 23684
rect 40132 23588 40184 23594
rect 40132 23530 40184 23536
rect 40144 23322 40172 23530
rect 40224 23520 40276 23526
rect 40224 23462 40276 23468
rect 40132 23316 40184 23322
rect 40132 23258 40184 23264
rect 40144 23186 40172 23258
rect 40132 23180 40184 23186
rect 40132 23122 40184 23128
rect 40052 23038 40172 23066
rect 39764 22976 39816 22982
rect 39764 22918 39816 22924
rect 39776 22438 39804 22918
rect 39948 22636 40000 22642
rect 39948 22578 40000 22584
rect 39764 22432 39816 22438
rect 39762 22400 39764 22409
rect 39816 22400 39818 22409
rect 39762 22335 39818 22344
rect 39672 21412 39724 21418
rect 39672 21354 39724 21360
rect 39856 20800 39908 20806
rect 39856 20742 39908 20748
rect 39868 20534 39896 20742
rect 39856 20528 39908 20534
rect 39856 20470 39908 20476
rect 39500 18902 39528 19110
rect 39592 19094 39896 19122
rect 39868 18970 39896 19094
rect 39764 18964 39816 18970
rect 39764 18906 39816 18912
rect 39856 18964 39908 18970
rect 39856 18906 39908 18912
rect 39488 18896 39540 18902
rect 39488 18838 39540 18844
rect 39500 18222 39528 18838
rect 39776 18766 39804 18906
rect 39764 18760 39816 18766
rect 39764 18702 39816 18708
rect 39580 18692 39632 18698
rect 39580 18634 39632 18640
rect 39592 18290 39620 18634
rect 39776 18290 39804 18702
rect 39580 18284 39632 18290
rect 39580 18226 39632 18232
rect 39672 18284 39724 18290
rect 39672 18226 39724 18232
rect 39764 18284 39816 18290
rect 39764 18226 39816 18232
rect 39488 18216 39540 18222
rect 39488 18158 39540 18164
rect 39408 17836 39528 17864
rect 39304 17332 39356 17338
rect 39304 17274 39356 17280
rect 39210 16688 39266 16697
rect 39210 16623 39266 16632
rect 39120 15632 39172 15638
rect 39120 15574 39172 15580
rect 39028 15496 39080 15502
rect 39028 15438 39080 15444
rect 38568 15156 38620 15162
rect 38568 15098 38620 15104
rect 39040 15026 39068 15438
rect 39224 15434 39252 16623
rect 39316 15434 39344 17274
rect 39396 17060 39448 17066
rect 39396 17002 39448 17008
rect 39408 16454 39436 17002
rect 39396 16448 39448 16454
rect 39396 16390 39448 16396
rect 39408 15978 39436 16390
rect 39500 16182 39528 17836
rect 39684 16454 39712 18226
rect 39868 18170 39896 18906
rect 39776 18142 39896 18170
rect 39776 17338 39804 18142
rect 39960 17882 39988 22578
rect 40040 21004 40092 21010
rect 40040 20946 40092 20952
rect 40052 19378 40080 20946
rect 40040 19372 40092 19378
rect 40040 19314 40092 19320
rect 40144 18426 40172 23038
rect 40236 20602 40264 23462
rect 40604 23322 40632 25638
rect 40774 24168 40830 24177
rect 40774 24103 40776 24112
rect 40828 24103 40830 24112
rect 40776 24074 40828 24080
rect 40682 24032 40738 24041
rect 40682 23967 40738 23976
rect 40592 23316 40644 23322
rect 40592 23258 40644 23264
rect 40408 22024 40460 22030
rect 40460 21984 40540 22012
rect 40408 21966 40460 21972
rect 40316 21412 40368 21418
rect 40316 21354 40368 21360
rect 40224 20596 40276 20602
rect 40224 20538 40276 20544
rect 40224 19372 40276 19378
rect 40224 19314 40276 19320
rect 40040 18420 40092 18426
rect 40040 18362 40092 18368
rect 40132 18420 40184 18426
rect 40132 18362 40184 18368
rect 39948 17876 40000 17882
rect 39948 17818 40000 17824
rect 40052 17746 40080 18362
rect 40132 18284 40184 18290
rect 40132 18226 40184 18232
rect 40040 17740 40092 17746
rect 40040 17682 40092 17688
rect 39856 17604 39908 17610
rect 39856 17546 39908 17552
rect 39764 17332 39816 17338
rect 39764 17274 39816 17280
rect 39762 17232 39818 17241
rect 39762 17167 39764 17176
rect 39816 17167 39818 17176
rect 39764 17138 39816 17144
rect 39672 16448 39724 16454
rect 39672 16390 39724 16396
rect 39868 16250 39896 17546
rect 40144 17542 40172 18226
rect 40236 18222 40264 19314
rect 40328 18290 40356 21354
rect 40512 20942 40540 21984
rect 40592 21072 40644 21078
rect 40592 21014 40644 21020
rect 40500 20936 40552 20942
rect 40500 20878 40552 20884
rect 40512 20398 40540 20878
rect 40500 20392 40552 20398
rect 40500 20334 40552 20340
rect 40512 19514 40540 20334
rect 40500 19508 40552 19514
rect 40500 19450 40552 19456
rect 40408 19236 40460 19242
rect 40408 19178 40460 19184
rect 40316 18284 40368 18290
rect 40316 18226 40368 18232
rect 40224 18216 40276 18222
rect 40224 18158 40276 18164
rect 40132 17536 40184 17542
rect 40132 17478 40184 17484
rect 40420 17338 40448 19178
rect 40500 18760 40552 18766
rect 40500 18702 40552 18708
rect 40512 18290 40540 18702
rect 40500 18284 40552 18290
rect 40500 18226 40552 18232
rect 40604 17762 40632 21014
rect 40696 19446 40724 23967
rect 40788 22094 40816 24074
rect 40880 24041 40908 25910
rect 41972 25832 42024 25838
rect 41972 25774 42024 25780
rect 41512 25492 41564 25498
rect 41512 25434 41564 25440
rect 41236 25356 41288 25362
rect 41288 25316 41460 25344
rect 41236 25298 41288 25304
rect 41432 25226 41460 25316
rect 41420 25220 41472 25226
rect 41420 25162 41472 25168
rect 40960 25152 41012 25158
rect 40960 25094 41012 25100
rect 40972 24818 41000 25094
rect 41432 24818 41460 25162
rect 41524 25158 41552 25434
rect 41984 25401 42012 25774
rect 41970 25392 42026 25401
rect 42076 25362 42104 26386
rect 42156 26240 42208 26246
rect 42156 26182 42208 26188
rect 41970 25327 41972 25336
rect 42024 25327 42026 25336
rect 42064 25356 42116 25362
rect 41972 25298 42024 25304
rect 42064 25298 42116 25304
rect 42062 25256 42118 25265
rect 42062 25191 42118 25200
rect 41512 25152 41564 25158
rect 41512 25094 41564 25100
rect 40960 24812 41012 24818
rect 40960 24754 41012 24760
rect 41420 24812 41472 24818
rect 41420 24754 41472 24760
rect 41788 24812 41840 24818
rect 41788 24754 41840 24760
rect 41328 24744 41380 24750
rect 41328 24686 41380 24692
rect 41340 24206 41368 24686
rect 41800 24614 41828 24754
rect 41788 24608 41840 24614
rect 41788 24550 41840 24556
rect 41512 24336 41564 24342
rect 41512 24278 41564 24284
rect 41328 24200 41380 24206
rect 41328 24142 41380 24148
rect 41420 24132 41472 24138
rect 41420 24074 41472 24080
rect 40866 24032 40922 24041
rect 40922 23990 41000 24018
rect 40866 23967 40922 23976
rect 40788 22066 40908 22094
rect 40880 21078 40908 22066
rect 40868 21072 40920 21078
rect 40868 21014 40920 21020
rect 40972 19666 41000 23990
rect 41432 23118 41460 24074
rect 41524 23662 41552 24278
rect 41512 23656 41564 23662
rect 41512 23598 41564 23604
rect 41604 23248 41656 23254
rect 41602 23216 41604 23225
rect 41656 23216 41658 23225
rect 41602 23151 41658 23160
rect 41696 23180 41748 23186
rect 41616 23118 41644 23151
rect 41696 23122 41748 23128
rect 41420 23112 41472 23118
rect 41420 23054 41472 23060
rect 41604 23112 41656 23118
rect 41604 23054 41656 23060
rect 41604 22636 41656 22642
rect 41604 22578 41656 22584
rect 41512 22568 41564 22574
rect 41512 22510 41564 22516
rect 41144 22432 41196 22438
rect 41144 22374 41196 22380
rect 41156 22234 41184 22374
rect 41144 22228 41196 22234
rect 41144 22170 41196 22176
rect 41524 21554 41552 22510
rect 41616 21894 41644 22578
rect 41708 22094 41736 23122
rect 42076 22094 42104 25191
rect 42168 24818 42196 26182
rect 42352 25906 42380 26862
rect 42444 26450 42472 28698
rect 42432 26444 42484 26450
rect 42432 26386 42484 26392
rect 42536 26042 42564 29582
rect 42800 29572 42852 29578
rect 42800 29514 42852 29520
rect 42812 28558 42840 29514
rect 43364 29510 43392 30262
rect 44732 30184 44784 30190
rect 44732 30126 44784 30132
rect 44180 29708 44232 29714
rect 44180 29650 44232 29656
rect 43996 29572 44048 29578
rect 43996 29514 44048 29520
rect 43352 29504 43404 29510
rect 43352 29446 43404 29452
rect 42892 29300 42944 29306
rect 42892 29242 42944 29248
rect 42800 28552 42852 28558
rect 42800 28494 42852 28500
rect 42708 28212 42760 28218
rect 42708 28154 42760 28160
rect 42720 28082 42748 28154
rect 42798 28112 42854 28121
rect 42708 28076 42760 28082
rect 42904 28082 42932 29242
rect 42984 29232 43036 29238
rect 42984 29174 43036 29180
rect 42996 28744 43024 29174
rect 43076 28756 43128 28762
rect 42996 28716 43076 28744
rect 42798 28047 42800 28056
rect 42708 28018 42760 28024
rect 42852 28047 42854 28056
rect 42892 28076 42944 28082
rect 42800 28018 42852 28024
rect 42892 28018 42944 28024
rect 42616 27872 42668 27878
rect 42616 27814 42668 27820
rect 42708 27872 42760 27878
rect 42708 27814 42760 27820
rect 42524 26036 42576 26042
rect 42524 25978 42576 25984
rect 42340 25900 42392 25906
rect 42340 25842 42392 25848
rect 42352 25362 42380 25842
rect 42628 25702 42656 27814
rect 42720 26926 42748 27814
rect 42812 27470 42840 28018
rect 42996 27946 43024 28716
rect 43076 28698 43128 28704
rect 43168 28688 43220 28694
rect 43168 28630 43220 28636
rect 43180 28558 43208 28630
rect 43168 28552 43220 28558
rect 43260 28552 43312 28558
rect 43168 28494 43220 28500
rect 43258 28520 43260 28529
rect 43312 28520 43314 28529
rect 43076 28076 43128 28082
rect 43076 28018 43128 28024
rect 42984 27940 43036 27946
rect 42984 27882 43036 27888
rect 42892 27600 42944 27606
rect 42892 27542 42944 27548
rect 42800 27464 42852 27470
rect 42800 27406 42852 27412
rect 42812 27130 42840 27406
rect 42800 27124 42852 27130
rect 42800 27066 42852 27072
rect 42708 26920 42760 26926
rect 42708 26862 42760 26868
rect 42708 26784 42760 26790
rect 42708 26726 42760 26732
rect 42720 25974 42748 26726
rect 42904 26518 42932 27542
rect 42996 27470 43024 27882
rect 43088 27674 43116 28018
rect 43076 27668 43128 27674
rect 43076 27610 43128 27616
rect 43180 27470 43208 28494
rect 43258 28455 43314 28464
rect 42984 27464 43036 27470
rect 42984 27406 43036 27412
rect 43168 27464 43220 27470
rect 43168 27406 43220 27412
rect 43364 27418 43392 29446
rect 43904 29232 43956 29238
rect 43904 29174 43956 29180
rect 43720 29164 43772 29170
rect 43720 29106 43772 29112
rect 43536 29096 43588 29102
rect 43536 29038 43588 29044
rect 43444 28960 43496 28966
rect 43444 28902 43496 28908
rect 43456 28558 43484 28902
rect 43444 28552 43496 28558
rect 43444 28494 43496 28500
rect 43548 27538 43576 29038
rect 43732 28558 43760 29106
rect 43812 29028 43864 29034
rect 43812 28970 43864 28976
rect 43824 28558 43852 28970
rect 43720 28552 43772 28558
rect 43720 28494 43772 28500
rect 43812 28552 43864 28558
rect 43812 28494 43864 28500
rect 43732 28218 43760 28494
rect 43720 28212 43772 28218
rect 43720 28154 43772 28160
rect 43628 27872 43680 27878
rect 43628 27814 43680 27820
rect 43640 27674 43668 27814
rect 43628 27668 43680 27674
rect 43628 27610 43680 27616
rect 43536 27532 43588 27538
rect 43536 27474 43588 27480
rect 43364 27390 43576 27418
rect 42892 26512 42944 26518
rect 42892 26454 42944 26460
rect 43444 26512 43496 26518
rect 43444 26454 43496 26460
rect 42892 26376 42944 26382
rect 42892 26318 42944 26324
rect 42904 26042 42932 26318
rect 43352 26308 43404 26314
rect 43352 26250 43404 26256
rect 42892 26036 42944 26042
rect 42892 25978 42944 25984
rect 42708 25968 42760 25974
rect 42708 25910 42760 25916
rect 42616 25696 42668 25702
rect 42616 25638 42668 25644
rect 42340 25356 42392 25362
rect 42260 25316 42340 25344
rect 42156 24812 42208 24818
rect 42156 24754 42208 24760
rect 42168 24206 42196 24754
rect 42156 24200 42208 24206
rect 42156 24142 42208 24148
rect 42260 23225 42288 25316
rect 42340 25298 42392 25304
rect 42524 25288 42576 25294
rect 42524 25230 42576 25236
rect 42432 24948 42484 24954
rect 42432 24890 42484 24896
rect 42444 24614 42472 24890
rect 42536 24800 42564 25230
rect 42628 25226 42656 25638
rect 42720 25498 42748 25910
rect 42708 25492 42760 25498
rect 42708 25434 42760 25440
rect 42800 25424 42852 25430
rect 42706 25392 42762 25401
rect 42762 25372 42800 25378
rect 42762 25366 42852 25372
rect 42762 25350 42840 25366
rect 42706 25327 42762 25336
rect 42904 25294 42932 25978
rect 43364 25498 43392 26250
rect 43456 25838 43484 26454
rect 43444 25832 43496 25838
rect 43444 25774 43496 25780
rect 43352 25492 43404 25498
rect 43272 25452 43352 25480
rect 42892 25288 42944 25294
rect 42892 25230 42944 25236
rect 42616 25220 42668 25226
rect 42616 25162 42668 25168
rect 42708 25220 42760 25226
rect 42708 25162 42760 25168
rect 42720 24954 42748 25162
rect 42708 24948 42760 24954
rect 42708 24890 42760 24896
rect 42708 24812 42760 24818
rect 42536 24772 42708 24800
rect 42708 24754 42760 24760
rect 42432 24608 42484 24614
rect 42432 24550 42484 24556
rect 42444 24138 42472 24550
rect 42720 24410 42748 24754
rect 42904 24750 42932 25230
rect 42892 24744 42944 24750
rect 42892 24686 42944 24692
rect 42984 24744 43036 24750
rect 42984 24686 43036 24692
rect 42800 24676 42852 24682
rect 42800 24618 42852 24624
rect 42708 24404 42760 24410
rect 42708 24346 42760 24352
rect 42524 24336 42576 24342
rect 42524 24278 42576 24284
rect 42432 24132 42484 24138
rect 42432 24074 42484 24080
rect 42246 23216 42302 23225
rect 42444 23186 42472 24074
rect 42536 23798 42564 24278
rect 42524 23792 42576 23798
rect 42524 23734 42576 23740
rect 42720 23730 42748 24346
rect 42812 23730 42840 24618
rect 42904 23798 42932 24686
rect 42996 24614 43024 24686
rect 42984 24608 43036 24614
rect 42984 24550 43036 24556
rect 42996 24449 43024 24550
rect 42982 24440 43038 24449
rect 42982 24375 43038 24384
rect 43272 24138 43300 25452
rect 43352 25434 43404 25440
rect 43350 24576 43406 24585
rect 43548 24562 43576 27390
rect 43640 26994 43668 27610
rect 43732 27538 43760 28154
rect 43720 27532 43772 27538
rect 43720 27474 43772 27480
rect 43824 27130 43852 28494
rect 43916 28422 43944 29174
rect 44008 28642 44036 29514
rect 44192 29510 44220 29650
rect 44364 29640 44416 29646
rect 44364 29582 44416 29588
rect 44180 29504 44232 29510
rect 44180 29446 44232 29452
rect 44192 29170 44220 29446
rect 44180 29164 44232 29170
rect 44180 29106 44232 29112
rect 44376 29102 44404 29582
rect 44744 29170 44772 30126
rect 49700 29640 49752 29646
rect 49700 29582 49752 29588
rect 45376 29572 45428 29578
rect 45376 29514 45428 29520
rect 47124 29572 47176 29578
rect 47124 29514 47176 29520
rect 45388 29306 45416 29514
rect 47136 29306 47164 29514
rect 47400 29504 47452 29510
rect 47400 29446 47452 29452
rect 45376 29300 45428 29306
rect 45376 29242 45428 29248
rect 47124 29300 47176 29306
rect 47124 29242 47176 29248
rect 44732 29164 44784 29170
rect 44732 29106 44784 29112
rect 46112 29164 46164 29170
rect 46112 29106 46164 29112
rect 44364 29096 44416 29102
rect 44364 29038 44416 29044
rect 44376 28694 44404 29038
rect 44364 28688 44416 28694
rect 44008 28614 44128 28642
rect 44364 28630 44416 28636
rect 43996 28552 44048 28558
rect 43996 28494 44048 28500
rect 43904 28416 43956 28422
rect 43904 28358 43956 28364
rect 44008 28082 44036 28494
rect 43996 28076 44048 28082
rect 43996 28018 44048 28024
rect 43904 27668 43956 27674
rect 43904 27610 43956 27616
rect 43812 27124 43864 27130
rect 43812 27066 43864 27072
rect 43916 26994 43944 27610
rect 44008 27402 44036 28018
rect 44100 27538 44128 28614
rect 44744 28490 44772 29106
rect 45928 29096 45980 29102
rect 45928 29038 45980 29044
rect 45192 28756 45244 28762
rect 45192 28698 45244 28704
rect 44824 28688 44876 28694
rect 44824 28630 44876 28636
rect 44180 28484 44232 28490
rect 44732 28484 44784 28490
rect 44180 28426 44232 28432
rect 44652 28444 44732 28472
rect 44192 28218 44220 28426
rect 44272 28416 44324 28422
rect 44272 28358 44324 28364
rect 44180 28212 44232 28218
rect 44180 28154 44232 28160
rect 44284 27674 44312 28358
rect 44652 28014 44680 28444
rect 44732 28426 44784 28432
rect 44836 28014 44864 28630
rect 45204 28558 45232 28698
rect 45192 28552 45244 28558
rect 45284 28552 45336 28558
rect 45192 28494 45244 28500
rect 45282 28520 45284 28529
rect 45652 28552 45704 28558
rect 45336 28520 45338 28529
rect 45652 28494 45704 28500
rect 45282 28455 45338 28464
rect 44916 28212 44968 28218
rect 44916 28154 44968 28160
rect 44640 28008 44692 28014
rect 44640 27950 44692 27956
rect 44732 28008 44784 28014
rect 44732 27950 44784 27956
rect 44824 28008 44876 28014
rect 44824 27950 44876 27956
rect 44744 27674 44772 27950
rect 44272 27668 44324 27674
rect 44272 27610 44324 27616
rect 44732 27668 44784 27674
rect 44732 27610 44784 27616
rect 44088 27532 44140 27538
rect 44088 27474 44140 27480
rect 43996 27396 44048 27402
rect 43996 27338 44048 27344
rect 43628 26988 43680 26994
rect 43628 26930 43680 26936
rect 43904 26988 43956 26994
rect 43904 26930 43956 26936
rect 43628 26784 43680 26790
rect 43628 26726 43680 26732
rect 43640 26246 43668 26726
rect 44180 26580 44232 26586
rect 44180 26522 44232 26528
rect 43628 26240 43680 26246
rect 43628 26182 43680 26188
rect 43812 25968 43864 25974
rect 43810 25936 43812 25945
rect 43864 25936 43866 25945
rect 44192 25906 44220 26522
rect 44928 26314 44956 28154
rect 45664 27946 45692 28494
rect 45940 27946 45968 29038
rect 46124 28762 46152 29106
rect 46112 28756 46164 28762
rect 46112 28698 46164 28704
rect 45652 27940 45704 27946
rect 45928 27940 45980 27946
rect 45652 27882 45704 27888
rect 45756 27900 45928 27928
rect 45100 27328 45152 27334
rect 45100 27270 45152 27276
rect 44916 26308 44968 26314
rect 44916 26250 44968 26256
rect 43810 25871 43866 25880
rect 44180 25900 44232 25906
rect 44180 25842 44232 25848
rect 43812 25696 43864 25702
rect 43812 25638 43864 25644
rect 43824 25498 43852 25638
rect 43812 25492 43864 25498
rect 43812 25434 43864 25440
rect 43996 25492 44048 25498
rect 43996 25434 44048 25440
rect 43824 25362 43852 25434
rect 43812 25356 43864 25362
rect 43812 25298 43864 25304
rect 43628 25288 43680 25294
rect 43628 25230 43680 25236
rect 43640 24682 43668 25230
rect 44008 25158 44036 25434
rect 43996 25152 44048 25158
rect 43996 25094 44048 25100
rect 43812 24744 43864 24750
rect 43810 24712 43812 24721
rect 43864 24712 43866 24721
rect 43628 24676 43680 24682
rect 43810 24647 43866 24656
rect 43628 24618 43680 24624
rect 43720 24608 43772 24614
rect 43548 24534 43668 24562
rect 43720 24550 43772 24556
rect 43350 24511 43406 24520
rect 42984 24132 43036 24138
rect 42984 24074 43036 24080
rect 43260 24132 43312 24138
rect 43260 24074 43312 24080
rect 42996 24041 43024 24074
rect 43168 24064 43220 24070
rect 42982 24032 43038 24041
rect 43038 24012 43168 24018
rect 43038 24006 43220 24012
rect 43038 23990 43208 24006
rect 42982 23967 43038 23976
rect 43166 23896 43222 23905
rect 43166 23831 43222 23840
rect 43180 23798 43208 23831
rect 42892 23792 42944 23798
rect 42892 23734 42944 23740
rect 43168 23792 43220 23798
rect 43168 23734 43220 23740
rect 42708 23724 42760 23730
rect 42708 23666 42760 23672
rect 42800 23724 42852 23730
rect 42800 23666 42852 23672
rect 42246 23151 42302 23160
rect 42432 23180 42484 23186
rect 42154 23080 42210 23089
rect 42154 23015 42156 23024
rect 42208 23015 42210 23024
rect 42156 22986 42208 22992
rect 42260 22982 42288 23151
rect 42432 23122 42484 23128
rect 42812 23118 42840 23666
rect 43272 23662 43300 24074
rect 43260 23656 43312 23662
rect 43260 23598 43312 23604
rect 42800 23112 42852 23118
rect 42800 23054 42852 23060
rect 42340 23044 42392 23050
rect 42340 22986 42392 22992
rect 42248 22976 42300 22982
rect 42248 22918 42300 22924
rect 42352 22778 42380 22986
rect 42340 22772 42392 22778
rect 42340 22714 42392 22720
rect 42708 22772 42760 22778
rect 42708 22714 42760 22720
rect 42248 22636 42300 22642
rect 42248 22578 42300 22584
rect 42616 22636 42668 22642
rect 42616 22578 42668 22584
rect 42156 22432 42208 22438
rect 42156 22374 42208 22380
rect 41708 22066 41828 22094
rect 41604 21888 41656 21894
rect 41604 21830 41656 21836
rect 41512 21548 41564 21554
rect 41512 21490 41564 21496
rect 41236 21412 41288 21418
rect 41236 21354 41288 21360
rect 41248 20262 41276 21354
rect 41328 20392 41380 20398
rect 41328 20334 41380 20340
rect 41236 20256 41288 20262
rect 41236 20198 41288 20204
rect 41248 20058 41276 20198
rect 41340 20058 41368 20334
rect 41236 20052 41288 20058
rect 41236 19994 41288 20000
rect 41328 20052 41380 20058
rect 41328 19994 41380 20000
rect 41524 19854 41552 21490
rect 41512 19848 41564 19854
rect 41512 19790 41564 19796
rect 41052 19780 41104 19786
rect 41052 19722 41104 19728
rect 40788 19638 41000 19666
rect 40684 19440 40736 19446
rect 40684 19382 40736 19388
rect 40684 18148 40736 18154
rect 40684 18090 40736 18096
rect 40696 17882 40724 18090
rect 40684 17876 40736 17882
rect 40684 17818 40736 17824
rect 40604 17734 40724 17762
rect 40592 17672 40644 17678
rect 40592 17614 40644 17620
rect 40604 17338 40632 17614
rect 40696 17338 40724 17734
rect 40408 17332 40460 17338
rect 40408 17274 40460 17280
rect 40592 17332 40644 17338
rect 40592 17274 40644 17280
rect 40684 17332 40736 17338
rect 40684 17274 40736 17280
rect 39948 17196 40000 17202
rect 40316 17196 40368 17202
rect 39948 17138 40000 17144
rect 40236 17156 40316 17184
rect 39960 16794 39988 17138
rect 40236 16833 40264 17156
rect 40316 17138 40368 17144
rect 40592 17128 40644 17134
rect 40592 17070 40644 17076
rect 40222 16824 40278 16833
rect 39948 16788 40000 16794
rect 40222 16759 40278 16768
rect 39948 16730 40000 16736
rect 40132 16720 40184 16726
rect 40052 16668 40132 16674
rect 40052 16662 40184 16668
rect 40052 16646 40172 16662
rect 40052 16590 40080 16646
rect 40040 16584 40092 16590
rect 40040 16526 40092 16532
rect 40132 16516 40184 16522
rect 40132 16458 40184 16464
rect 39856 16244 39908 16250
rect 39856 16186 39908 16192
rect 39488 16176 39540 16182
rect 39488 16118 39540 16124
rect 39396 15972 39448 15978
rect 39396 15914 39448 15920
rect 39500 15722 39528 16118
rect 39948 16108 40000 16114
rect 39948 16050 40000 16056
rect 39672 15972 39724 15978
rect 39672 15914 39724 15920
rect 39500 15694 39620 15722
rect 39488 15632 39540 15638
rect 39488 15574 39540 15580
rect 39212 15428 39264 15434
rect 39212 15370 39264 15376
rect 39304 15428 39356 15434
rect 39304 15370 39356 15376
rect 39500 15162 39528 15574
rect 39592 15366 39620 15694
rect 39580 15360 39632 15366
rect 39580 15302 39632 15308
rect 39684 15201 39712 15914
rect 39960 15609 39988 16050
rect 39946 15600 40002 15609
rect 39946 15535 40002 15544
rect 40040 15564 40092 15570
rect 40040 15506 40092 15512
rect 39854 15464 39910 15473
rect 39854 15399 39856 15408
rect 39908 15399 39910 15408
rect 39856 15370 39908 15376
rect 39670 15192 39726 15201
rect 39488 15156 39540 15162
rect 39670 15127 39672 15136
rect 39488 15098 39540 15104
rect 39724 15127 39726 15136
rect 39672 15098 39724 15104
rect 39028 15020 39080 15026
rect 39028 14962 39080 14968
rect 38384 14952 38436 14958
rect 38384 14894 38436 14900
rect 40052 14890 40080 15506
rect 40144 14958 40172 16458
rect 40236 15502 40264 16759
rect 40316 16448 40368 16454
rect 40316 16390 40368 16396
rect 40328 16182 40356 16390
rect 40316 16176 40368 16182
rect 40316 16118 40368 16124
rect 40408 16040 40460 16046
rect 40408 15982 40460 15988
rect 40316 15700 40368 15706
rect 40316 15642 40368 15648
rect 40328 15502 40356 15642
rect 40224 15496 40276 15502
rect 40224 15438 40276 15444
rect 40316 15496 40368 15502
rect 40316 15438 40368 15444
rect 40132 14952 40184 14958
rect 40328 14929 40356 15438
rect 40132 14894 40184 14900
rect 40314 14920 40370 14929
rect 40040 14884 40092 14890
rect 40040 14826 40092 14832
rect 37832 14816 37884 14822
rect 37832 14758 37884 14764
rect 38200 14816 38252 14822
rect 38200 14758 38252 14764
rect 38212 14618 38240 14758
rect 38200 14612 38252 14618
rect 38200 14554 38252 14560
rect 40144 14414 40172 14894
rect 40314 14855 40370 14864
rect 40420 14482 40448 15982
rect 40500 15428 40552 15434
rect 40500 15370 40552 15376
rect 40408 14476 40460 14482
rect 40408 14418 40460 14424
rect 40132 14408 40184 14414
rect 40132 14350 40184 14356
rect 38476 14272 38528 14278
rect 38476 14214 38528 14220
rect 40132 14272 40184 14278
rect 40132 14214 40184 14220
rect 37740 13864 37792 13870
rect 37740 13806 37792 13812
rect 37648 13796 37700 13802
rect 37648 13738 37700 13744
rect 37660 13530 37688 13738
rect 37752 13530 37780 13806
rect 37648 13524 37700 13530
rect 37648 13466 37700 13472
rect 37740 13524 37792 13530
rect 37740 13466 37792 13472
rect 37660 13326 37688 13466
rect 37648 13320 37700 13326
rect 37648 13262 37700 13268
rect 37464 13252 37516 13258
rect 37464 13194 37516 13200
rect 37556 13184 37608 13190
rect 37556 13126 37608 13132
rect 37568 11898 37596 13126
rect 37752 12986 37780 13466
rect 38488 13462 38516 14214
rect 38568 14000 38620 14006
rect 38568 13942 38620 13948
rect 37832 13456 37884 13462
rect 37832 13398 37884 13404
rect 38476 13456 38528 13462
rect 38476 13398 38528 13404
rect 37740 12980 37792 12986
rect 37740 12922 37792 12928
rect 37648 12844 37700 12850
rect 37648 12786 37700 12792
rect 37660 12753 37688 12786
rect 37740 12776 37792 12782
rect 37646 12744 37702 12753
rect 37740 12718 37792 12724
rect 37646 12679 37702 12688
rect 37660 12442 37688 12679
rect 37752 12442 37780 12718
rect 37648 12436 37700 12442
rect 37648 12378 37700 12384
rect 37740 12436 37792 12442
rect 37740 12378 37792 12384
rect 37844 12238 37872 13398
rect 37924 13252 37976 13258
rect 37924 13194 37976 13200
rect 37936 12714 37964 13194
rect 38488 12850 38516 13398
rect 38580 13326 38608 13942
rect 38936 13864 38988 13870
rect 38936 13806 38988 13812
rect 38948 13530 38976 13806
rect 38936 13524 38988 13530
rect 38936 13466 38988 13472
rect 40040 13456 40092 13462
rect 40040 13398 40092 13404
rect 38568 13320 38620 13326
rect 38568 13262 38620 13268
rect 39764 13320 39816 13326
rect 39764 13262 39816 13268
rect 38580 12986 38608 13262
rect 39212 13184 39264 13190
rect 39212 13126 39264 13132
rect 39224 12986 39252 13126
rect 38568 12980 38620 12986
rect 38568 12922 38620 12928
rect 39212 12980 39264 12986
rect 39212 12922 39264 12928
rect 38476 12844 38528 12850
rect 38476 12786 38528 12792
rect 38752 12844 38804 12850
rect 38752 12786 38804 12792
rect 38844 12844 38896 12850
rect 38844 12786 38896 12792
rect 39304 12844 39356 12850
rect 39304 12786 39356 12792
rect 39580 12844 39632 12850
rect 39580 12786 39632 12792
rect 38660 12776 38712 12782
rect 38660 12718 38712 12724
rect 37924 12708 37976 12714
rect 37924 12650 37976 12656
rect 37832 12232 37884 12238
rect 37832 12174 37884 12180
rect 37740 12096 37792 12102
rect 37740 12038 37792 12044
rect 37556 11892 37608 11898
rect 37556 11834 37608 11840
rect 37752 11762 37780 12038
rect 37936 11762 37964 12650
rect 38672 12374 38700 12718
rect 38660 12368 38712 12374
rect 38660 12310 38712 12316
rect 38764 12238 38792 12786
rect 38752 12232 38804 12238
rect 38672 12192 38752 12220
rect 38672 12102 38700 12192
rect 38752 12174 38804 12180
rect 38856 12102 38884 12786
rect 39120 12776 39172 12782
rect 38934 12744 38990 12753
rect 39316 12730 39344 12786
rect 39172 12724 39344 12730
rect 39120 12718 39344 12724
rect 39132 12702 39344 12718
rect 38934 12679 38990 12688
rect 38660 12096 38712 12102
rect 38660 12038 38712 12044
rect 38844 12096 38896 12102
rect 38844 12038 38896 12044
rect 38384 11892 38436 11898
rect 38384 11834 38436 11840
rect 38396 11801 38424 11834
rect 38382 11792 38438 11801
rect 37740 11756 37792 11762
rect 37740 11698 37792 11704
rect 37924 11756 37976 11762
rect 37924 11698 37976 11704
rect 38292 11756 38344 11762
rect 38382 11727 38438 11736
rect 38476 11756 38528 11762
rect 38292 11698 38344 11704
rect 38476 11698 38528 11704
rect 37832 11552 37884 11558
rect 37832 11494 37884 11500
rect 37844 11286 37872 11494
rect 37936 11354 37964 11698
rect 37924 11348 37976 11354
rect 37924 11290 37976 11296
rect 37832 11280 37884 11286
rect 37462 11248 37518 11257
rect 37832 11222 37884 11228
rect 38304 11234 38332 11698
rect 37462 11183 37518 11192
rect 37372 11008 37424 11014
rect 37200 10968 37320 10996
rect 37096 10804 37148 10810
rect 37096 10746 37148 10752
rect 37188 10736 37240 10742
rect 37188 10678 37240 10684
rect 37292 10690 37320 10968
rect 37372 10950 37424 10956
rect 37384 10810 37412 10950
rect 37372 10804 37424 10810
rect 37372 10746 37424 10752
rect 37200 10062 37228 10678
rect 37292 10662 37412 10690
rect 37004 10056 37056 10062
rect 37188 10056 37240 10062
rect 37004 9998 37056 10004
rect 37108 10016 37188 10044
rect 36912 9648 36964 9654
rect 36912 9590 36964 9596
rect 36820 9376 36872 9382
rect 36820 9318 36872 9324
rect 36636 9172 36688 9178
rect 36636 9114 36688 9120
rect 36728 9172 36780 9178
rect 36728 9114 36780 9120
rect 36740 9042 36768 9114
rect 36832 9042 36860 9318
rect 36728 9036 36780 9042
rect 36728 8978 36780 8984
rect 36820 9036 36872 9042
rect 36820 8978 36872 8984
rect 36464 8906 36584 8922
rect 36464 8900 36596 8906
rect 36464 8894 36544 8900
rect 36084 8560 36136 8566
rect 36084 8502 36136 8508
rect 32496 8492 32548 8498
rect 32496 8434 32548 8440
rect 35808 8492 35860 8498
rect 35808 8434 35860 8440
rect 35992 8492 36044 8498
rect 35992 8434 36044 8440
rect 32220 8424 32272 8430
rect 32220 8366 32272 8372
rect 32508 8294 32536 8434
rect 32496 8288 32548 8294
rect 32496 8230 32548 8236
rect 32680 8288 32732 8294
rect 32680 8230 32732 8236
rect 32128 8084 32180 8090
rect 32128 8026 32180 8032
rect 32508 8022 32536 8230
rect 32496 8016 32548 8022
rect 32496 7958 32548 7964
rect 32692 7886 32720 8230
rect 34934 8188 35242 8197
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8123 35242 8132
rect 33784 8016 33836 8022
rect 33784 7958 33836 7964
rect 32680 7880 32732 7886
rect 32680 7822 32732 7828
rect 31852 7540 31904 7546
rect 31852 7482 31904 7488
rect 32404 7336 32456 7342
rect 32404 7278 32456 7284
rect 32416 7002 32444 7278
rect 32404 6996 32456 7002
rect 32404 6938 32456 6944
rect 32692 6662 32720 7822
rect 32864 7472 32916 7478
rect 32864 7414 32916 7420
rect 32876 7002 32904 7414
rect 32956 7200 33008 7206
rect 32956 7142 33008 7148
rect 33140 7200 33192 7206
rect 33140 7142 33192 7148
rect 32864 6996 32916 7002
rect 32864 6938 32916 6944
rect 32968 6882 32996 7142
rect 33048 6928 33100 6934
rect 32876 6876 33048 6882
rect 32876 6870 33100 6876
rect 32876 6866 33088 6870
rect 32864 6860 33088 6866
rect 32916 6854 33088 6860
rect 32864 6802 32916 6808
rect 33152 6798 33180 7142
rect 33140 6792 33192 6798
rect 33140 6734 33192 6740
rect 32680 6656 32732 6662
rect 32680 6598 32732 6604
rect 31852 6316 31904 6322
rect 31852 6258 31904 6264
rect 31760 6248 31812 6254
rect 31760 6190 31812 6196
rect 31864 5914 31892 6258
rect 31852 5908 31904 5914
rect 31852 5850 31904 5856
rect 31864 5710 31892 5850
rect 31852 5704 31904 5710
rect 31852 5646 31904 5652
rect 31944 5568 31996 5574
rect 31944 5510 31996 5516
rect 31956 5370 31984 5510
rect 31944 5364 31996 5370
rect 31944 5306 31996 5312
rect 31668 5296 31720 5302
rect 31668 5238 31720 5244
rect 31392 5160 31444 5166
rect 31392 5102 31444 5108
rect 30748 4616 30800 4622
rect 30748 4558 30800 4564
rect 30760 3738 30788 4558
rect 31404 3738 31432 5102
rect 31484 4684 31536 4690
rect 31484 4626 31536 4632
rect 30748 3732 30800 3738
rect 30748 3674 30800 3680
rect 31392 3732 31444 3738
rect 31392 3674 31444 3680
rect 30656 2848 30708 2854
rect 30656 2790 30708 2796
rect 30392 2746 30604 2774
rect 29000 2644 29052 2650
rect 29000 2586 29052 2592
rect 29368 2644 29420 2650
rect 29368 2586 29420 2592
rect 30104 2644 30156 2650
rect 30104 2586 30156 2592
rect 30288 2644 30340 2650
rect 30288 2586 30340 2592
rect 29000 2508 29052 2514
rect 29000 2450 29052 2456
rect 23388 2440 23440 2446
rect 23388 2382 23440 2388
rect 22652 2372 22704 2378
rect 22652 2314 22704 2320
rect 23204 2304 23256 2310
rect 23204 2246 23256 2252
rect 23216 800 23244 2246
rect 29012 800 29040 2450
rect 30116 2446 30144 2586
rect 30300 2446 30328 2586
rect 30392 2582 30420 2746
rect 30380 2576 30432 2582
rect 30380 2518 30432 2524
rect 30760 2446 30788 3674
rect 31496 3602 31524 4626
rect 31484 3596 31536 3602
rect 31484 3538 31536 3544
rect 31496 2990 31524 3538
rect 32312 3460 32364 3466
rect 32312 3402 32364 3408
rect 32324 3126 32352 3402
rect 32404 3392 32456 3398
rect 32404 3334 32456 3340
rect 32416 3126 32444 3334
rect 32692 3194 32720 6598
rect 33796 6254 33824 7958
rect 35820 7954 35848 8434
rect 34428 7948 34480 7954
rect 34428 7890 34480 7896
rect 34520 7948 34572 7954
rect 34520 7890 34572 7896
rect 35808 7948 35860 7954
rect 35808 7890 35860 7896
rect 33876 7880 33928 7886
rect 33876 7822 33928 7828
rect 33888 7546 33916 7822
rect 33876 7540 33928 7546
rect 33876 7482 33928 7488
rect 34440 6798 34468 7890
rect 34532 6934 34560 7890
rect 35594 7644 35902 7653
rect 35594 7642 35600 7644
rect 35656 7642 35680 7644
rect 35736 7642 35760 7644
rect 35816 7642 35840 7644
rect 35896 7642 35902 7644
rect 35656 7590 35658 7642
rect 35838 7590 35840 7642
rect 35594 7588 35600 7590
rect 35656 7588 35680 7590
rect 35736 7588 35760 7590
rect 35816 7588 35840 7590
rect 35896 7588 35902 7590
rect 35594 7579 35902 7588
rect 34796 7472 34848 7478
rect 34796 7414 34848 7420
rect 34612 6996 34664 7002
rect 34612 6938 34664 6944
rect 34520 6928 34572 6934
rect 34520 6870 34572 6876
rect 33968 6792 34020 6798
rect 33968 6734 34020 6740
rect 34428 6792 34480 6798
rect 34428 6734 34480 6740
rect 33980 6254 34008 6734
rect 34520 6316 34572 6322
rect 34520 6258 34572 6264
rect 33784 6248 33836 6254
rect 33784 6190 33836 6196
rect 33968 6248 34020 6254
rect 33968 6190 34020 6196
rect 32772 5704 32824 5710
rect 32772 5646 32824 5652
rect 32784 4690 32812 5646
rect 33324 5636 33376 5642
rect 33324 5578 33376 5584
rect 32864 5568 32916 5574
rect 32864 5510 32916 5516
rect 32772 4684 32824 4690
rect 32772 4626 32824 4632
rect 32876 4622 32904 5510
rect 33336 5370 33364 5578
rect 33324 5364 33376 5370
rect 33324 5306 33376 5312
rect 33796 5166 33824 6190
rect 34532 5914 34560 6258
rect 34520 5908 34572 5914
rect 34520 5850 34572 5856
rect 33784 5160 33836 5166
rect 33784 5102 33836 5108
rect 34152 5160 34204 5166
rect 34152 5102 34204 5108
rect 32864 4616 32916 4622
rect 32864 4558 32916 4564
rect 32876 3466 32904 4558
rect 32864 3460 32916 3466
rect 32864 3402 32916 3408
rect 32680 3188 32732 3194
rect 32680 3130 32732 3136
rect 32876 3126 32904 3402
rect 33796 3194 33824 5102
rect 34164 4826 34192 5102
rect 34624 4826 34652 6938
rect 34808 6390 34836 7414
rect 35440 7336 35492 7342
rect 35440 7278 35492 7284
rect 35348 7200 35400 7206
rect 35348 7142 35400 7148
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 35360 6866 35388 7142
rect 35348 6860 35400 6866
rect 35348 6802 35400 6808
rect 35452 6730 35480 7278
rect 36004 6730 36032 8434
rect 36360 8356 36412 8362
rect 36360 8298 36412 8304
rect 36268 8288 36320 8294
rect 36268 8230 36320 8236
rect 36280 8022 36308 8230
rect 36268 8016 36320 8022
rect 36268 7958 36320 7964
rect 36176 7200 36228 7206
rect 36176 7142 36228 7148
rect 36188 6798 36216 7142
rect 36176 6792 36228 6798
rect 36176 6734 36228 6740
rect 35440 6724 35492 6730
rect 35440 6666 35492 6672
rect 35992 6724 36044 6730
rect 35992 6666 36044 6672
rect 36280 6662 36308 7958
rect 36372 7886 36400 8298
rect 36360 7880 36412 7886
rect 36360 7822 36412 7828
rect 36360 7336 36412 7342
rect 36464 7290 36492 8894
rect 36544 8842 36596 8848
rect 36728 8832 36780 8838
rect 36728 8774 36780 8780
rect 36740 8498 36768 8774
rect 36636 8492 36688 8498
rect 36636 8434 36688 8440
rect 36728 8492 36780 8498
rect 36728 8434 36780 8440
rect 36648 7954 36676 8434
rect 36912 8424 36964 8430
rect 36912 8366 36964 8372
rect 36636 7948 36688 7954
rect 36636 7890 36688 7896
rect 36648 7546 36676 7890
rect 36636 7540 36688 7546
rect 36636 7482 36688 7488
rect 36544 7404 36596 7410
rect 36544 7346 36596 7352
rect 36412 7284 36492 7290
rect 36360 7278 36492 7284
rect 36372 7262 36492 7278
rect 35348 6656 35400 6662
rect 35348 6598 35400 6604
rect 36268 6656 36320 6662
rect 36268 6598 36320 6604
rect 35360 6390 35388 6598
rect 35594 6556 35902 6565
rect 35594 6554 35600 6556
rect 35656 6554 35680 6556
rect 35736 6554 35760 6556
rect 35816 6554 35840 6556
rect 35896 6554 35902 6556
rect 35656 6502 35658 6554
rect 35838 6502 35840 6554
rect 35594 6500 35600 6502
rect 35656 6500 35680 6502
rect 35736 6500 35760 6502
rect 35816 6500 35840 6502
rect 35896 6500 35902 6502
rect 35594 6491 35902 6500
rect 36372 6458 36400 7262
rect 36556 7002 36584 7346
rect 36544 6996 36596 7002
rect 36544 6938 36596 6944
rect 36648 6730 36676 7482
rect 36728 7404 36780 7410
rect 36728 7346 36780 7352
rect 36740 7002 36768 7346
rect 36728 6996 36780 7002
rect 36728 6938 36780 6944
rect 36924 6798 36952 8366
rect 37016 7954 37044 9998
rect 37108 9926 37136 10016
rect 37188 9998 37240 10004
rect 37280 9988 37332 9994
rect 37280 9930 37332 9936
rect 37096 9920 37148 9926
rect 37096 9862 37148 9868
rect 37108 9586 37136 9862
rect 37292 9586 37320 9930
rect 37096 9580 37148 9586
rect 37096 9522 37148 9528
rect 37280 9580 37332 9586
rect 37280 9522 37332 9528
rect 37096 8968 37148 8974
rect 37096 8910 37148 8916
rect 37004 7948 37056 7954
rect 37004 7890 37056 7896
rect 37004 7404 37056 7410
rect 37004 7346 37056 7352
rect 37016 7274 37044 7346
rect 37004 7268 37056 7274
rect 37004 7210 37056 7216
rect 36912 6792 36964 6798
rect 36912 6734 36964 6740
rect 36636 6724 36688 6730
rect 36636 6666 36688 6672
rect 36360 6452 36412 6458
rect 36360 6394 36412 6400
rect 34796 6384 34848 6390
rect 34796 6326 34848 6332
rect 35348 6384 35400 6390
rect 35348 6326 35400 6332
rect 36176 6316 36228 6322
rect 36176 6258 36228 6264
rect 36268 6316 36320 6322
rect 36268 6258 36320 6264
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 36188 5914 36216 6258
rect 36176 5908 36228 5914
rect 36176 5850 36228 5856
rect 36188 5574 36216 5850
rect 36280 5710 36308 6258
rect 36636 6248 36688 6254
rect 36636 6190 36688 6196
rect 36648 5914 36676 6190
rect 37004 6112 37056 6118
rect 37004 6054 37056 6060
rect 36636 5908 36688 5914
rect 36636 5850 36688 5856
rect 36268 5704 36320 5710
rect 36268 5646 36320 5652
rect 34704 5568 34756 5574
rect 34704 5510 34756 5516
rect 36176 5568 36228 5574
rect 36176 5510 36228 5516
rect 34716 5370 34744 5510
rect 35594 5468 35902 5477
rect 35594 5466 35600 5468
rect 35656 5466 35680 5468
rect 35736 5466 35760 5468
rect 35816 5466 35840 5468
rect 35896 5466 35902 5468
rect 35656 5414 35658 5466
rect 35838 5414 35840 5466
rect 35594 5412 35600 5414
rect 35656 5412 35680 5414
rect 35736 5412 35760 5414
rect 35816 5412 35840 5414
rect 35896 5412 35902 5414
rect 35594 5403 35902 5412
rect 34704 5364 34756 5370
rect 34704 5306 34756 5312
rect 34796 5024 34848 5030
rect 34796 4966 34848 4972
rect 34808 4826 34836 4966
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 36188 4826 36216 5510
rect 36280 5370 36308 5646
rect 36268 5364 36320 5370
rect 36268 5306 36320 5312
rect 37016 5302 37044 6054
rect 37004 5296 37056 5302
rect 37004 5238 37056 5244
rect 37108 5234 37136 8910
rect 37292 8634 37320 9522
rect 37280 8628 37332 8634
rect 37280 8570 37332 8576
rect 37384 8498 37412 10662
rect 37476 10470 37504 11183
rect 37844 10470 37872 11222
rect 38304 11206 38424 11234
rect 38292 11144 38344 11150
rect 38198 11112 38254 11121
rect 38108 11076 38160 11082
rect 38292 11086 38344 11092
rect 38198 11047 38254 11056
rect 38108 11018 38160 11024
rect 37464 10464 37516 10470
rect 37464 10406 37516 10412
rect 37556 10464 37608 10470
rect 37556 10406 37608 10412
rect 37832 10464 37884 10470
rect 37832 10406 37884 10412
rect 37568 9994 37596 10406
rect 38120 10266 38148 11018
rect 38212 10742 38240 11047
rect 38200 10736 38252 10742
rect 38200 10678 38252 10684
rect 38304 10606 38332 11086
rect 38396 10742 38424 11206
rect 38384 10736 38436 10742
rect 38384 10678 38436 10684
rect 38488 10674 38516 11698
rect 38672 11354 38700 12038
rect 38750 11792 38806 11801
rect 38750 11727 38752 11736
rect 38804 11727 38806 11736
rect 38752 11698 38804 11704
rect 38660 11348 38712 11354
rect 38660 11290 38712 11296
rect 38856 11257 38884 12038
rect 38948 11762 38976 12679
rect 39212 12232 39264 12238
rect 39212 12174 39264 12180
rect 38936 11756 38988 11762
rect 38936 11698 38988 11704
rect 39028 11688 39080 11694
rect 39028 11630 39080 11636
rect 39120 11688 39172 11694
rect 39120 11630 39172 11636
rect 39040 11558 39068 11630
rect 39028 11552 39080 11558
rect 39028 11494 39080 11500
rect 39132 11354 39160 11630
rect 39224 11558 39252 12174
rect 39212 11552 39264 11558
rect 39212 11494 39264 11500
rect 39120 11348 39172 11354
rect 39120 11290 39172 11296
rect 39212 11348 39264 11354
rect 39212 11290 39264 11296
rect 39224 11257 39252 11290
rect 38842 11248 38898 11257
rect 38842 11183 38898 11192
rect 39210 11248 39266 11257
rect 39210 11183 39266 11192
rect 38568 11144 38620 11150
rect 38568 11086 38620 11092
rect 39212 11144 39264 11150
rect 39212 11086 39264 11092
rect 38476 10668 38528 10674
rect 38476 10610 38528 10616
rect 38292 10600 38344 10606
rect 38292 10542 38344 10548
rect 38580 10266 38608 11086
rect 39224 11014 39252 11086
rect 39212 11008 39264 11014
rect 39212 10950 39264 10956
rect 39316 10674 39344 12702
rect 39592 12434 39620 12786
rect 39776 12714 39804 13262
rect 39948 12776 40000 12782
rect 39948 12718 40000 12724
rect 39764 12708 39816 12714
rect 39764 12650 39816 12656
rect 39500 12406 39620 12434
rect 39672 12436 39724 12442
rect 39500 12238 39528 12406
rect 39672 12378 39724 12384
rect 39488 12232 39540 12238
rect 39488 12174 39540 12180
rect 39396 12096 39448 12102
rect 39396 12038 39448 12044
rect 39408 11898 39436 12038
rect 39396 11892 39448 11898
rect 39396 11834 39448 11840
rect 39500 11014 39528 12174
rect 39684 12170 39712 12378
rect 39960 12238 39988 12718
rect 39948 12232 40000 12238
rect 39948 12174 40000 12180
rect 39672 12164 39724 12170
rect 39672 12106 39724 12112
rect 39684 11694 39712 12106
rect 40052 11830 40080 13398
rect 40144 13394 40172 14214
rect 40420 13870 40448 14418
rect 40512 14006 40540 15370
rect 40500 14000 40552 14006
rect 40500 13942 40552 13948
rect 40604 13870 40632 17070
rect 40696 16726 40724 17274
rect 40788 16726 40816 19638
rect 40960 19372 41012 19378
rect 40960 19314 41012 19320
rect 40972 19174 41000 19314
rect 40960 19168 41012 19174
rect 40960 19110 41012 19116
rect 40868 18624 40920 18630
rect 40868 18566 40920 18572
rect 40880 18290 40908 18566
rect 40972 18426 41000 19110
rect 40960 18420 41012 18426
rect 40960 18362 41012 18368
rect 40868 18284 40920 18290
rect 40868 18226 40920 18232
rect 40960 18284 41012 18290
rect 40960 18226 41012 18232
rect 40880 17921 40908 18226
rect 40972 18193 41000 18226
rect 40958 18184 41014 18193
rect 40958 18119 41014 18128
rect 40960 18080 41012 18086
rect 40960 18022 41012 18028
rect 40866 17912 40922 17921
rect 40866 17847 40922 17856
rect 40866 17368 40922 17377
rect 40866 17303 40922 17312
rect 40880 17202 40908 17303
rect 40868 17196 40920 17202
rect 40868 17138 40920 17144
rect 40868 17060 40920 17066
rect 40868 17002 40920 17008
rect 40684 16720 40736 16726
rect 40684 16662 40736 16668
rect 40776 16720 40828 16726
rect 40776 16662 40828 16668
rect 40880 16658 40908 17002
rect 40972 16658 41000 18022
rect 41064 17202 41092 19722
rect 41616 19530 41644 21830
rect 41696 21344 41748 21350
rect 41696 21286 41748 21292
rect 41708 21010 41736 21286
rect 41696 21004 41748 21010
rect 41696 20946 41748 20952
rect 41696 19848 41748 19854
rect 41696 19790 41748 19796
rect 41432 19502 41644 19530
rect 41328 19440 41380 19446
rect 41328 19382 41380 19388
rect 41236 19304 41288 19310
rect 41236 19246 41288 19252
rect 41144 19236 41196 19242
rect 41144 19178 41196 19184
rect 41156 18057 41184 19178
rect 41248 18766 41276 19246
rect 41340 18902 41368 19382
rect 41328 18896 41380 18902
rect 41328 18838 41380 18844
rect 41236 18760 41288 18766
rect 41236 18702 41288 18708
rect 41142 18048 41198 18057
rect 41142 17983 41198 17992
rect 41248 17678 41276 18702
rect 41340 18086 41368 18838
rect 41328 18080 41380 18086
rect 41328 18022 41380 18028
rect 41236 17672 41288 17678
rect 41142 17640 41198 17649
rect 41236 17614 41288 17620
rect 41142 17575 41198 17584
rect 41156 17542 41184 17575
rect 41144 17536 41196 17542
rect 41144 17478 41196 17484
rect 41144 17264 41196 17270
rect 41144 17206 41196 17212
rect 41052 17196 41104 17202
rect 41052 17138 41104 17144
rect 41156 16726 41184 17206
rect 41052 16720 41104 16726
rect 41052 16662 41104 16668
rect 41144 16720 41196 16726
rect 41144 16662 41196 16668
rect 40868 16652 40920 16658
rect 40868 16594 40920 16600
rect 40960 16652 41012 16658
rect 40960 16594 41012 16600
rect 40776 16584 40828 16590
rect 40776 16526 40828 16532
rect 40880 16538 40908 16594
rect 41064 16538 41092 16662
rect 41142 16552 41198 16561
rect 40788 16266 40816 16526
rect 40880 16510 41000 16538
rect 41064 16510 41142 16538
rect 40696 16238 40816 16266
rect 40696 15706 40724 16238
rect 40868 16176 40920 16182
rect 40868 16118 40920 16124
rect 40972 16130 41000 16510
rect 41142 16487 41198 16496
rect 41156 16454 41184 16487
rect 41144 16448 41196 16454
rect 41144 16390 41196 16396
rect 41248 16250 41276 17614
rect 41328 17536 41380 17542
rect 41328 17478 41380 17484
rect 41340 16794 41368 17478
rect 41432 16946 41460 19502
rect 41602 18320 41658 18329
rect 41602 18255 41604 18264
rect 41656 18255 41658 18264
rect 41604 18226 41656 18232
rect 41512 18080 41564 18086
rect 41512 18022 41564 18028
rect 41524 17746 41552 18022
rect 41512 17740 41564 17746
rect 41512 17682 41564 17688
rect 41616 17066 41644 18226
rect 41604 17060 41656 17066
rect 41604 17002 41656 17008
rect 41432 16918 41644 16946
rect 41328 16788 41380 16794
rect 41328 16730 41380 16736
rect 41512 16720 41564 16726
rect 41510 16688 41512 16697
rect 41564 16688 41566 16697
rect 41328 16652 41380 16658
rect 41510 16623 41566 16632
rect 41328 16594 41380 16600
rect 41236 16244 41288 16250
rect 41236 16186 41288 16192
rect 40684 15700 40736 15706
rect 40684 15642 40736 15648
rect 40682 15600 40738 15609
rect 40682 15535 40738 15544
rect 40696 15366 40724 15535
rect 40880 15434 40908 16118
rect 40972 16102 41276 16130
rect 40958 15464 41014 15473
rect 40868 15428 40920 15434
rect 40958 15399 40960 15408
rect 40868 15370 40920 15376
rect 41012 15399 41014 15408
rect 40960 15370 41012 15376
rect 40684 15360 40736 15366
rect 40684 15302 40736 15308
rect 41248 15026 41276 16102
rect 41236 15020 41288 15026
rect 41236 14962 41288 14968
rect 41142 14920 41198 14929
rect 40960 14884 41012 14890
rect 41142 14855 41198 14864
rect 40960 14826 41012 14832
rect 40972 14414 41000 14826
rect 41156 14414 41184 14855
rect 41340 14618 41368 16594
rect 41524 15366 41552 16623
rect 41512 15360 41564 15366
rect 41512 15302 41564 15308
rect 41512 15088 41564 15094
rect 41432 15036 41512 15042
rect 41432 15030 41564 15036
rect 41432 15014 41552 15030
rect 41432 14958 41460 15014
rect 41420 14952 41472 14958
rect 41420 14894 41472 14900
rect 41512 14952 41564 14958
rect 41512 14894 41564 14900
rect 41328 14612 41380 14618
rect 41328 14554 41380 14560
rect 41328 14476 41380 14482
rect 41328 14418 41380 14424
rect 40960 14408 41012 14414
rect 40960 14350 41012 14356
rect 41144 14408 41196 14414
rect 41144 14350 41196 14356
rect 41340 14074 41368 14418
rect 40684 14068 40736 14074
rect 40684 14010 40736 14016
rect 41328 14068 41380 14074
rect 41328 14010 41380 14016
rect 40408 13864 40460 13870
rect 40408 13806 40460 13812
rect 40592 13864 40644 13870
rect 40592 13806 40644 13812
rect 40132 13388 40184 13394
rect 40132 13330 40184 13336
rect 40316 13252 40368 13258
rect 40316 13194 40368 13200
rect 40328 12238 40356 13194
rect 40604 12918 40632 13806
rect 40696 13394 40724 14010
rect 41524 14006 41552 14894
rect 41512 14000 41564 14006
rect 41512 13942 41564 13948
rect 41050 13560 41106 13569
rect 41524 13530 41552 13942
rect 41050 13495 41052 13504
rect 41104 13495 41106 13504
rect 41512 13524 41564 13530
rect 41052 13466 41104 13472
rect 41512 13466 41564 13472
rect 40684 13388 40736 13394
rect 40684 13330 40736 13336
rect 40592 12912 40644 12918
rect 40592 12854 40644 12860
rect 40316 12232 40368 12238
rect 40316 12174 40368 12180
rect 40592 12232 40644 12238
rect 40592 12174 40644 12180
rect 40040 11824 40092 11830
rect 40040 11766 40092 11772
rect 39856 11756 39908 11762
rect 39856 11698 39908 11704
rect 39948 11756 40000 11762
rect 39948 11698 40000 11704
rect 39672 11688 39724 11694
rect 39672 11630 39724 11636
rect 39868 11354 39896 11698
rect 39856 11348 39908 11354
rect 39856 11290 39908 11296
rect 39960 11257 39988 11698
rect 39946 11248 40002 11257
rect 40328 11218 40356 12174
rect 40604 11626 40632 12174
rect 40696 12102 40724 13330
rect 41064 13326 41092 13466
rect 41052 13320 41104 13326
rect 41052 13262 41104 13268
rect 40868 12436 40920 12442
rect 40868 12378 40920 12384
rect 40880 12238 40908 12378
rect 40868 12232 40920 12238
rect 40868 12174 40920 12180
rect 40960 12232 41012 12238
rect 40960 12174 41012 12180
rect 40776 12164 40828 12170
rect 40776 12106 40828 12112
rect 40684 12096 40736 12102
rect 40684 12038 40736 12044
rect 40788 11898 40816 12106
rect 40776 11892 40828 11898
rect 40776 11834 40828 11840
rect 40972 11830 41000 12174
rect 40960 11824 41012 11830
rect 40960 11766 41012 11772
rect 40592 11620 40644 11626
rect 40592 11562 40644 11568
rect 39946 11183 40002 11192
rect 40316 11212 40368 11218
rect 40316 11154 40368 11160
rect 39580 11076 39632 11082
rect 39580 11018 39632 11024
rect 39488 11008 39540 11014
rect 39488 10950 39540 10956
rect 39592 10810 39620 11018
rect 39580 10804 39632 10810
rect 39580 10746 39632 10752
rect 39304 10668 39356 10674
rect 39304 10610 39356 10616
rect 40592 10668 40644 10674
rect 40592 10610 40644 10616
rect 38108 10260 38160 10266
rect 38108 10202 38160 10208
rect 38568 10260 38620 10266
rect 38568 10202 38620 10208
rect 40604 10130 40632 10610
rect 39212 10124 39264 10130
rect 39212 10066 39264 10072
rect 40132 10124 40184 10130
rect 40132 10066 40184 10072
rect 40592 10124 40644 10130
rect 40592 10066 40644 10072
rect 37556 9988 37608 9994
rect 37556 9930 37608 9936
rect 39224 9654 39252 10066
rect 40040 10056 40092 10062
rect 40040 9998 40092 10004
rect 39212 9648 39264 9654
rect 39212 9590 39264 9596
rect 39396 9376 39448 9382
rect 39396 9318 39448 9324
rect 38016 9172 38068 9178
rect 38016 9114 38068 9120
rect 38028 8906 38056 9114
rect 39408 8906 39436 9318
rect 40052 9042 40080 9998
rect 40144 9722 40172 10066
rect 40132 9716 40184 9722
rect 40132 9658 40184 9664
rect 40040 9036 40092 9042
rect 40040 8978 40092 8984
rect 38016 8900 38068 8906
rect 38016 8842 38068 8848
rect 39396 8900 39448 8906
rect 39396 8842 39448 8848
rect 37832 8628 37884 8634
rect 37832 8570 37884 8576
rect 37372 8492 37424 8498
rect 37372 8434 37424 8440
rect 37188 7744 37240 7750
rect 37188 7686 37240 7692
rect 37200 7478 37228 7686
rect 37188 7472 37240 7478
rect 37188 7414 37240 7420
rect 37384 5914 37412 8434
rect 37556 8288 37608 8294
rect 37556 8230 37608 8236
rect 37568 7886 37596 8230
rect 37844 8090 37872 8570
rect 38028 8566 38056 8842
rect 40052 8566 40080 8978
rect 38016 8560 38068 8566
rect 37936 8508 38016 8514
rect 37936 8502 38068 8508
rect 40040 8560 40092 8566
rect 40040 8502 40092 8508
rect 37936 8486 38056 8502
rect 37832 8084 37884 8090
rect 37832 8026 37884 8032
rect 37556 7880 37608 7886
rect 37556 7822 37608 7828
rect 37648 7880 37700 7886
rect 37648 7822 37700 7828
rect 37660 7342 37688 7822
rect 37936 7478 37964 8486
rect 40052 7886 40080 8502
rect 40316 8424 40368 8430
rect 40316 8366 40368 8372
rect 40328 8090 40356 8366
rect 41064 8090 41092 13262
rect 41512 13252 41564 13258
rect 41512 13194 41564 13200
rect 41328 12300 41380 12306
rect 41328 12242 41380 12248
rect 41340 11762 41368 12242
rect 41328 11756 41380 11762
rect 41328 11698 41380 11704
rect 41236 10124 41288 10130
rect 41236 10066 41288 10072
rect 41248 9586 41276 10066
rect 41524 9994 41552 13194
rect 41616 12345 41644 16918
rect 41602 12336 41658 12345
rect 41602 12271 41658 12280
rect 41708 11082 41736 19790
rect 41800 17066 41828 22066
rect 41984 22066 42104 22094
rect 41880 21548 41932 21554
rect 41880 21490 41932 21496
rect 41892 21010 41920 21490
rect 41880 21004 41932 21010
rect 41880 20946 41932 20952
rect 41880 20324 41932 20330
rect 41880 20266 41932 20272
rect 41892 19854 41920 20266
rect 41880 19848 41932 19854
rect 41880 19790 41932 19796
rect 41984 17338 42012 22066
rect 42168 21593 42196 22374
rect 42260 22166 42288 22578
rect 42524 22568 42576 22574
rect 42524 22510 42576 22516
rect 42248 22160 42300 22166
rect 42248 22102 42300 22108
rect 42154 21584 42210 21593
rect 42154 21519 42210 21528
rect 42168 21418 42196 21519
rect 42156 21412 42208 21418
rect 42156 21354 42208 21360
rect 42432 20256 42484 20262
rect 42432 20198 42484 20204
rect 42064 19984 42116 19990
rect 42064 19926 42116 19932
rect 41972 17332 42024 17338
rect 41972 17274 42024 17280
rect 41788 17060 41840 17066
rect 41788 17002 41840 17008
rect 41788 16584 41840 16590
rect 41788 16526 41840 16532
rect 41800 15910 41828 16526
rect 41880 16516 41932 16522
rect 41984 16504 42012 17274
rect 41932 16476 42012 16504
rect 41880 16458 41932 16464
rect 42076 16454 42104 19926
rect 42444 19786 42472 20198
rect 42432 19780 42484 19786
rect 42432 19722 42484 19728
rect 42156 19372 42208 19378
rect 42156 19314 42208 19320
rect 42064 16448 42116 16454
rect 42064 16390 42116 16396
rect 41788 15904 41840 15910
rect 41788 15846 41840 15852
rect 41800 15502 41828 15846
rect 41788 15496 41840 15502
rect 41788 15438 41840 15444
rect 42168 15162 42196 19314
rect 42340 17196 42392 17202
rect 42340 17138 42392 17144
rect 42064 15156 42116 15162
rect 42064 15098 42116 15104
rect 42156 15156 42208 15162
rect 42156 15098 42208 15104
rect 42076 14657 42104 15098
rect 42168 14890 42196 15098
rect 42352 14890 42380 17138
rect 42536 16640 42564 22510
rect 42628 20602 42656 22578
rect 42720 21962 42748 22714
rect 42984 22636 43036 22642
rect 42984 22578 43036 22584
rect 42996 22438 43024 22578
rect 42984 22432 43036 22438
rect 42984 22374 43036 22380
rect 42708 21956 42760 21962
rect 42708 21898 42760 21904
rect 42720 20874 42748 21898
rect 42892 21684 42944 21690
rect 42892 21626 42944 21632
rect 42904 21146 42932 21626
rect 42984 21548 43036 21554
rect 42984 21490 43036 21496
rect 42892 21140 42944 21146
rect 42892 21082 42944 21088
rect 42904 20942 42932 21082
rect 42892 20936 42944 20942
rect 42892 20878 42944 20884
rect 42708 20868 42760 20874
rect 42708 20810 42760 20816
rect 42720 20602 42748 20810
rect 42996 20806 43024 21490
rect 43076 21480 43128 21486
rect 43076 21422 43128 21428
rect 42984 20800 43036 20806
rect 42984 20742 43036 20748
rect 42996 20641 43024 20742
rect 42982 20632 43038 20641
rect 42616 20596 42668 20602
rect 42616 20538 42668 20544
rect 42708 20596 42760 20602
rect 43088 20602 43116 21422
rect 42982 20567 43038 20576
rect 43076 20596 43128 20602
rect 42708 20538 42760 20544
rect 42628 20466 42656 20538
rect 42616 20460 42668 20466
rect 42616 20402 42668 20408
rect 42720 19786 42748 20538
rect 42800 20528 42852 20534
rect 42800 20470 42852 20476
rect 42890 20496 42946 20505
rect 42812 20262 42840 20470
rect 42996 20466 43024 20567
rect 43076 20538 43128 20544
rect 43168 20596 43220 20602
rect 43168 20538 43220 20544
rect 42890 20431 42892 20440
rect 42944 20431 42946 20440
rect 42984 20460 43036 20466
rect 42892 20402 42944 20408
rect 42984 20402 43036 20408
rect 42800 20256 42852 20262
rect 42800 20198 42852 20204
rect 42708 19780 42760 19786
rect 42708 19722 42760 19728
rect 42904 19378 42932 20402
rect 43180 20330 43208 20538
rect 43168 20324 43220 20330
rect 43168 20266 43220 20272
rect 42892 19372 42944 19378
rect 42892 19314 42944 19320
rect 43364 18426 43392 24511
rect 43442 24304 43498 24313
rect 43442 24239 43498 24248
rect 43456 24041 43484 24239
rect 43442 24032 43498 24041
rect 43442 23967 43498 23976
rect 43444 23316 43496 23322
rect 43444 23258 43496 23264
rect 43456 23118 43484 23258
rect 43444 23112 43496 23118
rect 43444 23054 43496 23060
rect 43536 22704 43588 22710
rect 43536 22646 43588 22652
rect 43548 22234 43576 22646
rect 43640 22409 43668 24534
rect 43732 24206 43760 24550
rect 43720 24200 43772 24206
rect 43720 24142 43772 24148
rect 43812 23588 43864 23594
rect 43812 23530 43864 23536
rect 43626 22400 43682 22409
rect 43626 22335 43682 22344
rect 43536 22228 43588 22234
rect 43536 22170 43588 22176
rect 43548 20466 43576 22170
rect 43824 22001 43852 23530
rect 44192 23322 44220 25842
rect 44272 25696 44324 25702
rect 44272 25638 44324 25644
rect 44456 25696 44508 25702
rect 44456 25638 44508 25644
rect 44180 23316 44232 23322
rect 44180 23258 44232 23264
rect 43904 22976 43956 22982
rect 43904 22918 43956 22924
rect 43810 21992 43866 22001
rect 43810 21927 43866 21936
rect 43536 20460 43588 20466
rect 43536 20402 43588 20408
rect 43548 20262 43576 20402
rect 43536 20256 43588 20262
rect 43536 20198 43588 20204
rect 43548 19334 43576 20198
rect 43720 19372 43772 19378
rect 43548 19306 43668 19334
rect 43720 19314 43772 19320
rect 43352 18420 43404 18426
rect 43352 18362 43404 18368
rect 42984 18216 43036 18222
rect 42984 18158 43036 18164
rect 42706 17912 42762 17921
rect 42706 17847 42762 17856
rect 42616 17808 42668 17814
rect 42616 17750 42668 17756
rect 42628 17270 42656 17750
rect 42720 17270 42748 17847
rect 42996 17746 43024 18158
rect 42984 17740 43036 17746
rect 42984 17682 43036 17688
rect 43364 17678 43392 18362
rect 43076 17672 43128 17678
rect 43076 17614 43128 17620
rect 43352 17672 43404 17678
rect 43352 17614 43404 17620
rect 43444 17672 43496 17678
rect 43444 17614 43496 17620
rect 43088 17338 43116 17614
rect 43076 17332 43128 17338
rect 43076 17274 43128 17280
rect 42616 17264 42668 17270
rect 42616 17206 42668 17212
rect 42708 17264 42760 17270
rect 43456 17252 43484 17614
rect 43456 17224 43576 17252
rect 42708 17206 42760 17212
rect 42628 17066 42656 17206
rect 42984 17128 43036 17134
rect 42984 17070 43036 17076
rect 43444 17128 43496 17134
rect 43444 17070 43496 17076
rect 42616 17060 42668 17066
rect 42616 17002 42668 17008
rect 42444 16612 42564 16640
rect 42156 14884 42208 14890
rect 42156 14826 42208 14832
rect 42340 14884 42392 14890
rect 42340 14826 42392 14832
rect 42444 14822 42472 16612
rect 42996 16590 43024 17070
rect 43166 16824 43222 16833
rect 43166 16759 43222 16768
rect 43180 16590 43208 16759
rect 42800 16584 42852 16590
rect 42800 16526 42852 16532
rect 42984 16584 43036 16590
rect 42984 16526 43036 16532
rect 43076 16584 43128 16590
rect 43076 16526 43128 16532
rect 43168 16584 43220 16590
rect 43168 16526 43220 16532
rect 42616 16448 42668 16454
rect 42616 16390 42668 16396
rect 42628 15638 42656 16390
rect 42812 16182 42840 16526
rect 42800 16176 42852 16182
rect 42800 16118 42852 16124
rect 43088 15706 43116 16526
rect 43180 16028 43208 16526
rect 43260 16040 43312 16046
rect 43180 16000 43260 16028
rect 43260 15982 43312 15988
rect 43456 15910 43484 17070
rect 43548 16998 43576 17224
rect 43536 16992 43588 16998
rect 43536 16934 43588 16940
rect 43444 15904 43496 15910
rect 43444 15846 43496 15852
rect 43076 15700 43128 15706
rect 43076 15642 43128 15648
rect 42616 15632 42668 15638
rect 42616 15574 42668 15580
rect 43456 15570 43484 15846
rect 43444 15564 43496 15570
rect 43444 15506 43496 15512
rect 43548 15502 43576 16934
rect 43640 15910 43668 19306
rect 43628 15904 43680 15910
rect 43628 15846 43680 15852
rect 43640 15502 43668 15846
rect 43352 15496 43404 15502
rect 43352 15438 43404 15444
rect 43536 15496 43588 15502
rect 43536 15438 43588 15444
rect 43628 15496 43680 15502
rect 43628 15438 43680 15444
rect 42524 15428 42576 15434
rect 42524 15370 42576 15376
rect 42432 14816 42484 14822
rect 42432 14758 42484 14764
rect 42062 14648 42118 14657
rect 42536 14618 42564 15370
rect 43076 15156 43128 15162
rect 43128 15116 43300 15144
rect 43076 15098 43128 15104
rect 42616 15020 42668 15026
rect 42616 14962 42668 14968
rect 42800 15020 42852 15026
rect 42800 14962 42852 14968
rect 42062 14583 42118 14592
rect 42524 14612 42576 14618
rect 42524 14554 42576 14560
rect 42432 14408 42484 14414
rect 42352 14368 42432 14396
rect 42064 14272 42116 14278
rect 42064 14214 42116 14220
rect 42076 14006 42104 14214
rect 42064 14000 42116 14006
rect 42064 13942 42116 13948
rect 42352 13870 42380 14368
rect 42432 14350 42484 14356
rect 42628 14278 42656 14962
rect 42708 14816 42760 14822
rect 42708 14758 42760 14764
rect 42616 14272 42668 14278
rect 42616 14214 42668 14220
rect 42720 14006 42748 14758
rect 42812 14618 42840 14962
rect 43272 14890 43300 15116
rect 43260 14884 43312 14890
rect 43260 14826 43312 14832
rect 43076 14816 43128 14822
rect 43076 14758 43128 14764
rect 42800 14612 42852 14618
rect 42800 14554 42852 14560
rect 43088 14482 43116 14758
rect 43076 14476 43128 14482
rect 43076 14418 43128 14424
rect 42708 14000 42760 14006
rect 42708 13942 42760 13948
rect 43088 13870 43116 14418
rect 43364 14414 43392 15438
rect 43444 14952 43496 14958
rect 43444 14894 43496 14900
rect 43352 14408 43404 14414
rect 43352 14350 43404 14356
rect 43456 14006 43484 14894
rect 43444 14000 43496 14006
rect 43444 13942 43496 13948
rect 42340 13864 42392 13870
rect 42340 13806 42392 13812
rect 43076 13864 43128 13870
rect 43076 13806 43128 13812
rect 42432 13524 42484 13530
rect 42432 13466 42484 13472
rect 42444 12170 42472 13466
rect 42892 12776 42944 12782
rect 42892 12718 42944 12724
rect 42800 12640 42852 12646
rect 42800 12582 42852 12588
rect 42432 12164 42484 12170
rect 42432 12106 42484 12112
rect 42444 11898 42472 12106
rect 42432 11892 42484 11898
rect 42432 11834 42484 11840
rect 42812 11830 42840 12582
rect 42904 12209 42932 12718
rect 43732 12442 43760 19314
rect 43824 17882 43852 21927
rect 43916 21894 43944 22918
rect 43996 22568 44048 22574
rect 44048 22516 44220 22522
rect 43996 22510 44220 22516
rect 44008 22494 44220 22510
rect 44086 22400 44142 22409
rect 44086 22335 44142 22344
rect 43904 21888 43956 21894
rect 43904 21830 43956 21836
rect 43812 17876 43864 17882
rect 43812 17818 43864 17824
rect 43824 17678 43852 17818
rect 43812 17672 43864 17678
rect 43812 17614 43864 17620
rect 43916 17338 43944 21830
rect 43996 21684 44048 21690
rect 43996 21626 44048 21632
rect 44008 21078 44036 21626
rect 44100 21146 44128 22335
rect 44192 22098 44220 22494
rect 44180 22092 44232 22098
rect 44180 22034 44232 22040
rect 44192 21486 44220 22034
rect 44180 21480 44232 21486
rect 44180 21422 44232 21428
rect 44088 21140 44140 21146
rect 44088 21082 44140 21088
rect 43996 21072 44048 21078
rect 43996 21014 44048 21020
rect 44192 19922 44220 21422
rect 44284 21078 44312 25638
rect 44468 25430 44496 25638
rect 44456 25424 44508 25430
rect 44456 25366 44508 25372
rect 44824 24064 44876 24070
rect 44824 24006 44876 24012
rect 44836 23798 44864 24006
rect 44824 23792 44876 23798
rect 44824 23734 44876 23740
rect 45112 23526 45140 27270
rect 45560 26444 45612 26450
rect 45560 26386 45612 26392
rect 45572 25838 45600 26386
rect 45756 26042 45784 27900
rect 45928 27882 45980 27888
rect 46480 27872 46532 27878
rect 46480 27814 46532 27820
rect 46492 27674 46520 27814
rect 47412 27674 47440 29446
rect 49712 28150 49740 29582
rect 50620 28552 50672 28558
rect 50620 28494 50672 28500
rect 49884 28416 49936 28422
rect 49884 28358 49936 28364
rect 48136 28144 48188 28150
rect 48136 28086 48188 28092
rect 49700 28144 49752 28150
rect 49700 28086 49752 28092
rect 47584 28076 47636 28082
rect 47584 28018 47636 28024
rect 46480 27668 46532 27674
rect 46480 27610 46532 27616
rect 47400 27668 47452 27674
rect 47400 27610 47452 27616
rect 46296 27464 46348 27470
rect 46296 27406 46348 27412
rect 45836 26512 45888 26518
rect 45836 26454 45888 26460
rect 45744 26036 45796 26042
rect 45744 25978 45796 25984
rect 45560 25832 45612 25838
rect 45560 25774 45612 25780
rect 45572 25276 45600 25774
rect 45652 25288 45704 25294
rect 45572 25248 45652 25276
rect 45652 25230 45704 25236
rect 45664 24274 45692 25230
rect 45848 24954 45876 26454
rect 46308 26450 46336 27406
rect 47412 27402 47440 27610
rect 47400 27396 47452 27402
rect 47400 27338 47452 27344
rect 47596 27334 47624 28018
rect 48148 27674 48176 28086
rect 49608 28076 49660 28082
rect 49608 28018 49660 28024
rect 49424 27872 49476 27878
rect 49424 27814 49476 27820
rect 48136 27668 48188 27674
rect 48136 27610 48188 27616
rect 48228 27532 48280 27538
rect 48228 27474 48280 27480
rect 47584 27328 47636 27334
rect 47584 27270 47636 27276
rect 48240 26858 48268 27474
rect 49436 27062 49464 27814
rect 49424 27056 49476 27062
rect 49424 26998 49476 27004
rect 48320 26920 48372 26926
rect 48320 26862 48372 26868
rect 48688 26920 48740 26926
rect 48688 26862 48740 26868
rect 49148 26920 49200 26926
rect 49148 26862 49200 26868
rect 48228 26852 48280 26858
rect 48228 26794 48280 26800
rect 46848 26784 46900 26790
rect 46848 26726 46900 26732
rect 46860 26450 46888 26726
rect 46296 26444 46348 26450
rect 46296 26386 46348 26392
rect 46848 26444 46900 26450
rect 46848 26386 46900 26392
rect 48044 26444 48096 26450
rect 48044 26386 48096 26392
rect 47124 26308 47176 26314
rect 47124 26250 47176 26256
rect 45928 26240 45980 26246
rect 45928 26182 45980 26188
rect 45940 25974 45968 26182
rect 47136 26042 47164 26250
rect 47124 26036 47176 26042
rect 47124 25978 47176 25984
rect 45928 25968 45980 25974
rect 45928 25910 45980 25916
rect 47216 25968 47268 25974
rect 47216 25910 47268 25916
rect 46480 25356 46532 25362
rect 46480 25298 46532 25304
rect 45928 25220 45980 25226
rect 45928 25162 45980 25168
rect 45940 24954 45968 25162
rect 45836 24948 45888 24954
rect 45836 24890 45888 24896
rect 45928 24948 45980 24954
rect 45928 24890 45980 24896
rect 45652 24268 45704 24274
rect 45652 24210 45704 24216
rect 45284 24132 45336 24138
rect 45284 24074 45336 24080
rect 45296 23866 45324 24074
rect 45284 23860 45336 23866
rect 45284 23802 45336 23808
rect 45376 23792 45428 23798
rect 45296 23740 45376 23746
rect 45296 23734 45428 23740
rect 45192 23724 45244 23730
rect 45192 23666 45244 23672
rect 45296 23718 45416 23734
rect 44456 23520 44508 23526
rect 44456 23462 44508 23468
rect 45100 23520 45152 23526
rect 45100 23462 45152 23468
rect 44364 22976 44416 22982
rect 44364 22918 44416 22924
rect 44376 22710 44404 22918
rect 44364 22704 44416 22710
rect 44364 22646 44416 22652
rect 44468 22094 44496 23462
rect 45204 23118 45232 23666
rect 45192 23112 45244 23118
rect 45192 23054 45244 23060
rect 44376 22066 44496 22094
rect 44272 21072 44324 21078
rect 44272 21014 44324 21020
rect 44272 20936 44324 20942
rect 44272 20878 44324 20884
rect 44284 20602 44312 20878
rect 44376 20874 44404 22066
rect 45204 22030 45232 23054
rect 45296 23050 45324 23718
rect 45652 23588 45704 23594
rect 45652 23530 45704 23536
rect 45468 23316 45520 23322
rect 45468 23258 45520 23264
rect 45284 23044 45336 23050
rect 45284 22986 45336 22992
rect 45296 22166 45324 22986
rect 45284 22160 45336 22166
rect 45284 22102 45336 22108
rect 44456 22024 44508 22030
rect 44456 21966 44508 21972
rect 45192 22024 45244 22030
rect 45192 21966 45244 21972
rect 44468 21298 44496 21966
rect 44824 21956 44876 21962
rect 44824 21898 44876 21904
rect 44640 21684 44692 21690
rect 44640 21626 44692 21632
rect 44548 21344 44600 21350
rect 44468 21292 44548 21298
rect 44468 21286 44600 21292
rect 44468 21270 44588 21286
rect 44468 20942 44496 21270
rect 44652 20942 44680 21626
rect 44456 20936 44508 20942
rect 44456 20878 44508 20884
rect 44640 20936 44692 20942
rect 44640 20878 44692 20884
rect 44732 20936 44784 20942
rect 44732 20878 44784 20884
rect 44364 20868 44416 20874
rect 44364 20810 44416 20816
rect 44744 20806 44772 20878
rect 44732 20800 44784 20806
rect 44732 20742 44784 20748
rect 44272 20596 44324 20602
rect 44272 20538 44324 20544
rect 44836 20466 44864 21898
rect 45284 21888 45336 21894
rect 45284 21830 45336 21836
rect 45008 21480 45060 21486
rect 45008 21422 45060 21428
rect 45020 21146 45048 21422
rect 45008 21140 45060 21146
rect 45008 21082 45060 21088
rect 45296 20942 45324 21830
rect 45480 21593 45508 23258
rect 45664 23118 45692 23530
rect 45848 23322 45876 24890
rect 46492 24818 46520 25298
rect 47228 25226 47256 25910
rect 47952 25900 48004 25906
rect 48056 25888 48084 26386
rect 48136 26308 48188 26314
rect 48136 26250 48188 26256
rect 48148 25974 48176 26250
rect 48228 26240 48280 26246
rect 48228 26182 48280 26188
rect 48136 25968 48188 25974
rect 48136 25910 48188 25916
rect 48004 25860 48084 25888
rect 47952 25842 48004 25848
rect 47308 25832 47360 25838
rect 47308 25774 47360 25780
rect 47216 25220 47268 25226
rect 47216 25162 47268 25168
rect 46940 25152 46992 25158
rect 46940 25094 46992 25100
rect 46952 24857 46980 25094
rect 46938 24848 46994 24857
rect 46112 24812 46164 24818
rect 46112 24754 46164 24760
rect 46480 24812 46532 24818
rect 46938 24783 46994 24792
rect 46480 24754 46532 24760
rect 46124 23866 46152 24754
rect 46388 24608 46440 24614
rect 46388 24550 46440 24556
rect 47032 24608 47084 24614
rect 47032 24550 47084 24556
rect 47216 24608 47268 24614
rect 47216 24550 47268 24556
rect 46400 24138 46428 24550
rect 46848 24268 46900 24274
rect 46848 24210 46900 24216
rect 46388 24132 46440 24138
rect 46388 24074 46440 24080
rect 46112 23860 46164 23866
rect 46112 23802 46164 23808
rect 46400 23497 46428 24074
rect 46664 23792 46716 23798
rect 46664 23734 46716 23740
rect 46386 23488 46442 23497
rect 46386 23423 46442 23432
rect 45836 23316 45888 23322
rect 45836 23258 45888 23264
rect 46020 23248 46072 23254
rect 46020 23190 46072 23196
rect 45652 23112 45704 23118
rect 45652 23054 45704 23060
rect 45560 22976 45612 22982
rect 45560 22918 45612 22924
rect 45572 22234 45600 22918
rect 45560 22228 45612 22234
rect 45560 22170 45612 22176
rect 45560 21956 45612 21962
rect 45560 21898 45612 21904
rect 45572 21690 45600 21898
rect 45560 21684 45612 21690
rect 45560 21626 45612 21632
rect 45466 21584 45522 21593
rect 45466 21519 45522 21528
rect 45480 21146 45508 21519
rect 45468 21140 45520 21146
rect 45468 21082 45520 21088
rect 45284 20936 45336 20942
rect 45284 20878 45336 20884
rect 44916 20868 44968 20874
rect 44916 20810 44968 20816
rect 44928 20641 44956 20810
rect 44914 20632 44970 20641
rect 44914 20567 44970 20576
rect 45100 20596 45152 20602
rect 44928 20534 44956 20567
rect 45100 20538 45152 20544
rect 44916 20528 44968 20534
rect 44916 20470 44968 20476
rect 44364 20460 44416 20466
rect 44364 20402 44416 20408
rect 44824 20460 44876 20466
rect 44824 20402 44876 20408
rect 44180 19916 44232 19922
rect 44180 19858 44232 19864
rect 44376 19718 44404 20402
rect 44364 19712 44416 19718
rect 44364 19654 44416 19660
rect 44376 19310 44404 19654
rect 44364 19304 44416 19310
rect 44364 19246 44416 19252
rect 45008 18760 45060 18766
rect 45008 18702 45060 18708
rect 44088 18692 44140 18698
rect 44088 18634 44140 18640
rect 44100 17610 44128 18634
rect 45020 17746 45048 18702
rect 45008 17740 45060 17746
rect 45008 17682 45060 17688
rect 44088 17604 44140 17610
rect 44088 17546 44140 17552
rect 44100 17338 44128 17546
rect 43904 17332 43956 17338
rect 43904 17274 43956 17280
rect 44088 17332 44140 17338
rect 44088 17274 44140 17280
rect 44548 17332 44600 17338
rect 44548 17274 44600 17280
rect 43812 17128 43864 17134
rect 43812 17070 43864 17076
rect 43824 16454 43852 17070
rect 44100 16946 44128 17274
rect 44008 16918 44128 16946
rect 44008 16726 44036 16918
rect 43996 16720 44048 16726
rect 43996 16662 44048 16668
rect 43904 16584 43956 16590
rect 43904 16526 43956 16532
rect 43812 16448 43864 16454
rect 43812 16390 43864 16396
rect 43810 14648 43866 14657
rect 43810 14583 43812 14592
rect 43864 14583 43866 14592
rect 43812 14554 43864 14560
rect 43916 14278 43944 16526
rect 44008 16114 44036 16662
rect 44180 16584 44232 16590
rect 44180 16526 44232 16532
rect 44192 16250 44220 16526
rect 44180 16244 44232 16250
rect 44180 16186 44232 16192
rect 43996 16108 44048 16114
rect 43996 16050 44048 16056
rect 44560 16046 44588 17274
rect 44732 16108 44784 16114
rect 44652 16068 44732 16096
rect 44548 16040 44600 16046
rect 44468 16000 44548 16028
rect 44088 15496 44140 15502
rect 44088 15438 44140 15444
rect 43996 15428 44048 15434
rect 43996 15370 44048 15376
rect 44008 15162 44036 15370
rect 43996 15156 44048 15162
rect 43996 15098 44048 15104
rect 43904 14272 43956 14278
rect 43904 14214 43956 14220
rect 43916 13920 43944 14214
rect 44008 14056 44036 15098
rect 44100 14929 44128 15438
rect 44180 14952 44232 14958
rect 44086 14920 44142 14929
rect 44180 14894 44232 14900
rect 44272 14952 44324 14958
rect 44272 14894 44324 14900
rect 44086 14855 44142 14864
rect 44088 14816 44140 14822
rect 44088 14758 44140 14764
rect 44100 14482 44128 14758
rect 44088 14476 44140 14482
rect 44088 14418 44140 14424
rect 44192 14346 44220 14894
rect 44180 14340 44232 14346
rect 44180 14282 44232 14288
rect 44284 14074 44312 14894
rect 44468 14550 44496 16000
rect 44548 15982 44600 15988
rect 44548 15360 44600 15366
rect 44548 15302 44600 15308
rect 44456 14544 44508 14550
rect 44456 14486 44508 14492
rect 44088 14068 44140 14074
rect 44008 14028 44088 14056
rect 44088 14010 44140 14016
rect 44272 14068 44324 14074
rect 44272 14010 44324 14016
rect 44560 13938 44588 15302
rect 44652 14822 44680 16068
rect 44732 16050 44784 16056
rect 44916 15564 44968 15570
rect 44916 15506 44968 15512
rect 44928 15026 44956 15506
rect 44916 15020 44968 15026
rect 44916 14962 44968 14968
rect 44640 14816 44692 14822
rect 44640 14758 44692 14764
rect 44652 13938 44680 14758
rect 43996 13932 44048 13938
rect 43916 13892 43996 13920
rect 43996 13874 44048 13880
rect 44456 13932 44508 13938
rect 44456 13874 44508 13880
rect 44548 13932 44600 13938
rect 44548 13874 44600 13880
rect 44640 13932 44692 13938
rect 44640 13874 44692 13880
rect 44468 13326 44496 13874
rect 44928 13394 44956 14962
rect 45112 14822 45140 20538
rect 45664 20330 45692 23054
rect 45652 20324 45704 20330
rect 45652 20266 45704 20272
rect 45192 20256 45244 20262
rect 45192 20198 45244 20204
rect 45560 20256 45612 20262
rect 45560 20198 45612 20204
rect 45204 19854 45232 20198
rect 45192 19848 45244 19854
rect 45192 19790 45244 19796
rect 45376 19848 45428 19854
rect 45376 19790 45428 19796
rect 45468 19848 45520 19854
rect 45468 19790 45520 19796
rect 45284 19168 45336 19174
rect 45284 19110 45336 19116
rect 45296 18834 45324 19110
rect 45284 18828 45336 18834
rect 45284 18770 45336 18776
rect 45284 16992 45336 16998
rect 45284 16934 45336 16940
rect 45296 16590 45324 16934
rect 45388 16794 45416 19790
rect 45480 19514 45508 19790
rect 45572 19786 45600 20198
rect 45560 19780 45612 19786
rect 45560 19722 45612 19728
rect 45468 19508 45520 19514
rect 45468 19450 45520 19456
rect 45468 19304 45520 19310
rect 45468 19246 45520 19252
rect 45480 18426 45508 19246
rect 45572 18737 45600 19722
rect 45558 18728 45614 18737
rect 45558 18663 45614 18672
rect 45468 18420 45520 18426
rect 45468 18362 45520 18368
rect 46032 17202 46060 23190
rect 46296 23112 46348 23118
rect 46296 23054 46348 23060
rect 46308 22438 46336 23054
rect 46296 22432 46348 22438
rect 46296 22374 46348 22380
rect 46112 21344 46164 21350
rect 46112 21286 46164 21292
rect 46124 20942 46152 21286
rect 46112 20936 46164 20942
rect 46112 20878 46164 20884
rect 46296 20800 46348 20806
rect 46296 20742 46348 20748
rect 46308 17202 46336 20742
rect 46400 19922 46428 23423
rect 46676 23322 46704 23734
rect 46756 23724 46808 23730
rect 46756 23666 46808 23672
rect 46664 23316 46716 23322
rect 46664 23258 46716 23264
rect 46676 23050 46704 23258
rect 46664 23044 46716 23050
rect 46664 22986 46716 22992
rect 46676 22642 46704 22986
rect 46768 22982 46796 23666
rect 46756 22976 46808 22982
rect 46756 22918 46808 22924
rect 46664 22636 46716 22642
rect 46664 22578 46716 22584
rect 46860 22098 46888 24210
rect 46940 24132 46992 24138
rect 46940 24074 46992 24080
rect 46952 23730 46980 24074
rect 47044 23730 47072 24550
rect 47124 24064 47176 24070
rect 47124 24006 47176 24012
rect 46940 23724 46992 23730
rect 46940 23666 46992 23672
rect 47032 23724 47084 23730
rect 47032 23666 47084 23672
rect 47136 23526 47164 24006
rect 47228 23905 47256 24550
rect 47320 24138 47348 25774
rect 47964 25362 47992 25842
rect 48240 25498 48268 26182
rect 48332 26042 48360 26862
rect 48700 26586 48728 26862
rect 48688 26580 48740 26586
rect 48688 26522 48740 26528
rect 48700 26382 48728 26522
rect 48688 26376 48740 26382
rect 48688 26318 48740 26324
rect 49160 26314 49188 26862
rect 49620 26586 49648 28018
rect 49712 27470 49740 28086
rect 49896 28082 49924 28358
rect 49884 28076 49936 28082
rect 49884 28018 49936 28024
rect 50068 28076 50120 28082
rect 50068 28018 50120 28024
rect 50080 27878 50108 28018
rect 49792 27872 49844 27878
rect 49792 27814 49844 27820
rect 50068 27872 50120 27878
rect 50068 27814 50120 27820
rect 49804 27538 49832 27814
rect 49792 27532 49844 27538
rect 49792 27474 49844 27480
rect 49700 27464 49752 27470
rect 49700 27406 49752 27412
rect 49712 26790 49740 27406
rect 49884 27124 49936 27130
rect 49884 27066 49936 27072
rect 49700 26784 49752 26790
rect 49700 26726 49752 26732
rect 49608 26580 49660 26586
rect 49608 26522 49660 26528
rect 49516 26512 49568 26518
rect 49514 26480 49516 26489
rect 49568 26480 49570 26489
rect 49514 26415 49570 26424
rect 49528 26382 49556 26415
rect 49516 26376 49568 26382
rect 49516 26318 49568 26324
rect 48780 26308 48832 26314
rect 48780 26250 48832 26256
rect 49148 26308 49200 26314
rect 49148 26250 49200 26256
rect 49332 26308 49384 26314
rect 49332 26250 49384 26256
rect 49700 26308 49752 26314
rect 49700 26250 49752 26256
rect 49792 26308 49844 26314
rect 49792 26250 49844 26256
rect 48320 26036 48372 26042
rect 48320 25978 48372 25984
rect 48688 25900 48740 25906
rect 48608 25860 48688 25888
rect 48228 25492 48280 25498
rect 48228 25434 48280 25440
rect 47952 25356 48004 25362
rect 47952 25298 48004 25304
rect 47492 25220 47544 25226
rect 47492 25162 47544 25168
rect 47400 24948 47452 24954
rect 47400 24890 47452 24896
rect 47412 24410 47440 24890
rect 47400 24404 47452 24410
rect 47400 24346 47452 24352
rect 47308 24132 47360 24138
rect 47308 24074 47360 24080
rect 47214 23896 47270 23905
rect 47214 23831 47270 23840
rect 47124 23520 47176 23526
rect 47124 23462 47176 23468
rect 46848 22092 46900 22098
rect 46848 22034 46900 22040
rect 46480 21956 46532 21962
rect 46480 21898 46532 21904
rect 46388 19916 46440 19922
rect 46388 19858 46440 19864
rect 46388 19372 46440 19378
rect 46388 19314 46440 19320
rect 46492 19334 46520 21898
rect 46860 21554 46888 22034
rect 47136 22001 47164 23462
rect 47216 22976 47268 22982
rect 47216 22918 47268 22924
rect 47228 22574 47256 22918
rect 47216 22568 47268 22574
rect 47216 22510 47268 22516
rect 47216 22024 47268 22030
rect 47122 21992 47178 22001
rect 47216 21966 47268 21972
rect 47306 21992 47362 22001
rect 47122 21927 47178 21936
rect 46848 21548 46900 21554
rect 46848 21490 46900 21496
rect 46848 20936 46900 20942
rect 46846 20904 46848 20913
rect 46900 20904 46902 20913
rect 46846 20839 46902 20848
rect 47136 20602 47164 21927
rect 47228 21865 47256 21966
rect 47306 21927 47362 21936
rect 47320 21894 47348 21927
rect 47308 21888 47360 21894
rect 47214 21856 47270 21865
rect 47308 21830 47360 21836
rect 47214 21791 47270 21800
rect 47124 20596 47176 20602
rect 47124 20538 47176 20544
rect 46756 20528 46808 20534
rect 46756 20470 46808 20476
rect 46664 19848 46716 19854
rect 46664 19790 46716 19796
rect 46676 19718 46704 19790
rect 46664 19712 46716 19718
rect 46664 19654 46716 19660
rect 46676 19446 46704 19654
rect 46664 19440 46716 19446
rect 46664 19382 46716 19388
rect 46020 17196 46072 17202
rect 46020 17138 46072 17144
rect 46204 17196 46256 17202
rect 46204 17138 46256 17144
rect 46296 17196 46348 17202
rect 46296 17138 46348 17144
rect 45376 16788 45428 16794
rect 45376 16730 45428 16736
rect 45284 16584 45336 16590
rect 45284 16526 45336 16532
rect 45388 16046 45416 16730
rect 45376 16040 45428 16046
rect 45376 15982 45428 15988
rect 46110 16008 46166 16017
rect 45100 14816 45152 14822
rect 45100 14758 45152 14764
rect 45388 13530 45416 15982
rect 46110 15943 46166 15952
rect 45652 15904 45704 15910
rect 45652 15846 45704 15852
rect 45928 15904 45980 15910
rect 45928 15846 45980 15852
rect 45664 14346 45692 15846
rect 45940 15434 45968 15846
rect 45928 15428 45980 15434
rect 45928 15370 45980 15376
rect 46020 15088 46072 15094
rect 46020 15030 46072 15036
rect 46032 14482 46060 15030
rect 46020 14476 46072 14482
rect 46020 14418 46072 14424
rect 45652 14340 45704 14346
rect 45652 14282 45704 14288
rect 45664 13938 45692 14282
rect 46032 14278 46060 14418
rect 46020 14272 46072 14278
rect 46020 14214 46072 14220
rect 46032 14074 46060 14214
rect 46020 14068 46072 14074
rect 46020 14010 46072 14016
rect 45652 13932 45704 13938
rect 45652 13874 45704 13880
rect 45376 13524 45428 13530
rect 45376 13466 45428 13472
rect 44916 13388 44968 13394
rect 44916 13330 44968 13336
rect 44456 13320 44508 13326
rect 44456 13262 44508 13268
rect 44928 12850 44956 13330
rect 45928 13320 45980 13326
rect 45928 13262 45980 13268
rect 45468 13184 45520 13190
rect 45468 13126 45520 13132
rect 45480 12918 45508 13126
rect 45468 12912 45520 12918
rect 45468 12854 45520 12860
rect 44916 12844 44968 12850
rect 44916 12786 44968 12792
rect 44272 12776 44324 12782
rect 44272 12718 44324 12724
rect 43720 12436 43772 12442
rect 43720 12378 43772 12384
rect 42890 12200 42946 12209
rect 42890 12135 42946 12144
rect 44284 11898 44312 12718
rect 45940 12646 45968 13262
rect 46124 12866 46152 15943
rect 46216 14006 46244 17138
rect 46308 16658 46336 17138
rect 46296 16652 46348 16658
rect 46296 16594 46348 16600
rect 46400 15094 46428 19314
rect 46492 19306 46525 19334
rect 46497 19224 46525 19306
rect 46492 19196 46525 19224
rect 46662 19272 46718 19281
rect 46662 19207 46718 19216
rect 46492 17202 46520 19196
rect 46572 17264 46624 17270
rect 46572 17206 46624 17212
rect 46480 17196 46532 17202
rect 46480 17138 46532 17144
rect 46492 16794 46520 17138
rect 46480 16788 46532 16794
rect 46480 16730 46532 16736
rect 46584 16232 46612 17206
rect 46492 16204 46612 16232
rect 46388 15088 46440 15094
rect 46388 15030 46440 15036
rect 46296 14272 46348 14278
rect 46296 14214 46348 14220
rect 46204 14000 46256 14006
rect 46204 13942 46256 13948
rect 46308 13394 46336 14214
rect 46492 13938 46520 16204
rect 46572 16108 46624 16114
rect 46572 16050 46624 16056
rect 46584 15162 46612 16050
rect 46676 15366 46704 19207
rect 46768 18970 46796 20470
rect 47136 20398 47164 20538
rect 47124 20392 47176 20398
rect 47124 20334 47176 20340
rect 47032 20324 47084 20330
rect 47032 20266 47084 20272
rect 46848 19916 46900 19922
rect 46848 19858 46900 19864
rect 46860 19718 46888 19858
rect 46848 19712 46900 19718
rect 46848 19654 46900 19660
rect 46860 19242 46888 19654
rect 46940 19508 46992 19514
rect 46940 19450 46992 19456
rect 46952 19417 46980 19450
rect 46938 19408 46994 19417
rect 47044 19378 47072 20266
rect 46938 19343 46994 19352
rect 47032 19372 47084 19378
rect 47032 19314 47084 19320
rect 46848 19236 46900 19242
rect 46848 19178 46900 19184
rect 46756 18964 46808 18970
rect 46756 18906 46808 18912
rect 46768 18290 46796 18906
rect 46756 18284 46808 18290
rect 46756 18226 46808 18232
rect 46756 17604 46808 17610
rect 46756 17546 46808 17552
rect 46768 17338 46796 17546
rect 46756 17332 46808 17338
rect 46756 17274 46808 17280
rect 46860 16726 46888 19178
rect 47044 19174 47072 19314
rect 47124 19304 47176 19310
rect 47124 19246 47176 19252
rect 47032 19168 47084 19174
rect 47032 19110 47084 19116
rect 46848 16720 46900 16726
rect 46848 16662 46900 16668
rect 46860 16522 46888 16662
rect 46848 16516 46900 16522
rect 46848 16458 46900 16464
rect 46664 15360 46716 15366
rect 46664 15302 46716 15308
rect 46572 15156 46624 15162
rect 46572 15098 46624 15104
rect 46676 15026 46704 15302
rect 46664 15020 46716 15026
rect 46716 14980 46888 15008
rect 46664 14962 46716 14968
rect 46572 14408 46624 14414
rect 46572 14350 46624 14356
rect 46756 14408 46808 14414
rect 46756 14350 46808 14356
rect 46584 14074 46612 14350
rect 46664 14340 46716 14346
rect 46664 14282 46716 14288
rect 46572 14068 46624 14074
rect 46572 14010 46624 14016
rect 46676 14006 46704 14282
rect 46664 14000 46716 14006
rect 46664 13942 46716 13948
rect 46480 13932 46532 13938
rect 46480 13874 46532 13880
rect 46572 13932 46624 13938
rect 46572 13874 46624 13880
rect 46296 13388 46348 13394
rect 46296 13330 46348 13336
rect 46124 12838 46244 12866
rect 45928 12640 45980 12646
rect 45928 12582 45980 12588
rect 45940 12306 45968 12582
rect 46216 12442 46244 12838
rect 46584 12646 46612 13874
rect 46768 13870 46796 14350
rect 46756 13864 46808 13870
rect 46756 13806 46808 13812
rect 46860 13394 46888 14980
rect 47044 14618 47072 19110
rect 47136 18970 47164 19246
rect 47124 18964 47176 18970
rect 47124 18906 47176 18912
rect 47228 15201 47256 21791
rect 47320 20874 47348 21830
rect 47308 20868 47360 20874
rect 47308 20810 47360 20816
rect 47412 19242 47440 24346
rect 47504 23746 47532 25162
rect 47768 25152 47820 25158
rect 47768 25094 47820 25100
rect 47780 24138 47808 25094
rect 47584 24132 47636 24138
rect 47584 24074 47636 24080
rect 47768 24132 47820 24138
rect 47768 24074 47820 24080
rect 47596 23905 47624 24074
rect 47780 24018 47808 24074
rect 47688 23990 47808 24018
rect 47582 23896 47638 23905
rect 47582 23831 47638 23840
rect 47504 23718 47624 23746
rect 47688 23730 47716 23990
rect 47860 23860 47912 23866
rect 47860 23802 47912 23808
rect 47872 23730 47900 23802
rect 47964 23730 47992 25298
rect 48608 25226 48636 25860
rect 48688 25842 48740 25848
rect 48792 25786 48820 26250
rect 49056 26240 49108 26246
rect 49056 26182 49108 26188
rect 48700 25758 48820 25786
rect 48596 25220 48648 25226
rect 48516 25180 48596 25208
rect 48412 24268 48464 24274
rect 48412 24210 48464 24216
rect 48318 24168 48374 24177
rect 48318 24103 48374 24112
rect 48332 24070 48360 24103
rect 48136 24064 48188 24070
rect 48136 24006 48188 24012
rect 48320 24064 48372 24070
rect 48320 24006 48372 24012
rect 48042 23896 48098 23905
rect 48042 23831 48098 23840
rect 47492 23656 47544 23662
rect 47492 23598 47544 23604
rect 47504 23186 47532 23598
rect 47492 23180 47544 23186
rect 47492 23122 47544 23128
rect 47596 23050 47624 23718
rect 47676 23724 47728 23730
rect 47676 23666 47728 23672
rect 47768 23724 47820 23730
rect 47768 23666 47820 23672
rect 47860 23724 47912 23730
rect 47860 23666 47912 23672
rect 47952 23724 48004 23730
rect 47952 23666 48004 23672
rect 47780 23322 47808 23666
rect 47768 23316 47820 23322
rect 47768 23258 47820 23264
rect 47584 23044 47636 23050
rect 47584 22986 47636 22992
rect 47676 22568 47728 22574
rect 47676 22510 47728 22516
rect 47492 21480 47544 21486
rect 47492 21422 47544 21428
rect 47504 21146 47532 21422
rect 47492 21140 47544 21146
rect 47492 21082 47544 21088
rect 47584 21072 47636 21078
rect 47584 21014 47636 21020
rect 47492 20936 47544 20942
rect 47492 20878 47544 20884
rect 47504 20806 47532 20878
rect 47492 20800 47544 20806
rect 47492 20742 47544 20748
rect 47504 20346 47532 20742
rect 47596 20466 47624 21014
rect 47688 20942 47716 22510
rect 47860 22228 47912 22234
rect 47860 22170 47912 22176
rect 47872 21962 47900 22170
rect 47964 22030 47992 23666
rect 48056 22522 48084 23831
rect 48148 23662 48176 24006
rect 48136 23656 48188 23662
rect 48188 23604 48268 23610
rect 48136 23598 48268 23604
rect 48148 23582 48268 23598
rect 48136 23520 48188 23526
rect 48136 23462 48188 23468
rect 48148 22710 48176 23462
rect 48136 22704 48188 22710
rect 48136 22646 48188 22652
rect 48056 22494 48176 22522
rect 48044 22432 48096 22438
rect 48044 22374 48096 22380
rect 48056 22166 48084 22374
rect 48044 22160 48096 22166
rect 48044 22102 48096 22108
rect 47952 22024 48004 22030
rect 47952 21966 48004 21972
rect 47860 21956 47912 21962
rect 47860 21898 47912 21904
rect 47768 21888 47820 21894
rect 47768 21830 47820 21836
rect 47780 20942 47808 21830
rect 47952 21616 48004 21622
rect 47952 21558 48004 21564
rect 47964 21486 47992 21558
rect 47952 21480 48004 21486
rect 47952 21422 48004 21428
rect 47950 21176 48006 21185
rect 48056 21162 48084 22102
rect 48006 21134 48084 21162
rect 47950 21111 47952 21120
rect 48004 21111 48006 21120
rect 47952 21082 48004 21088
rect 47676 20936 47728 20942
rect 47676 20878 47728 20884
rect 47768 20936 47820 20942
rect 47768 20878 47820 20884
rect 47858 20632 47914 20641
rect 47858 20567 47860 20576
rect 47912 20567 47914 20576
rect 47964 20602 48084 20618
rect 47964 20596 48096 20602
rect 47964 20590 48044 20596
rect 47860 20538 47912 20544
rect 47872 20466 47900 20538
rect 47584 20460 47636 20466
rect 47584 20402 47636 20408
rect 47768 20460 47820 20466
rect 47768 20402 47820 20408
rect 47860 20460 47912 20466
rect 47860 20402 47912 20408
rect 47504 20318 47624 20346
rect 47492 19780 47544 19786
rect 47492 19722 47544 19728
rect 47400 19236 47452 19242
rect 47400 19178 47452 19184
rect 47412 18902 47440 19178
rect 47504 19174 47532 19722
rect 47492 19168 47544 19174
rect 47492 19110 47544 19116
rect 47400 18896 47452 18902
rect 47400 18838 47452 18844
rect 47504 17882 47532 19110
rect 47492 17876 47544 17882
rect 47492 17818 47544 17824
rect 47504 17082 47532 17818
rect 47596 17542 47624 20318
rect 47676 20324 47728 20330
rect 47676 20266 47728 20272
rect 47584 17536 47636 17542
rect 47584 17478 47636 17484
rect 47504 17054 47624 17082
rect 47492 16992 47544 16998
rect 47492 16934 47544 16940
rect 47504 16590 47532 16934
rect 47492 16584 47544 16590
rect 47492 16526 47544 16532
rect 47596 16522 47624 17054
rect 47584 16516 47636 16522
rect 47584 16458 47636 16464
rect 47596 16250 47624 16458
rect 47688 16250 47716 20266
rect 47780 20262 47808 20402
rect 47768 20256 47820 20262
rect 47768 20198 47820 20204
rect 47768 19848 47820 19854
rect 47768 19790 47820 19796
rect 47780 19242 47808 19790
rect 47964 19718 47992 20590
rect 48044 20538 48096 20544
rect 48148 20482 48176 22494
rect 48240 20602 48268 23582
rect 48320 23588 48372 23594
rect 48320 23530 48372 23536
rect 48332 22234 48360 23530
rect 48424 23186 48452 24210
rect 48516 23322 48544 25180
rect 48596 25162 48648 25168
rect 48700 25106 48728 25758
rect 48964 25288 49016 25294
rect 49068 25276 49096 26182
rect 49148 25832 49200 25838
rect 49148 25774 49200 25780
rect 49160 25294 49188 25774
rect 49344 25294 49372 26250
rect 49712 26042 49740 26250
rect 49700 26036 49752 26042
rect 49700 25978 49752 25984
rect 49516 25900 49568 25906
rect 49516 25842 49568 25848
rect 49016 25248 49096 25276
rect 48964 25230 49016 25236
rect 48608 25078 48728 25106
rect 48780 25152 48832 25158
rect 48780 25094 48832 25100
rect 48608 24154 48636 25078
rect 48792 24886 48820 25094
rect 48780 24880 48832 24886
rect 48964 24880 49016 24886
rect 48832 24840 48912 24868
rect 48780 24822 48832 24828
rect 48688 24404 48740 24410
rect 48688 24346 48740 24352
rect 48780 24404 48832 24410
rect 48780 24346 48832 24352
rect 48700 24274 48728 24346
rect 48688 24268 48740 24274
rect 48688 24210 48740 24216
rect 48608 24126 48728 24154
rect 48596 24064 48648 24070
rect 48596 24006 48648 24012
rect 48608 23730 48636 24006
rect 48596 23724 48648 23730
rect 48596 23666 48648 23672
rect 48504 23316 48556 23322
rect 48504 23258 48556 23264
rect 48412 23180 48464 23186
rect 48412 23122 48464 23128
rect 48320 22228 48372 22234
rect 48320 22170 48372 22176
rect 48320 22024 48372 22030
rect 48516 22012 48544 23258
rect 48372 21984 48544 22012
rect 48320 21966 48372 21972
rect 48332 21146 48360 21966
rect 48504 21888 48556 21894
rect 48504 21830 48556 21836
rect 48516 21593 48544 21830
rect 48502 21584 48558 21593
rect 48502 21519 48558 21528
rect 48608 21468 48636 23666
rect 48700 22438 48728 24126
rect 48792 23866 48820 24346
rect 48780 23860 48832 23866
rect 48780 23802 48832 23808
rect 48884 23168 48912 24840
rect 48964 24822 49016 24828
rect 48976 24614 49004 24822
rect 48964 24608 49016 24614
rect 48962 24576 48964 24585
rect 49016 24576 49018 24585
rect 48962 24511 49018 24520
rect 48964 24268 49016 24274
rect 48964 24210 49016 24216
rect 48976 23662 49004 24210
rect 48964 23656 49016 23662
rect 48964 23598 49016 23604
rect 48792 23140 48912 23168
rect 48688 22432 48740 22438
rect 48688 22374 48740 22380
rect 48688 22024 48740 22030
rect 48688 21966 48740 21972
rect 48700 21690 48728 21966
rect 48688 21684 48740 21690
rect 48688 21626 48740 21632
rect 48424 21440 48636 21468
rect 48320 21140 48372 21146
rect 48320 21082 48372 21088
rect 48424 21078 48452 21440
rect 48412 21072 48464 21078
rect 48412 21014 48464 21020
rect 48594 21040 48650 21049
rect 48228 20596 48280 20602
rect 48228 20538 48280 20544
rect 48056 20454 48176 20482
rect 48424 20482 48452 21014
rect 48594 20975 48650 20984
rect 48608 20942 48636 20975
rect 48700 20942 48728 21626
rect 48792 21468 48820 23140
rect 48976 23050 49004 23598
rect 49068 23508 49096 25248
rect 49148 25288 49200 25294
rect 49148 25230 49200 25236
rect 49332 25288 49384 25294
rect 49332 25230 49384 25236
rect 49424 25288 49476 25294
rect 49424 25230 49476 25236
rect 49436 24954 49464 25230
rect 49424 24948 49476 24954
rect 49424 24890 49476 24896
rect 49240 24744 49292 24750
rect 49238 24712 49240 24721
rect 49292 24712 49294 24721
rect 49294 24670 49372 24698
rect 49238 24647 49294 24656
rect 49146 24032 49202 24041
rect 49146 23967 49202 23976
rect 49160 23866 49188 23967
rect 49148 23860 49200 23866
rect 49148 23802 49200 23808
rect 49148 23520 49200 23526
rect 49068 23480 49148 23508
rect 49148 23462 49200 23468
rect 49240 23520 49292 23526
rect 49240 23462 49292 23468
rect 48872 23044 48924 23050
rect 48872 22986 48924 22992
rect 48964 23044 49016 23050
rect 48964 22986 49016 22992
rect 48884 22778 48912 22986
rect 48976 22953 49004 22986
rect 48962 22944 49018 22953
rect 48962 22879 49018 22888
rect 48872 22772 48924 22778
rect 48872 22714 48924 22720
rect 49056 22772 49108 22778
rect 49056 22714 49108 22720
rect 48872 22432 48924 22438
rect 48872 22374 48924 22380
rect 48884 21894 48912 22374
rect 49068 22030 49096 22714
rect 49056 22024 49108 22030
rect 49056 21966 49108 21972
rect 48872 21888 48924 21894
rect 48872 21830 48924 21836
rect 49056 21888 49108 21894
rect 49056 21830 49108 21836
rect 48884 21690 48912 21830
rect 48872 21684 48924 21690
rect 48872 21626 48924 21632
rect 49068 21593 49096 21830
rect 49054 21584 49110 21593
rect 49054 21519 49110 21528
rect 48872 21480 48924 21486
rect 48792 21440 48872 21468
rect 48792 20942 48820 21440
rect 48872 21422 48924 21428
rect 49056 21412 49108 21418
rect 49056 21354 49108 21360
rect 49068 21128 49096 21354
rect 48884 21100 49096 21128
rect 48884 21010 48912 21100
rect 48872 21004 48924 21010
rect 48872 20946 48924 20952
rect 49160 20942 49188 23462
rect 49252 23322 49280 23462
rect 49240 23316 49292 23322
rect 49240 23258 49292 23264
rect 49240 22636 49292 22642
rect 49240 22578 49292 22584
rect 49252 21593 49280 22578
rect 49344 22114 49372 24670
rect 49424 24608 49476 24614
rect 49424 24550 49476 24556
rect 49436 24206 49464 24550
rect 49528 24410 49556 25842
rect 49804 25838 49832 26250
rect 49792 25832 49844 25838
rect 49792 25774 49844 25780
rect 49608 25764 49660 25770
rect 49608 25706 49660 25712
rect 49620 25265 49648 25706
rect 49606 25256 49662 25265
rect 49606 25191 49662 25200
rect 49792 25152 49844 25158
rect 49792 25094 49844 25100
rect 49608 24676 49660 24682
rect 49608 24618 49660 24624
rect 49620 24426 49648 24618
rect 49620 24410 49740 24426
rect 49516 24404 49568 24410
rect 49620 24404 49752 24410
rect 49620 24398 49700 24404
rect 49516 24346 49568 24352
rect 49700 24346 49752 24352
rect 49424 24200 49476 24206
rect 49424 24142 49476 24148
rect 49700 23724 49752 23730
rect 49700 23666 49752 23672
rect 49712 23322 49740 23666
rect 49700 23316 49752 23322
rect 49700 23258 49752 23264
rect 49700 22772 49752 22778
rect 49700 22714 49752 22720
rect 49712 22234 49740 22714
rect 49700 22228 49752 22234
rect 49700 22170 49752 22176
rect 49344 22086 49648 22114
rect 49332 22024 49384 22030
rect 49332 21966 49384 21972
rect 49344 21729 49372 21966
rect 49330 21720 49386 21729
rect 49330 21655 49386 21664
rect 49332 21616 49384 21622
rect 49238 21584 49294 21593
rect 49332 21558 49384 21564
rect 49238 21519 49294 21528
rect 49252 21321 49280 21519
rect 49238 21312 49294 21321
rect 49238 21247 49294 21256
rect 49344 21146 49372 21558
rect 49424 21480 49476 21486
rect 49424 21422 49476 21428
rect 49332 21140 49384 21146
rect 49332 21082 49384 21088
rect 49238 21040 49294 21049
rect 49238 20975 49294 20984
rect 48596 20936 48648 20942
rect 48596 20878 48648 20884
rect 48688 20936 48740 20942
rect 48688 20878 48740 20884
rect 48780 20936 48832 20942
rect 48780 20878 48832 20884
rect 48964 20936 49016 20942
rect 48964 20878 49016 20884
rect 49056 20936 49108 20942
rect 49056 20878 49108 20884
rect 49148 20936 49200 20942
rect 49148 20878 49200 20884
rect 48792 20777 48820 20878
rect 48872 20800 48924 20806
rect 48778 20768 48834 20777
rect 48872 20742 48924 20748
rect 48778 20703 48834 20712
rect 48884 20602 48912 20742
rect 48872 20596 48924 20602
rect 48872 20538 48924 20544
rect 48594 20496 48650 20505
rect 48424 20454 48508 20482
rect 47952 19712 48004 19718
rect 47952 19654 48004 19660
rect 48056 19514 48084 20454
rect 48136 20392 48188 20398
rect 48480 20380 48508 20454
rect 48650 20466 48728 20482
rect 48650 20460 48740 20466
rect 48650 20454 48688 20460
rect 48594 20431 48650 20440
rect 48688 20402 48740 20408
rect 48780 20460 48832 20466
rect 48780 20402 48832 20408
rect 48480 20352 48544 20380
rect 48136 20334 48188 20340
rect 48148 19854 48176 20334
rect 48320 20324 48372 20330
rect 48320 20266 48372 20272
rect 48332 20058 48360 20266
rect 48320 20052 48372 20058
rect 48320 19994 48372 20000
rect 48228 19984 48280 19990
rect 48228 19926 48280 19932
rect 48136 19848 48188 19854
rect 48136 19790 48188 19796
rect 48240 19786 48268 19926
rect 48412 19848 48464 19854
rect 48412 19790 48464 19796
rect 48228 19780 48280 19786
rect 48228 19722 48280 19728
rect 48044 19508 48096 19514
rect 48044 19450 48096 19456
rect 47768 19236 47820 19242
rect 47768 19178 47820 19184
rect 47860 18692 47912 18698
rect 48240 18680 48268 19722
rect 48318 19544 48374 19553
rect 48318 19479 48374 19488
rect 48332 18850 48360 19479
rect 48424 18970 48452 19790
rect 48412 18964 48464 18970
rect 48412 18906 48464 18912
rect 48332 18822 48452 18850
rect 48320 18692 48372 18698
rect 48240 18652 48320 18680
rect 47860 18634 47912 18640
rect 48320 18634 48372 18640
rect 47872 17678 47900 18634
rect 48424 17921 48452 18822
rect 48410 17912 48466 17921
rect 48410 17847 48466 17856
rect 47952 17808 48004 17814
rect 47952 17750 48004 17756
rect 48226 17776 48282 17785
rect 47860 17672 47912 17678
rect 47860 17614 47912 17620
rect 47872 16794 47900 17614
rect 47860 16788 47912 16794
rect 47860 16730 47912 16736
rect 47768 16584 47820 16590
rect 47768 16526 47820 16532
rect 47584 16244 47636 16250
rect 47584 16186 47636 16192
rect 47676 16244 47728 16250
rect 47676 16186 47728 16192
rect 47400 16108 47452 16114
rect 47400 16050 47452 16056
rect 47308 15428 47360 15434
rect 47308 15370 47360 15376
rect 47214 15192 47270 15201
rect 47214 15127 47270 15136
rect 47216 15020 47268 15026
rect 47216 14962 47268 14968
rect 47228 14822 47256 14962
rect 47124 14816 47176 14822
rect 47124 14758 47176 14764
rect 47216 14816 47268 14822
rect 47216 14758 47268 14764
rect 47032 14612 47084 14618
rect 47032 14554 47084 14560
rect 47044 14346 47072 14554
rect 47032 14340 47084 14346
rect 47032 14282 47084 14288
rect 47136 13938 47164 14758
rect 47228 14346 47256 14758
rect 47216 14340 47268 14346
rect 47216 14282 47268 14288
rect 47124 13932 47176 13938
rect 47124 13874 47176 13880
rect 47228 13870 47256 14282
rect 47216 13864 47268 13870
rect 47216 13806 47268 13812
rect 46848 13388 46900 13394
rect 46848 13330 46900 13336
rect 47320 13258 47348 15370
rect 47412 15366 47440 16050
rect 47688 15706 47716 16186
rect 47780 16114 47808 16526
rect 47768 16108 47820 16114
rect 47768 16050 47820 16056
rect 47676 15700 47728 15706
rect 47676 15642 47728 15648
rect 47872 15434 47900 16730
rect 47964 16658 47992 17750
rect 48516 17762 48544 20352
rect 48596 20324 48648 20330
rect 48596 20266 48648 20272
rect 48608 19961 48636 20266
rect 48792 20233 48820 20402
rect 48872 20324 48924 20330
rect 48872 20266 48924 20272
rect 48778 20224 48834 20233
rect 48778 20159 48834 20168
rect 48686 20088 48742 20097
rect 48686 20023 48742 20032
rect 48594 19952 48650 19961
rect 48594 19887 48650 19896
rect 48594 19816 48650 19825
rect 48594 19751 48650 19760
rect 48608 17882 48636 19751
rect 48596 17876 48648 17882
rect 48596 17818 48648 17824
rect 48516 17734 48636 17762
rect 48226 17711 48282 17720
rect 48240 17542 48268 17711
rect 48412 17604 48464 17610
rect 48412 17546 48464 17552
rect 48228 17536 48280 17542
rect 48228 17478 48280 17484
rect 48320 17536 48372 17542
rect 48320 17478 48372 17484
rect 48332 17202 48360 17478
rect 48320 17196 48372 17202
rect 48320 17138 48372 17144
rect 48320 16992 48372 16998
rect 48240 16940 48320 16946
rect 48240 16934 48372 16940
rect 48240 16918 48360 16934
rect 48044 16788 48096 16794
rect 48044 16730 48096 16736
rect 48056 16658 48084 16730
rect 47952 16652 48004 16658
rect 47952 16594 48004 16600
rect 48044 16652 48096 16658
rect 48044 16594 48096 16600
rect 47964 15570 47992 16594
rect 48240 16561 48268 16918
rect 48320 16788 48372 16794
rect 48424 16776 48452 17546
rect 48504 17264 48556 17270
rect 48504 17206 48556 17212
rect 48516 17105 48544 17206
rect 48502 17096 48558 17105
rect 48502 17031 48558 17040
rect 48504 16992 48556 16998
rect 48504 16934 48556 16940
rect 48372 16748 48452 16776
rect 48320 16730 48372 16736
rect 48516 16726 48544 16934
rect 48504 16720 48556 16726
rect 48504 16662 48556 16668
rect 48226 16552 48282 16561
rect 48044 16516 48096 16522
rect 48226 16487 48282 16496
rect 48320 16516 48372 16522
rect 48044 16458 48096 16464
rect 48056 15978 48084 16458
rect 48240 16454 48268 16487
rect 48320 16458 48372 16464
rect 48228 16448 48280 16454
rect 48228 16390 48280 16396
rect 48228 16040 48280 16046
rect 48228 15982 48280 15988
rect 48044 15972 48096 15978
rect 48044 15914 48096 15920
rect 48044 15632 48096 15638
rect 48042 15600 48044 15609
rect 48096 15600 48098 15609
rect 47952 15564 48004 15570
rect 48042 15535 48098 15544
rect 47952 15506 48004 15512
rect 47860 15428 47912 15434
rect 47860 15370 47912 15376
rect 47400 15360 47452 15366
rect 47400 15302 47452 15308
rect 47412 14346 47440 15302
rect 47872 15094 47900 15370
rect 47860 15088 47912 15094
rect 47860 15030 47912 15036
rect 47964 15026 47992 15506
rect 47952 15020 48004 15026
rect 47952 14962 48004 14968
rect 48240 14906 48268 15982
rect 48148 14878 48268 14906
rect 47584 14408 47636 14414
rect 47584 14350 47636 14356
rect 47400 14340 47452 14346
rect 47400 14282 47452 14288
rect 47412 14006 47440 14282
rect 47596 14074 47624 14350
rect 47584 14068 47636 14074
rect 47584 14010 47636 14016
rect 47400 14000 47452 14006
rect 47400 13942 47452 13948
rect 48148 13326 48176 14878
rect 48228 14816 48280 14822
rect 48332 14770 48360 16458
rect 48412 16244 48464 16250
rect 48412 16186 48464 16192
rect 48424 15978 48452 16186
rect 48412 15972 48464 15978
rect 48412 15914 48464 15920
rect 48516 15065 48544 16662
rect 48608 16590 48636 17734
rect 48596 16584 48648 16590
rect 48596 16526 48648 16532
rect 48596 16448 48648 16454
rect 48700 16436 48728 20023
rect 48780 19712 48832 19718
rect 48780 19654 48832 19660
rect 48792 19378 48820 19654
rect 48780 19372 48832 19378
rect 48780 19314 48832 19320
rect 48884 19258 48912 20266
rect 48976 20097 49004 20878
rect 48962 20088 49018 20097
rect 49068 20058 49096 20878
rect 49160 20777 49188 20878
rect 49252 20806 49280 20975
rect 49332 20936 49384 20942
rect 49436 20924 49464 21422
rect 49516 21072 49568 21078
rect 49516 21014 49568 21020
rect 49384 20896 49464 20924
rect 49332 20878 49384 20884
rect 49240 20800 49292 20806
rect 49146 20768 49202 20777
rect 49240 20742 49292 20748
rect 49146 20703 49202 20712
rect 49332 20596 49384 20602
rect 49528 20584 49556 21014
rect 49620 20602 49648 22086
rect 49804 22001 49832 25094
rect 49896 24274 49924 27066
rect 49976 26376 50028 26382
rect 49976 26318 50028 26324
rect 49988 26246 50016 26318
rect 49976 26240 50028 26246
rect 49976 26182 50028 26188
rect 49976 25696 50028 25702
rect 49976 25638 50028 25644
rect 49988 24954 50016 25638
rect 49976 24948 50028 24954
rect 49976 24890 50028 24896
rect 49976 24812 50028 24818
rect 49976 24754 50028 24760
rect 49884 24268 49936 24274
rect 49884 24210 49936 24216
rect 49988 24138 50016 24754
rect 49976 24132 50028 24138
rect 49976 24074 50028 24080
rect 49976 23792 50028 23798
rect 49976 23734 50028 23740
rect 49884 23724 49936 23730
rect 49884 23666 49936 23672
rect 49896 23322 49924 23666
rect 49884 23316 49936 23322
rect 49884 23258 49936 23264
rect 49884 23112 49936 23118
rect 49884 23054 49936 23060
rect 49790 21992 49846 22001
rect 49712 21950 49790 21978
rect 49332 20538 49384 20544
rect 49436 20556 49556 20584
rect 49608 20596 49660 20602
rect 49344 20466 49372 20538
rect 49332 20460 49384 20466
rect 49332 20402 49384 20408
rect 49436 20398 49464 20556
rect 49608 20538 49660 20544
rect 49514 20496 49570 20505
rect 49514 20431 49570 20440
rect 49424 20392 49476 20398
rect 49424 20334 49476 20340
rect 49528 20330 49556 20431
rect 49516 20324 49568 20330
rect 49516 20266 49568 20272
rect 49238 20224 49294 20233
rect 49238 20159 49294 20168
rect 49252 20058 49280 20159
rect 48962 20023 49018 20032
rect 49056 20052 49108 20058
rect 49056 19994 49108 20000
rect 49240 20052 49292 20058
rect 49240 19994 49292 20000
rect 49056 19848 49108 19854
rect 49056 19790 49108 19796
rect 49068 19689 49096 19790
rect 49054 19680 49110 19689
rect 49054 19615 49110 19624
rect 49252 19281 49280 19994
rect 49424 19848 49476 19854
rect 49424 19790 49476 19796
rect 49332 19508 49384 19514
rect 49332 19450 49384 19456
rect 49238 19272 49294 19281
rect 48884 19230 49004 19258
rect 48976 18766 49004 19230
rect 49238 19207 49294 19216
rect 49148 19168 49200 19174
rect 49148 19110 49200 19116
rect 49240 19168 49292 19174
rect 49240 19110 49292 19116
rect 49056 18964 49108 18970
rect 49056 18906 49108 18912
rect 49068 18766 49096 18906
rect 48964 18760 49016 18766
rect 48964 18702 49016 18708
rect 49056 18760 49108 18766
rect 49056 18702 49108 18708
rect 48976 18630 49004 18702
rect 48964 18624 49016 18630
rect 48964 18566 49016 18572
rect 49068 18222 49096 18702
rect 49056 18216 49108 18222
rect 49056 18158 49108 18164
rect 48778 17912 48834 17921
rect 48778 17847 48834 17856
rect 48792 17241 48820 17847
rect 48964 17740 49016 17746
rect 48964 17682 49016 17688
rect 48778 17232 48834 17241
rect 48778 17167 48834 17176
rect 48872 17196 48924 17202
rect 48872 17138 48924 17144
rect 48780 17128 48832 17134
rect 48780 17070 48832 17076
rect 48648 16408 48728 16436
rect 48596 16390 48648 16396
rect 48594 16280 48650 16289
rect 48594 16215 48650 16224
rect 48608 16114 48636 16215
rect 48596 16108 48648 16114
rect 48596 16050 48648 16056
rect 48688 16108 48740 16114
rect 48688 16050 48740 16056
rect 48608 15638 48636 16050
rect 48700 15638 48728 16050
rect 48792 15706 48820 17070
rect 48884 16794 48912 17138
rect 48872 16788 48924 16794
rect 48872 16730 48924 16736
rect 48872 16584 48924 16590
rect 48872 16526 48924 16532
rect 48884 16096 48912 16526
rect 48976 16232 49004 17682
rect 49056 17672 49108 17678
rect 49056 17614 49108 17620
rect 49068 17338 49096 17614
rect 49056 17332 49108 17338
rect 49056 17274 49108 17280
rect 49056 17196 49108 17202
rect 49056 17138 49108 17144
rect 49068 16969 49096 17138
rect 49054 16960 49110 16969
rect 49054 16895 49110 16904
rect 49160 16708 49188 19110
rect 49252 18902 49280 19110
rect 49240 18896 49292 18902
rect 49240 18838 49292 18844
rect 49344 18578 49372 19450
rect 49436 19310 49464 19790
rect 49516 19712 49568 19718
rect 49516 19654 49568 19660
rect 49528 19514 49556 19654
rect 49516 19508 49568 19514
rect 49516 19450 49568 19456
rect 49620 19334 49648 20538
rect 49712 19394 49740 21950
rect 49790 21927 49846 21936
rect 49792 21888 49844 21894
rect 49792 21830 49844 21836
rect 49804 21321 49832 21830
rect 49790 21312 49846 21321
rect 49790 21247 49846 21256
rect 49804 20942 49832 21247
rect 49792 20936 49844 20942
rect 49792 20878 49844 20884
rect 49792 20800 49844 20806
rect 49792 20742 49844 20748
rect 49804 19825 49832 20742
rect 49896 20534 49924 23054
rect 49988 20942 50016 23734
rect 50080 23497 50108 27814
rect 50436 27396 50488 27402
rect 50436 27338 50488 27344
rect 50528 27396 50580 27402
rect 50528 27338 50580 27344
rect 50448 27130 50476 27338
rect 50436 27124 50488 27130
rect 50436 27066 50488 27072
rect 50540 26994 50568 27338
rect 50528 26988 50580 26994
rect 50528 26930 50580 26936
rect 50632 26926 50660 28494
rect 50896 28008 50948 28014
rect 50896 27950 50948 27956
rect 50804 26988 50856 26994
rect 50804 26930 50856 26936
rect 50620 26920 50672 26926
rect 50620 26862 50672 26868
rect 50632 26602 50660 26862
rect 50540 26574 50660 26602
rect 50816 26586 50844 26930
rect 50804 26580 50856 26586
rect 50434 26480 50490 26489
rect 50434 26415 50436 26424
rect 50488 26415 50490 26424
rect 50436 26386 50488 26392
rect 50540 26382 50568 26574
rect 50804 26522 50856 26528
rect 50620 26512 50672 26518
rect 50620 26454 50672 26460
rect 50528 26376 50580 26382
rect 50528 26318 50580 26324
rect 50436 26308 50488 26314
rect 50436 26250 50488 26256
rect 50448 26042 50476 26250
rect 50436 26036 50488 26042
rect 50436 25978 50488 25984
rect 50540 25974 50568 26318
rect 50528 25968 50580 25974
rect 50528 25910 50580 25916
rect 50344 25900 50396 25906
rect 50344 25842 50396 25848
rect 50160 25832 50212 25838
rect 50160 25774 50212 25780
rect 50172 25498 50200 25774
rect 50160 25492 50212 25498
rect 50160 25434 50212 25440
rect 50252 25424 50304 25430
rect 50252 25366 50304 25372
rect 50160 25288 50212 25294
rect 50158 25256 50160 25265
rect 50212 25256 50214 25265
rect 50158 25191 50214 25200
rect 50160 24880 50212 24886
rect 50160 24822 50212 24828
rect 50066 23488 50122 23497
rect 50066 23423 50122 23432
rect 50172 22386 50200 24822
rect 50264 24818 50292 25366
rect 50252 24812 50304 24818
rect 50252 24754 50304 24760
rect 50356 23594 50384 25842
rect 50434 25800 50490 25809
rect 50434 25735 50436 25744
rect 50488 25735 50490 25744
rect 50436 25706 50488 25712
rect 50540 24954 50568 25910
rect 50632 25294 50660 26454
rect 50712 25832 50764 25838
rect 50712 25774 50764 25780
rect 50724 25294 50752 25774
rect 50620 25288 50672 25294
rect 50620 25230 50672 25236
rect 50712 25288 50764 25294
rect 50712 25230 50764 25236
rect 50802 25256 50858 25265
rect 50802 25191 50858 25200
rect 50816 25158 50844 25191
rect 50804 25152 50856 25158
rect 50804 25094 50856 25100
rect 50528 24948 50580 24954
rect 50528 24890 50580 24896
rect 50712 24880 50764 24886
rect 50710 24848 50712 24857
rect 50764 24848 50766 24857
rect 50620 24812 50672 24818
rect 50540 24772 50620 24800
rect 50540 24410 50568 24772
rect 50710 24783 50766 24792
rect 50620 24754 50672 24760
rect 50908 24682 50936 27950
rect 52460 27668 52512 27674
rect 52460 27610 52512 27616
rect 50988 27532 51040 27538
rect 50988 27474 51040 27480
rect 51908 27532 51960 27538
rect 51908 27474 51960 27480
rect 51000 26790 51028 27474
rect 50988 26784 51040 26790
rect 50988 26726 51040 26732
rect 51000 26450 51028 26726
rect 51920 26518 51948 27474
rect 52000 27328 52052 27334
rect 52000 27270 52052 27276
rect 52012 26994 52040 27270
rect 52472 27130 52500 27610
rect 52460 27124 52512 27130
rect 52460 27066 52512 27072
rect 53288 27056 53340 27062
rect 53288 26998 53340 27004
rect 52000 26988 52052 26994
rect 52000 26930 52052 26936
rect 53012 26920 53064 26926
rect 53012 26862 53064 26868
rect 52184 26852 52236 26858
rect 52184 26794 52236 26800
rect 51908 26512 51960 26518
rect 51908 26454 51960 26460
rect 50988 26444 51040 26450
rect 50988 26386 51040 26392
rect 50896 24676 50948 24682
rect 50896 24618 50948 24624
rect 51000 24410 51028 26386
rect 51920 25974 51948 26454
rect 51908 25968 51960 25974
rect 51908 25910 51960 25916
rect 51356 25900 51408 25906
rect 51356 25842 51408 25848
rect 51632 25900 51684 25906
rect 51632 25842 51684 25848
rect 51368 25702 51396 25842
rect 51356 25696 51408 25702
rect 51356 25638 51408 25644
rect 51368 24818 51396 25638
rect 51356 24812 51408 24818
rect 51356 24754 51408 24760
rect 51644 24750 51672 25842
rect 51816 25696 51868 25702
rect 51816 25638 51868 25644
rect 51828 25294 51856 25638
rect 52196 25362 52224 26794
rect 53024 26586 53052 26862
rect 53012 26580 53064 26586
rect 53012 26522 53064 26528
rect 52644 26376 52696 26382
rect 52644 26318 52696 26324
rect 52656 26042 52684 26318
rect 53012 26240 53064 26246
rect 53012 26182 53064 26188
rect 52644 26036 52696 26042
rect 52644 25978 52696 25984
rect 53024 25974 53052 26182
rect 53012 25968 53064 25974
rect 53012 25910 53064 25916
rect 52644 25900 52696 25906
rect 52644 25842 52696 25848
rect 52656 25498 52684 25842
rect 52644 25492 52696 25498
rect 52644 25434 52696 25440
rect 52184 25356 52236 25362
rect 52184 25298 52236 25304
rect 51816 25288 51868 25294
rect 51816 25230 51868 25236
rect 52000 25288 52052 25294
rect 52000 25230 52052 25236
rect 52012 24954 52040 25230
rect 52000 24948 52052 24954
rect 52000 24890 52052 24896
rect 51632 24744 51684 24750
rect 51632 24686 51684 24692
rect 50528 24404 50580 24410
rect 50528 24346 50580 24352
rect 50988 24404 51040 24410
rect 50988 24346 51040 24352
rect 50344 23588 50396 23594
rect 50344 23530 50396 23536
rect 50080 22358 50200 22386
rect 49976 20936 50028 20942
rect 49976 20878 50028 20884
rect 49988 20534 50016 20878
rect 49884 20528 49936 20534
rect 49884 20470 49936 20476
rect 49976 20528 50028 20534
rect 49976 20470 50028 20476
rect 49896 20058 49924 20470
rect 49884 20052 49936 20058
rect 49884 19994 49936 20000
rect 49790 19816 49846 19825
rect 49790 19751 49846 19760
rect 49792 19712 49844 19718
rect 49790 19680 49792 19689
rect 49844 19680 49846 19689
rect 49790 19615 49846 19624
rect 49884 19508 49936 19514
rect 49884 19450 49936 19456
rect 49712 19366 49832 19394
rect 49424 19304 49476 19310
rect 49424 19246 49476 19252
rect 49528 19306 49648 19334
rect 49436 18698 49464 19246
rect 49424 18692 49476 18698
rect 49424 18634 49476 18640
rect 49344 18550 49464 18578
rect 49332 17876 49384 17882
rect 49332 17818 49384 17824
rect 49344 17202 49372 17818
rect 49332 17196 49384 17202
rect 49332 17138 49384 17144
rect 49068 16680 49188 16708
rect 49068 16522 49096 16680
rect 49436 16590 49464 18550
rect 49528 17954 49556 19306
rect 49700 19304 49752 19310
rect 49700 19246 49752 19252
rect 49608 19236 49660 19242
rect 49608 19178 49660 19184
rect 49620 18902 49648 19178
rect 49712 18970 49740 19246
rect 49700 18964 49752 18970
rect 49700 18906 49752 18912
rect 49608 18896 49660 18902
rect 49608 18838 49660 18844
rect 49528 17926 49648 17954
rect 49516 17876 49568 17882
rect 49516 17818 49568 17824
rect 49528 17338 49556 17818
rect 49516 17332 49568 17338
rect 49516 17274 49568 17280
rect 49620 16590 49648 17926
rect 49712 17814 49740 18906
rect 49700 17808 49752 17814
rect 49700 17750 49752 17756
rect 49700 17672 49752 17678
rect 49700 17614 49752 17620
rect 49712 17338 49740 17614
rect 49804 17338 49832 19366
rect 49700 17332 49752 17338
rect 49700 17274 49752 17280
rect 49792 17332 49844 17338
rect 49792 17274 49844 17280
rect 49896 17218 49924 19450
rect 49988 19394 50016 20470
rect 50080 20466 50108 22358
rect 50252 22092 50304 22098
rect 50540 22094 50568 24346
rect 50712 24336 50764 24342
rect 50712 24278 50764 24284
rect 50724 24206 50752 24278
rect 50712 24200 50764 24206
rect 50712 24142 50764 24148
rect 50804 24200 50856 24206
rect 50804 24142 50856 24148
rect 50712 24064 50764 24070
rect 50712 24006 50764 24012
rect 50724 23798 50752 24006
rect 50712 23792 50764 23798
rect 50712 23734 50764 23740
rect 50816 23322 50844 24142
rect 50804 23316 50856 23322
rect 50804 23258 50856 23264
rect 50712 23112 50764 23118
rect 50712 23054 50764 23060
rect 50252 22034 50304 22040
rect 50448 22066 50568 22094
rect 50264 21486 50292 22034
rect 50252 21480 50304 21486
rect 50252 21422 50304 21428
rect 50158 21040 50214 21049
rect 50158 20975 50214 20984
rect 50172 20874 50200 20975
rect 50160 20868 50212 20874
rect 50160 20810 50212 20816
rect 50264 20806 50292 21422
rect 50252 20800 50304 20806
rect 50252 20742 50304 20748
rect 50158 20632 50214 20641
rect 50158 20567 50214 20576
rect 50068 20460 50120 20466
rect 50068 20402 50120 20408
rect 50080 19514 50108 20402
rect 50068 19508 50120 19514
rect 50068 19450 50120 19456
rect 49988 19366 50108 19394
rect 49976 19304 50028 19310
rect 49976 19246 50028 19252
rect 49988 18970 50016 19246
rect 49976 18964 50028 18970
rect 49976 18906 50028 18912
rect 49976 18284 50028 18290
rect 49976 18226 50028 18232
rect 49988 17746 50016 18226
rect 49976 17740 50028 17746
rect 49976 17682 50028 17688
rect 50080 17270 50108 19366
rect 50068 17264 50120 17270
rect 49804 17190 49924 17218
rect 49974 17232 50030 17241
rect 49804 17134 49832 17190
rect 50068 17206 50120 17212
rect 49974 17167 50030 17176
rect 49792 17128 49844 17134
rect 49792 17070 49844 17076
rect 49332 16584 49384 16590
rect 49332 16526 49384 16532
rect 49424 16584 49476 16590
rect 49424 16526 49476 16532
rect 49608 16584 49660 16590
rect 49608 16526 49660 16532
rect 49056 16516 49108 16522
rect 49056 16458 49108 16464
rect 49148 16516 49200 16522
rect 49148 16458 49200 16464
rect 48976 16204 49096 16232
rect 48964 16108 49016 16114
rect 48884 16068 48964 16096
rect 48964 16050 49016 16056
rect 49068 15978 49096 16204
rect 49056 15972 49108 15978
rect 49056 15914 49108 15920
rect 48780 15700 48832 15706
rect 48780 15642 48832 15648
rect 48596 15632 48648 15638
rect 48596 15574 48648 15580
rect 48688 15632 48740 15638
rect 48688 15574 48740 15580
rect 48780 15496 48832 15502
rect 49160 15450 49188 16458
rect 49240 15700 49292 15706
rect 49240 15642 49292 15648
rect 48780 15438 48832 15444
rect 48688 15360 48740 15366
rect 48688 15302 48740 15308
rect 48502 15056 48558 15065
rect 48502 14991 48558 15000
rect 48700 14929 48728 15302
rect 48410 14920 48466 14929
rect 48410 14855 48466 14864
rect 48686 14920 48742 14929
rect 48686 14855 48742 14864
rect 48424 14822 48452 14855
rect 48280 14764 48360 14770
rect 48228 14758 48360 14764
rect 48413 14816 48465 14822
rect 48413 14758 48465 14764
rect 48502 14784 48558 14793
rect 48240 14742 48360 14758
rect 48228 14476 48280 14482
rect 48228 14418 48280 14424
rect 48240 13326 48268 14418
rect 48332 13938 48360 14742
rect 48502 14719 48558 14728
rect 48320 13932 48372 13938
rect 48320 13874 48372 13880
rect 48332 13394 48360 13874
rect 48516 13530 48544 14719
rect 48792 14618 48820 15438
rect 48976 15422 49188 15450
rect 48780 14612 48832 14618
rect 48780 14554 48832 14560
rect 48976 14550 49004 15422
rect 49056 15360 49108 15366
rect 49056 15302 49108 15308
rect 48964 14544 49016 14550
rect 48964 14486 49016 14492
rect 48976 14414 49004 14486
rect 48780 14408 48832 14414
rect 48778 14376 48780 14385
rect 48964 14408 49016 14414
rect 48832 14376 48834 14385
rect 48964 14350 49016 14356
rect 48778 14311 48834 14320
rect 48596 14272 48648 14278
rect 48596 14214 48648 14220
rect 48608 13870 48636 14214
rect 49068 13977 49096 15302
rect 49252 14618 49280 15642
rect 49344 15434 49372 16526
rect 49436 16114 49464 16526
rect 49620 16250 49648 16526
rect 49698 16280 49754 16289
rect 49608 16244 49660 16250
rect 49698 16215 49700 16224
rect 49608 16186 49660 16192
rect 49752 16215 49754 16224
rect 49700 16186 49752 16192
rect 49712 16114 49740 16186
rect 49424 16108 49476 16114
rect 49424 16050 49476 16056
rect 49700 16108 49752 16114
rect 49700 16050 49752 16056
rect 49884 15564 49936 15570
rect 49884 15506 49936 15512
rect 49332 15428 49384 15434
rect 49332 15370 49384 15376
rect 49240 14612 49292 14618
rect 49240 14554 49292 14560
rect 49148 14272 49200 14278
rect 49148 14214 49200 14220
rect 49054 13968 49110 13977
rect 48780 13932 48832 13938
rect 49160 13938 49188 14214
rect 49054 13903 49056 13912
rect 48780 13874 48832 13880
rect 49108 13903 49110 13912
rect 49148 13932 49200 13938
rect 49056 13874 49108 13880
rect 49148 13874 49200 13880
rect 48596 13864 48648 13870
rect 48596 13806 48648 13812
rect 48688 13728 48740 13734
rect 48688 13670 48740 13676
rect 48504 13524 48556 13530
rect 48504 13466 48556 13472
rect 48320 13388 48372 13394
rect 48320 13330 48372 13336
rect 48136 13320 48188 13326
rect 48136 13262 48188 13268
rect 48228 13320 48280 13326
rect 48228 13262 48280 13268
rect 47308 13252 47360 13258
rect 47308 13194 47360 13200
rect 47320 12918 47348 13194
rect 46756 12912 46808 12918
rect 46756 12854 46808 12860
rect 47308 12912 47360 12918
rect 47308 12854 47360 12860
rect 46572 12640 46624 12646
rect 46572 12582 46624 12588
rect 46768 12442 46796 12854
rect 48148 12782 48176 13262
rect 48516 13258 48544 13466
rect 48700 13326 48728 13670
rect 48792 13530 48820 13874
rect 49252 13734 49280 14554
rect 49344 14396 49372 15370
rect 49896 15162 49924 15506
rect 49988 15162 50016 17167
rect 50080 16726 50108 17206
rect 50068 16720 50120 16726
rect 50068 16662 50120 16668
rect 50172 16232 50200 20567
rect 50448 20262 50476 22066
rect 50724 21321 50752 23054
rect 50804 23044 50856 23050
rect 50804 22986 50856 22992
rect 50816 21690 50844 22986
rect 51000 22506 51028 24346
rect 52368 24268 52420 24274
rect 52368 24210 52420 24216
rect 52184 24200 52236 24206
rect 52184 24142 52236 24148
rect 52196 23866 52224 24142
rect 52184 23860 52236 23866
rect 52184 23802 52236 23808
rect 51448 23792 51500 23798
rect 51448 23734 51500 23740
rect 50988 22500 51040 22506
rect 50988 22442 51040 22448
rect 51356 21888 51408 21894
rect 51356 21830 51408 21836
rect 50804 21684 50856 21690
rect 50804 21626 50856 21632
rect 50988 21480 51040 21486
rect 50988 21422 51040 21428
rect 50710 21312 50766 21321
rect 50710 21247 50766 21256
rect 51000 21146 51028 21422
rect 51262 21176 51318 21185
rect 50988 21140 51040 21146
rect 51262 21111 51264 21120
rect 50988 21082 51040 21088
rect 51316 21111 51318 21120
rect 51264 21082 51316 21088
rect 50802 21040 50858 21049
rect 51368 21010 51396 21830
rect 51460 21622 51488 23734
rect 52380 23254 52408 24210
rect 52656 23662 52684 25434
rect 52828 25356 52880 25362
rect 52828 25298 52880 25304
rect 52840 24818 52868 25298
rect 52828 24812 52880 24818
rect 52828 24754 52880 24760
rect 53300 23798 53328 26998
rect 54484 26784 54536 26790
rect 54484 26726 54536 26732
rect 54496 26382 54524 26726
rect 57888 26512 57940 26518
rect 57888 26454 57940 26460
rect 54484 26376 54536 26382
rect 54484 26318 54536 26324
rect 54208 25968 54260 25974
rect 57900 25945 57928 26454
rect 58256 26376 58308 26382
rect 58256 26318 58308 26324
rect 54208 25910 54260 25916
rect 56690 25936 56746 25945
rect 53472 25900 53524 25906
rect 53472 25842 53524 25848
rect 53748 25900 53800 25906
rect 53748 25842 53800 25848
rect 53484 25362 53512 25842
rect 53472 25356 53524 25362
rect 53472 25298 53524 25304
rect 53380 25152 53432 25158
rect 53380 25094 53432 25100
rect 53392 24750 53420 25094
rect 53484 24818 53512 25298
rect 53760 25226 53788 25842
rect 54220 25226 54248 25910
rect 57886 25936 57942 25945
rect 56690 25871 56692 25880
rect 56744 25871 56746 25880
rect 56876 25900 56928 25906
rect 56692 25842 56744 25848
rect 57886 25871 57942 25880
rect 56876 25842 56928 25848
rect 55312 25832 55364 25838
rect 55312 25774 55364 25780
rect 55956 25832 56008 25838
rect 55956 25774 56008 25780
rect 56232 25832 56284 25838
rect 56232 25774 56284 25780
rect 55324 25294 55352 25774
rect 55968 25498 55996 25774
rect 55956 25492 56008 25498
rect 55956 25434 56008 25440
rect 56244 25430 56272 25774
rect 56508 25696 56560 25702
rect 56508 25638 56560 25644
rect 56232 25424 56284 25430
rect 56232 25366 56284 25372
rect 55312 25288 55364 25294
rect 55312 25230 55364 25236
rect 53748 25220 53800 25226
rect 53748 25162 53800 25168
rect 53840 25220 53892 25226
rect 53840 25162 53892 25168
rect 54208 25220 54260 25226
rect 54208 25162 54260 25168
rect 53472 24812 53524 24818
rect 53472 24754 53524 24760
rect 53380 24744 53432 24750
rect 53380 24686 53432 24692
rect 53380 24132 53432 24138
rect 53380 24074 53432 24080
rect 53392 23866 53420 24074
rect 53380 23860 53432 23866
rect 53380 23802 53432 23808
rect 53288 23792 53340 23798
rect 53288 23734 53340 23740
rect 52644 23656 52696 23662
rect 52644 23598 52696 23604
rect 52368 23248 52420 23254
rect 52368 23190 52420 23196
rect 51908 22976 51960 22982
rect 52460 22976 52512 22982
rect 51908 22918 51960 22924
rect 52380 22924 52460 22930
rect 52380 22918 52512 22924
rect 51920 22642 51948 22918
rect 52380 22902 52500 22918
rect 51908 22636 51960 22642
rect 51908 22578 51960 22584
rect 52092 21888 52144 21894
rect 52092 21830 52144 21836
rect 52000 21684 52052 21690
rect 52104 21672 52132 21830
rect 52052 21644 52132 21672
rect 52000 21626 52052 21632
rect 51448 21616 51500 21622
rect 51448 21558 51500 21564
rect 51460 21332 51488 21558
rect 51540 21344 51592 21350
rect 51460 21304 51540 21332
rect 50802 20975 50858 20984
rect 51356 21004 51408 21010
rect 50816 20942 50844 20975
rect 51356 20946 51408 20952
rect 50528 20936 50580 20942
rect 50528 20878 50580 20884
rect 50804 20936 50856 20942
rect 50804 20878 50856 20884
rect 50540 20466 50568 20878
rect 51264 20868 51316 20874
rect 51264 20810 51316 20816
rect 51276 20777 51304 20810
rect 51262 20768 51318 20777
rect 51262 20703 51318 20712
rect 50528 20460 50580 20466
rect 50528 20402 50580 20408
rect 50896 20392 50948 20398
rect 50896 20334 50948 20340
rect 50436 20256 50488 20262
rect 50436 20198 50488 20204
rect 50448 20058 50476 20198
rect 50436 20052 50488 20058
rect 50436 19994 50488 20000
rect 50448 19854 50476 19994
rect 50908 19854 50936 20334
rect 51264 20052 51316 20058
rect 51264 19994 51316 20000
rect 50988 19984 51040 19990
rect 50988 19926 51040 19932
rect 51000 19854 51028 19926
rect 50436 19848 50488 19854
rect 50436 19790 50488 19796
rect 50712 19848 50764 19854
rect 50712 19790 50764 19796
rect 50896 19848 50948 19854
rect 50896 19790 50948 19796
rect 50988 19848 51040 19854
rect 50988 19790 51040 19796
rect 50436 19712 50488 19718
rect 50436 19654 50488 19660
rect 50252 19440 50304 19446
rect 50304 19400 50384 19428
rect 50252 19382 50304 19388
rect 50356 18766 50384 19400
rect 50344 18760 50396 18766
rect 50344 18702 50396 18708
rect 50252 18284 50304 18290
rect 50252 18226 50304 18232
rect 50264 17202 50292 18226
rect 50356 17320 50384 18702
rect 50448 18290 50476 19654
rect 50528 18352 50580 18358
rect 50528 18294 50580 18300
rect 50436 18284 50488 18290
rect 50436 18226 50488 18232
rect 50356 17292 50476 17320
rect 50252 17196 50304 17202
rect 50252 17138 50304 17144
rect 50344 17196 50396 17202
rect 50344 17138 50396 17144
rect 50356 16522 50384 17138
rect 50448 17105 50476 17292
rect 50434 17096 50490 17105
rect 50434 17031 50490 17040
rect 50344 16516 50396 16522
rect 50344 16458 50396 16464
rect 50252 16244 50304 16250
rect 50172 16204 50252 16232
rect 50068 16108 50120 16114
rect 50068 16050 50120 16056
rect 49884 15156 49936 15162
rect 49712 15116 49884 15144
rect 49712 14958 49740 15116
rect 49884 15098 49936 15104
rect 49976 15156 50028 15162
rect 49976 15098 50028 15104
rect 49700 14952 49752 14958
rect 49700 14894 49752 14900
rect 49608 14408 49660 14414
rect 49344 14368 49608 14396
rect 49608 14350 49660 14356
rect 49712 14278 49740 14894
rect 49792 14476 49844 14482
rect 49792 14418 49844 14424
rect 49804 14278 49832 14418
rect 49988 14414 50016 15098
rect 50080 14958 50108 16050
rect 50172 16046 50200 16204
rect 50252 16186 50304 16192
rect 50540 16130 50568 18294
rect 50620 18284 50672 18290
rect 50620 18226 50672 18232
rect 50632 18068 50660 18226
rect 50724 18170 50752 19790
rect 51080 19780 51132 19786
rect 51132 19740 51212 19768
rect 51080 19722 51132 19728
rect 51184 19310 51212 19740
rect 51172 19304 51224 19310
rect 51172 19246 51224 19252
rect 51080 18692 51132 18698
rect 51080 18634 51132 18640
rect 50724 18142 51028 18170
rect 50896 18080 50948 18086
rect 50632 18040 50752 18068
rect 50620 17604 50672 17610
rect 50620 17546 50672 17552
rect 50632 17338 50660 17546
rect 50620 17332 50672 17338
rect 50620 17274 50672 17280
rect 50448 16102 50568 16130
rect 50160 16040 50212 16046
rect 50160 15982 50212 15988
rect 50068 14952 50120 14958
rect 50068 14894 50120 14900
rect 50080 14414 50108 14894
rect 49976 14408 50028 14414
rect 49976 14350 50028 14356
rect 50068 14408 50120 14414
rect 50448 14385 50476 16102
rect 50618 15328 50674 15337
rect 50724 15314 50752 18040
rect 50896 18022 50948 18028
rect 50908 17202 50936 18022
rect 50804 17196 50856 17202
rect 50804 17138 50856 17144
rect 50896 17196 50948 17202
rect 50896 17138 50948 17144
rect 50816 17105 50844 17138
rect 50802 17096 50858 17105
rect 50802 17031 50858 17040
rect 50816 15473 50844 17031
rect 50802 15464 50858 15473
rect 50802 15399 50858 15408
rect 50674 15286 50752 15314
rect 50618 15263 50674 15272
rect 50632 14414 50660 15263
rect 50528 14408 50580 14414
rect 50068 14350 50120 14356
rect 50434 14376 50490 14385
rect 50528 14350 50580 14356
rect 50620 14408 50672 14414
rect 50620 14350 50672 14356
rect 50434 14311 50436 14320
rect 50488 14311 50490 14320
rect 50436 14282 50488 14288
rect 49700 14272 49752 14278
rect 49700 14214 49752 14220
rect 49792 14272 49844 14278
rect 49792 14214 49844 14220
rect 50540 13938 50568 14350
rect 50804 14272 50856 14278
rect 50804 14214 50856 14220
rect 50816 14006 50844 14214
rect 50804 14000 50856 14006
rect 50804 13942 50856 13948
rect 49792 13932 49844 13938
rect 49792 13874 49844 13880
rect 50528 13932 50580 13938
rect 50528 13874 50580 13880
rect 49056 13728 49108 13734
rect 49056 13670 49108 13676
rect 49240 13728 49292 13734
rect 49240 13670 49292 13676
rect 48780 13524 48832 13530
rect 48780 13466 48832 13472
rect 48688 13320 48740 13326
rect 48688 13262 48740 13268
rect 48504 13252 48556 13258
rect 48504 13194 48556 13200
rect 49068 12918 49096 13670
rect 49804 13394 49832 13874
rect 49792 13388 49844 13394
rect 49792 13330 49844 13336
rect 49804 12986 49832 13330
rect 50160 13252 50212 13258
rect 50160 13194 50212 13200
rect 49792 12980 49844 12986
rect 49792 12922 49844 12928
rect 49056 12912 49108 12918
rect 49056 12854 49108 12860
rect 50172 12850 50200 13194
rect 50540 12986 50568 13874
rect 51000 13870 51028 18142
rect 51092 16998 51120 18634
rect 51276 18358 51304 19994
rect 51460 19446 51488 21304
rect 51540 21286 51592 21292
rect 51724 21344 51776 21350
rect 51724 21286 51776 21292
rect 51736 19922 51764 21286
rect 52104 20942 52132 21644
rect 52380 21418 52408 22902
rect 52656 21894 52684 23598
rect 52920 23044 52972 23050
rect 52920 22986 52972 22992
rect 52932 22166 52960 22986
rect 53300 22778 53328 23734
rect 53380 23044 53432 23050
rect 53380 22986 53432 22992
rect 53392 22778 53420 22986
rect 53288 22772 53340 22778
rect 53288 22714 53340 22720
rect 53380 22772 53432 22778
rect 53380 22714 53432 22720
rect 52920 22160 52972 22166
rect 52920 22102 52972 22108
rect 52644 21888 52696 21894
rect 52644 21830 52696 21836
rect 52550 21584 52606 21593
rect 52460 21548 52512 21554
rect 52550 21519 52606 21528
rect 52460 21490 52512 21496
rect 52368 21412 52420 21418
rect 52368 21354 52420 21360
rect 52184 21344 52236 21350
rect 52184 21286 52236 21292
rect 52196 21146 52224 21286
rect 52472 21146 52500 21490
rect 52184 21140 52236 21146
rect 52184 21082 52236 21088
rect 52460 21140 52512 21146
rect 52460 21082 52512 21088
rect 51908 20936 51960 20942
rect 51828 20896 51908 20924
rect 51828 20806 51856 20896
rect 51908 20878 51960 20884
rect 52092 20936 52144 20942
rect 52184 20936 52236 20942
rect 52092 20878 52144 20884
rect 52182 20904 52184 20913
rect 52460 20936 52512 20942
rect 52236 20904 52238 20913
rect 52460 20878 52512 20884
rect 52182 20839 52238 20848
rect 51816 20800 51868 20806
rect 51816 20742 51868 20748
rect 52472 20534 52500 20878
rect 52460 20528 52512 20534
rect 52460 20470 52512 20476
rect 51724 19916 51776 19922
rect 51724 19858 51776 19864
rect 51724 19780 51776 19786
rect 51724 19722 51776 19728
rect 51356 19440 51408 19446
rect 51356 19382 51408 19388
rect 51448 19440 51500 19446
rect 51448 19382 51500 19388
rect 51264 18352 51316 18358
rect 51264 18294 51316 18300
rect 51170 17776 51226 17785
rect 51170 17711 51226 17720
rect 51080 16992 51132 16998
rect 51080 16934 51132 16940
rect 51080 16040 51132 16046
rect 51080 15982 51132 15988
rect 51092 14074 51120 15982
rect 51184 14074 51212 17711
rect 51368 17610 51396 19382
rect 51540 19168 51592 19174
rect 51540 19110 51592 19116
rect 51552 18766 51580 19110
rect 51736 18970 51764 19722
rect 51816 19712 51868 19718
rect 51816 19654 51868 19660
rect 52092 19712 52144 19718
rect 52092 19654 52144 19660
rect 51724 18964 51776 18970
rect 51724 18906 51776 18912
rect 51828 18766 51856 19654
rect 52104 18766 52132 19654
rect 52564 18970 52592 21519
rect 52656 20942 52684 21830
rect 52644 20936 52696 20942
rect 52644 20878 52696 20884
rect 52932 19922 52960 22102
rect 53380 21888 53432 21894
rect 53380 21830 53432 21836
rect 53392 21690 53420 21830
rect 53380 21684 53432 21690
rect 53380 21626 53432 21632
rect 53484 20806 53512 24754
rect 53564 24200 53616 24206
rect 53564 24142 53616 24148
rect 53576 23730 53604 24142
rect 53564 23724 53616 23730
rect 53564 23666 53616 23672
rect 53760 23610 53788 25162
rect 53852 24342 53880 25162
rect 54116 24948 54168 24954
rect 54116 24890 54168 24896
rect 53840 24336 53892 24342
rect 53840 24278 53892 24284
rect 53852 24206 53880 24278
rect 54128 24274 54156 24890
rect 54220 24614 54248 25162
rect 55324 24954 55352 25230
rect 55680 25220 55732 25226
rect 55680 25162 55732 25168
rect 55312 24948 55364 24954
rect 55312 24890 55364 24896
rect 55692 24818 55720 25162
rect 56244 24886 56272 25366
rect 56416 25288 56468 25294
rect 56416 25230 56468 25236
rect 56232 24880 56284 24886
rect 56232 24822 56284 24828
rect 55404 24812 55456 24818
rect 55404 24754 55456 24760
rect 55680 24812 55732 24818
rect 55680 24754 55732 24760
rect 55312 24676 55364 24682
rect 55312 24618 55364 24624
rect 54208 24608 54260 24614
rect 54208 24550 54260 24556
rect 54116 24268 54168 24274
rect 54116 24210 54168 24216
rect 53840 24200 53892 24206
rect 53840 24142 53892 24148
rect 54024 24200 54076 24206
rect 54024 24142 54076 24148
rect 53668 23582 53788 23610
rect 53932 23656 53984 23662
rect 53932 23598 53984 23604
rect 53668 22982 53696 23582
rect 53748 23520 53800 23526
rect 53748 23462 53800 23468
rect 53838 23488 53894 23497
rect 53656 22976 53708 22982
rect 53656 22918 53708 22924
rect 53668 22710 53696 22918
rect 53656 22704 53708 22710
rect 53656 22646 53708 22652
rect 53564 22432 53616 22438
rect 53564 22374 53616 22380
rect 53576 21350 53604 22374
rect 53668 22166 53696 22646
rect 53760 22642 53788 23462
rect 53838 23423 53894 23432
rect 53852 23322 53880 23423
rect 53840 23316 53892 23322
rect 53840 23258 53892 23264
rect 53944 23118 53972 23598
rect 54036 23526 54064 24142
rect 54220 23866 54248 24550
rect 54392 24404 54444 24410
rect 54392 24346 54444 24352
rect 54404 24206 54432 24346
rect 55220 24268 55272 24274
rect 55220 24210 55272 24216
rect 54392 24200 54444 24206
rect 54392 24142 54444 24148
rect 54852 24200 54904 24206
rect 54852 24142 54904 24148
rect 54300 24064 54352 24070
rect 54300 24006 54352 24012
rect 54760 24064 54812 24070
rect 54760 24006 54812 24012
rect 54208 23860 54260 23866
rect 54208 23802 54260 23808
rect 54312 23662 54340 24006
rect 54668 23860 54720 23866
rect 54668 23802 54720 23808
rect 54300 23656 54352 23662
rect 54300 23598 54352 23604
rect 54024 23520 54076 23526
rect 54024 23462 54076 23468
rect 53932 23112 53984 23118
rect 53932 23054 53984 23060
rect 53748 22636 53800 22642
rect 53748 22578 53800 22584
rect 54392 22432 54444 22438
rect 54392 22374 54444 22380
rect 53656 22160 53708 22166
rect 53656 22102 53708 22108
rect 53668 21622 53696 22102
rect 54404 21690 54432 22374
rect 54484 22024 54536 22030
rect 54484 21966 54536 21972
rect 54392 21684 54444 21690
rect 54392 21626 54444 21632
rect 53656 21616 53708 21622
rect 53656 21558 53708 21564
rect 53564 21344 53616 21350
rect 53564 21286 53616 21292
rect 54404 20874 54432 21626
rect 54496 21554 54524 21966
rect 54680 21622 54708 23802
rect 54772 23798 54800 24006
rect 54760 23792 54812 23798
rect 54760 23734 54812 23740
rect 54864 22094 54892 24142
rect 54772 22066 54892 22094
rect 55232 22094 55260 24210
rect 55324 23866 55352 24618
rect 55312 23860 55364 23866
rect 55312 23802 55364 23808
rect 55416 23526 55444 24754
rect 56232 24744 56284 24750
rect 56232 24686 56284 24692
rect 55588 24676 55640 24682
rect 55588 24618 55640 24624
rect 55404 23520 55456 23526
rect 55404 23462 55456 23468
rect 55600 23118 55628 24618
rect 56244 24410 56272 24686
rect 56324 24608 56376 24614
rect 56324 24550 56376 24556
rect 56232 24404 56284 24410
rect 56232 24346 56284 24352
rect 56336 24206 56364 24550
rect 56428 24274 56456 25230
rect 56520 24886 56548 25638
rect 56704 24936 56732 25842
rect 56888 25809 56916 25842
rect 58268 25838 58296 26318
rect 58256 25832 58308 25838
rect 56874 25800 56930 25809
rect 58256 25774 58308 25780
rect 56874 25735 56930 25744
rect 57520 25696 57572 25702
rect 57520 25638 57572 25644
rect 57532 25294 57560 25638
rect 58268 25498 58296 25774
rect 58256 25492 58308 25498
rect 58256 25434 58308 25440
rect 57520 25288 57572 25294
rect 57520 25230 57572 25236
rect 56704 24908 56824 24936
rect 56508 24880 56560 24886
rect 56508 24822 56560 24828
rect 56416 24268 56468 24274
rect 56416 24210 56468 24216
rect 56324 24200 56376 24206
rect 56324 24142 56376 24148
rect 56520 24070 56548 24822
rect 56508 24064 56560 24070
rect 56508 24006 56560 24012
rect 56692 23656 56744 23662
rect 56692 23598 56744 23604
rect 55956 23520 56008 23526
rect 55956 23462 56008 23468
rect 55968 23186 55996 23462
rect 55956 23180 56008 23186
rect 55956 23122 56008 23128
rect 55588 23112 55640 23118
rect 56704 23089 56732 23598
rect 55588 23054 55640 23060
rect 56690 23080 56746 23089
rect 55600 22710 55628 23054
rect 56690 23015 56746 23024
rect 56600 22976 56652 22982
rect 56600 22918 56652 22924
rect 55588 22704 55640 22710
rect 55588 22646 55640 22652
rect 56140 22636 56192 22642
rect 56140 22578 56192 22584
rect 55864 22568 55916 22574
rect 55864 22510 55916 22516
rect 55232 22066 55352 22094
rect 54668 21616 54720 21622
rect 54668 21558 54720 21564
rect 54484 21548 54536 21554
rect 54484 21490 54536 21496
rect 54496 21350 54524 21490
rect 54576 21412 54628 21418
rect 54576 21354 54628 21360
rect 54484 21344 54536 21350
rect 54484 21286 54536 21292
rect 54496 21010 54524 21286
rect 54484 21004 54536 21010
rect 54484 20946 54536 20952
rect 54392 20868 54444 20874
rect 54392 20810 54444 20816
rect 53472 20800 53524 20806
rect 53472 20742 53524 20748
rect 54484 20800 54536 20806
rect 54484 20742 54536 20748
rect 53840 20460 53892 20466
rect 53840 20402 53892 20408
rect 53380 20324 53432 20330
rect 53380 20266 53432 20272
rect 53288 20256 53340 20262
rect 53288 20198 53340 20204
rect 52920 19916 52972 19922
rect 52920 19858 52972 19864
rect 52932 19514 52960 19858
rect 53300 19854 53328 20198
rect 53392 20097 53420 20266
rect 53656 20256 53708 20262
rect 53656 20198 53708 20204
rect 53378 20088 53434 20097
rect 53378 20023 53434 20032
rect 53392 19854 53420 20023
rect 53472 19916 53524 19922
rect 53472 19858 53524 19864
rect 53288 19848 53340 19854
rect 53288 19790 53340 19796
rect 53380 19848 53432 19854
rect 53380 19790 53432 19796
rect 53484 19718 53512 19858
rect 53472 19712 53524 19718
rect 53472 19654 53524 19660
rect 52920 19508 52972 19514
rect 52920 19450 52972 19456
rect 53668 19310 53696 20198
rect 53852 20058 53880 20402
rect 53932 20256 53984 20262
rect 53932 20198 53984 20204
rect 53840 20052 53892 20058
rect 53840 19994 53892 20000
rect 53944 19938 53972 20198
rect 53852 19910 53972 19938
rect 53748 19848 53800 19854
rect 53748 19790 53800 19796
rect 53656 19304 53708 19310
rect 53656 19246 53708 19252
rect 52552 18964 52604 18970
rect 52552 18906 52604 18912
rect 53288 18964 53340 18970
rect 53288 18906 53340 18912
rect 51540 18760 51592 18766
rect 51540 18702 51592 18708
rect 51816 18760 51868 18766
rect 51816 18702 51868 18708
rect 52092 18760 52144 18766
rect 52092 18702 52144 18708
rect 53012 18284 53064 18290
rect 53012 18226 53064 18232
rect 52736 18080 52788 18086
rect 52736 18022 52788 18028
rect 52828 18080 52880 18086
rect 52828 18022 52880 18028
rect 52748 17610 52776 18022
rect 51356 17604 51408 17610
rect 51356 17546 51408 17552
rect 52736 17604 52788 17610
rect 52736 17546 52788 17552
rect 51264 16992 51316 16998
rect 51264 16934 51316 16940
rect 51276 14618 51304 16934
rect 51368 16726 51396 17546
rect 52368 17536 52420 17542
rect 52840 17490 52868 18022
rect 52368 17478 52420 17484
rect 52380 17202 52408 17478
rect 52748 17462 52868 17490
rect 51632 17196 51684 17202
rect 51552 17156 51632 17184
rect 51552 17066 51580 17156
rect 51632 17138 51684 17144
rect 52368 17196 52420 17202
rect 52368 17138 52420 17144
rect 51540 17060 51592 17066
rect 51540 17002 51592 17008
rect 51816 17060 51868 17066
rect 51816 17002 51868 17008
rect 51356 16720 51408 16726
rect 51356 16662 51408 16668
rect 51356 16108 51408 16114
rect 51356 16050 51408 16056
rect 51368 15706 51396 16050
rect 51356 15700 51408 15706
rect 51356 15642 51408 15648
rect 51368 15502 51396 15642
rect 51356 15496 51408 15502
rect 51724 15496 51776 15502
rect 51356 15438 51408 15444
rect 51630 15464 51686 15473
rect 51828 15484 51856 17002
rect 51908 15632 51960 15638
rect 52460 15632 52512 15638
rect 51960 15580 52132 15586
rect 51908 15574 52132 15580
rect 52460 15574 52512 15580
rect 51920 15570 52132 15574
rect 51920 15564 52144 15570
rect 51920 15558 52092 15564
rect 52092 15506 52144 15512
rect 51776 15456 51856 15484
rect 51724 15438 51776 15444
rect 51630 15399 51686 15408
rect 51264 14612 51316 14618
rect 51264 14554 51316 14560
rect 51080 14068 51132 14074
rect 51080 14010 51132 14016
rect 51172 14068 51224 14074
rect 51172 14010 51224 14016
rect 51644 13977 51672 15399
rect 51724 15360 51776 15366
rect 51724 15302 51776 15308
rect 51736 14346 51764 15302
rect 51828 15026 51856 15456
rect 51908 15428 51960 15434
rect 51908 15370 51960 15376
rect 51816 15020 51868 15026
rect 51816 14962 51868 14968
rect 51816 14612 51868 14618
rect 51816 14554 51868 14560
rect 51724 14340 51776 14346
rect 51724 14282 51776 14288
rect 51630 13968 51686 13977
rect 51630 13903 51632 13912
rect 51684 13903 51686 13912
rect 51632 13874 51684 13880
rect 51828 13870 51856 14554
rect 51920 13938 51948 15370
rect 52366 15192 52422 15201
rect 52472 15162 52500 15574
rect 52552 15496 52604 15502
rect 52552 15438 52604 15444
rect 52366 15127 52422 15136
rect 52460 15156 52512 15162
rect 52380 15094 52408 15127
rect 52460 15098 52512 15104
rect 52368 15088 52420 15094
rect 52368 15030 52420 15036
rect 52000 14068 52052 14074
rect 52000 14010 52052 14016
rect 51908 13932 51960 13938
rect 51908 13874 51960 13880
rect 50988 13864 51040 13870
rect 50988 13806 51040 13812
rect 51816 13864 51868 13870
rect 51816 13806 51868 13812
rect 51724 13796 51776 13802
rect 51724 13738 51776 13744
rect 51448 13728 51500 13734
rect 51448 13670 51500 13676
rect 51460 13394 51488 13670
rect 51736 13462 51764 13738
rect 51920 13530 51948 13874
rect 52012 13530 52040 14010
rect 52380 14006 52408 15030
rect 52564 14958 52592 15438
rect 52748 15366 52776 17462
rect 53024 17338 53052 18226
rect 53104 17536 53156 17542
rect 53104 17478 53156 17484
rect 53012 17332 53064 17338
rect 53012 17274 53064 17280
rect 52920 17196 52972 17202
rect 52920 17138 52972 17144
rect 53012 17196 53064 17202
rect 53116 17184 53144 17478
rect 53064 17156 53144 17184
rect 53196 17196 53248 17202
rect 53012 17138 53064 17144
rect 53196 17138 53248 17144
rect 52932 16998 52960 17138
rect 52920 16992 52972 16998
rect 53024 16969 53052 17138
rect 53208 17066 53236 17138
rect 53196 17060 53248 17066
rect 53196 17002 53248 17008
rect 52920 16934 52972 16940
rect 53010 16960 53066 16969
rect 52932 15978 52960 16934
rect 53010 16895 53066 16904
rect 53300 16250 53328 18906
rect 53378 17504 53434 17513
rect 53378 17439 53434 17448
rect 53392 17270 53420 17439
rect 53472 17332 53524 17338
rect 53760 17320 53788 19790
rect 53852 18834 53880 19910
rect 54496 19854 54524 20742
rect 54588 20534 54616 21354
rect 54772 20806 54800 22066
rect 55324 21894 55352 22066
rect 55680 22092 55732 22098
rect 55680 22034 55732 22040
rect 55404 21956 55456 21962
rect 55404 21898 55456 21904
rect 55312 21888 55364 21894
rect 55416 21865 55444 21898
rect 55312 21830 55364 21836
rect 55402 21856 55458 21865
rect 55036 21684 55088 21690
rect 55036 21626 55088 21632
rect 55048 21554 55076 21626
rect 55128 21616 55180 21622
rect 55128 21558 55180 21564
rect 54944 21548 54996 21554
rect 54944 21490 54996 21496
rect 55036 21548 55088 21554
rect 55036 21490 55088 21496
rect 54956 21321 54984 21490
rect 54942 21312 54998 21321
rect 54942 21247 54998 21256
rect 54956 21010 54984 21247
rect 54944 21004 54996 21010
rect 54944 20946 54996 20952
rect 55140 20874 55168 21558
rect 55324 21350 55352 21830
rect 55402 21791 55458 21800
rect 55588 21548 55640 21554
rect 55588 21490 55640 21496
rect 55312 21344 55364 21350
rect 55312 21286 55364 21292
rect 55128 20868 55180 20874
rect 55128 20810 55180 20816
rect 54760 20800 54812 20806
rect 54760 20742 54812 20748
rect 54576 20528 54628 20534
rect 54576 20470 54628 20476
rect 54588 19961 54616 20470
rect 54944 20460 54996 20466
rect 54944 20402 54996 20408
rect 54852 20392 54904 20398
rect 54852 20334 54904 20340
rect 54574 19952 54630 19961
rect 54574 19887 54630 19896
rect 54588 19854 54616 19887
rect 54484 19848 54536 19854
rect 54484 19790 54536 19796
rect 54576 19848 54628 19854
rect 54576 19790 54628 19796
rect 54864 19786 54892 20334
rect 54956 19854 54984 20402
rect 55324 20330 55352 21286
rect 55600 20806 55628 21490
rect 55692 21350 55720 22034
rect 55876 21690 55904 22510
rect 56152 22030 56180 22578
rect 56140 22024 56192 22030
rect 56140 21966 56192 21972
rect 55864 21684 55916 21690
rect 55864 21626 55916 21632
rect 55680 21344 55732 21350
rect 55680 21286 55732 21292
rect 55588 20800 55640 20806
rect 55588 20742 55640 20748
rect 55404 20460 55456 20466
rect 55404 20402 55456 20408
rect 55312 20324 55364 20330
rect 55312 20266 55364 20272
rect 55220 20256 55272 20262
rect 55220 20198 55272 20204
rect 54944 19848 54996 19854
rect 54944 19790 54996 19796
rect 54852 19780 54904 19786
rect 54852 19722 54904 19728
rect 54864 19496 54892 19722
rect 54944 19508 54996 19514
rect 54864 19468 54944 19496
rect 54944 19450 54996 19456
rect 53932 19440 53984 19446
rect 53932 19382 53984 19388
rect 54116 19440 54168 19446
rect 54116 19382 54168 19388
rect 53840 18828 53892 18834
rect 53840 18770 53892 18776
rect 53852 18154 53880 18770
rect 53840 18148 53892 18154
rect 53840 18090 53892 18096
rect 53944 17746 53972 19382
rect 54128 18970 54156 19382
rect 54116 18964 54168 18970
rect 54116 18906 54168 18912
rect 54208 18216 54260 18222
rect 54208 18158 54260 18164
rect 53932 17740 53984 17746
rect 53932 17682 53984 17688
rect 53840 17672 53892 17678
rect 53840 17614 53892 17620
rect 53472 17274 53524 17280
rect 53576 17292 53788 17320
rect 53380 17264 53432 17270
rect 53380 17206 53432 17212
rect 53484 16998 53512 17274
rect 53576 17066 53604 17292
rect 53746 17232 53802 17241
rect 53746 17167 53748 17176
rect 53800 17167 53802 17176
rect 53748 17138 53800 17144
rect 53564 17060 53616 17066
rect 53564 17002 53616 17008
rect 53472 16992 53524 16998
rect 53472 16934 53524 16940
rect 53576 16726 53604 17002
rect 53852 16794 53880 17614
rect 53944 17134 53972 17682
rect 54220 17542 54248 18158
rect 54760 18148 54812 18154
rect 54760 18090 54812 18096
rect 54484 18080 54536 18086
rect 54484 18022 54536 18028
rect 54496 17814 54524 18022
rect 54484 17808 54536 17814
rect 54484 17750 54536 17756
rect 54496 17678 54524 17750
rect 54772 17746 54800 18090
rect 55232 17746 55260 20198
rect 55416 20058 55444 20402
rect 55588 20256 55640 20262
rect 55588 20198 55640 20204
rect 55404 20052 55456 20058
rect 55404 19994 55456 20000
rect 55600 19786 55628 20198
rect 55588 19780 55640 19786
rect 55588 19722 55640 19728
rect 54760 17740 54812 17746
rect 54760 17682 54812 17688
rect 55220 17740 55272 17746
rect 55220 17682 55272 17688
rect 54484 17672 54536 17678
rect 54484 17614 54536 17620
rect 54576 17672 54628 17678
rect 54576 17614 54628 17620
rect 54208 17536 54260 17542
rect 54206 17504 54208 17513
rect 54392 17536 54444 17542
rect 54260 17504 54262 17513
rect 54392 17478 54444 17484
rect 54206 17439 54262 17448
rect 54404 17270 54432 17478
rect 54588 17338 54616 17614
rect 54576 17332 54628 17338
rect 54576 17274 54628 17280
rect 54392 17264 54444 17270
rect 54392 17206 54444 17212
rect 53932 17128 53984 17134
rect 53932 17070 53984 17076
rect 53840 16788 53892 16794
rect 53840 16730 53892 16736
rect 53564 16720 53616 16726
rect 53564 16662 53616 16668
rect 53852 16574 53880 16730
rect 53760 16546 53880 16574
rect 53288 16244 53340 16250
rect 53288 16186 53340 16192
rect 53380 16244 53432 16250
rect 53380 16186 53432 16192
rect 52920 15972 52972 15978
rect 52920 15914 52972 15920
rect 52828 15904 52880 15910
rect 52828 15846 52880 15852
rect 52840 15502 52868 15846
rect 52828 15496 52880 15502
rect 52828 15438 52880 15444
rect 52736 15360 52788 15366
rect 52736 15302 52788 15308
rect 52552 14952 52604 14958
rect 52552 14894 52604 14900
rect 52564 14278 52592 14894
rect 52552 14272 52604 14278
rect 52552 14214 52604 14220
rect 52368 14000 52420 14006
rect 52368 13942 52420 13948
rect 52748 13734 52776 15302
rect 52840 15065 52868 15438
rect 52932 15434 52960 15914
rect 53392 15722 53420 16186
rect 53760 15910 53788 16546
rect 53944 16522 53972 17070
rect 54116 16584 54168 16590
rect 54116 16526 54168 16532
rect 53932 16516 53984 16522
rect 53932 16458 53984 16464
rect 53944 16046 53972 16458
rect 54128 16454 54156 16526
rect 54116 16448 54168 16454
rect 54116 16390 54168 16396
rect 53932 16040 53984 16046
rect 53932 15982 53984 15988
rect 53748 15904 53800 15910
rect 53748 15846 53800 15852
rect 53300 15694 53420 15722
rect 53300 15638 53328 15694
rect 53288 15632 53340 15638
rect 53288 15574 53340 15580
rect 53196 15496 53248 15502
rect 53564 15496 53616 15502
rect 53196 15438 53248 15444
rect 53562 15464 53564 15473
rect 53616 15464 53618 15473
rect 52920 15428 52972 15434
rect 52920 15370 52972 15376
rect 53208 15337 53236 15438
rect 53288 15428 53340 15434
rect 53562 15399 53618 15408
rect 53288 15370 53340 15376
rect 53194 15328 53250 15337
rect 53194 15263 53250 15272
rect 53300 15094 53328 15370
rect 53760 15094 53788 15846
rect 53840 15360 53892 15366
rect 53840 15302 53892 15308
rect 53288 15088 53340 15094
rect 52826 15056 52882 15065
rect 53288 15030 53340 15036
rect 53748 15088 53800 15094
rect 53748 15030 53800 15036
rect 52826 14991 52882 15000
rect 53760 14958 53788 15030
rect 53012 14952 53064 14958
rect 53012 14894 53064 14900
rect 53748 14952 53800 14958
rect 53748 14894 53800 14900
rect 53024 14482 53052 14894
rect 53012 14476 53064 14482
rect 53012 14418 53064 14424
rect 53760 14346 53788 14894
rect 53748 14340 53800 14346
rect 53748 14282 53800 14288
rect 53852 14090 53880 15302
rect 53944 15162 53972 15982
rect 54128 15570 54156 16390
rect 54772 16250 54800 17682
rect 54852 17264 54904 17270
rect 54852 17206 54904 17212
rect 54864 16794 54892 17206
rect 54852 16788 54904 16794
rect 54852 16730 54904 16736
rect 54760 16244 54812 16250
rect 54760 16186 54812 16192
rect 54758 16144 54814 16153
rect 54758 16079 54760 16088
rect 54812 16079 54814 16088
rect 54944 16108 54996 16114
rect 54760 16050 54812 16056
rect 54944 16050 54996 16056
rect 54760 15700 54812 15706
rect 54760 15642 54812 15648
rect 54116 15564 54168 15570
rect 54116 15506 54168 15512
rect 53932 15156 53984 15162
rect 53932 15098 53984 15104
rect 54772 14958 54800 15642
rect 54760 14952 54812 14958
rect 54760 14894 54812 14900
rect 53760 14074 53880 14090
rect 53748 14068 53880 14074
rect 53800 14062 53880 14068
rect 53748 14010 53800 14016
rect 52276 13728 52328 13734
rect 52276 13670 52328 13676
rect 52736 13728 52788 13734
rect 52736 13670 52788 13676
rect 51908 13524 51960 13530
rect 51908 13466 51960 13472
rect 52000 13524 52052 13530
rect 52000 13466 52052 13472
rect 51724 13456 51776 13462
rect 51724 13398 51776 13404
rect 51448 13388 51500 13394
rect 51448 13330 51500 13336
rect 52288 13190 52316 13670
rect 54956 13530 54984 16050
rect 55232 15366 55260 17682
rect 55692 17542 55720 21286
rect 56152 21010 56180 21966
rect 56612 21468 56640 22918
rect 56692 21616 56744 21622
rect 56690 21584 56692 21593
rect 56744 21584 56746 21593
rect 56690 21519 56746 21528
rect 56692 21480 56744 21486
rect 56612 21440 56692 21468
rect 56692 21422 56744 21428
rect 56140 21004 56192 21010
rect 56140 20946 56192 20952
rect 55956 20868 56008 20874
rect 55956 20810 56008 20816
rect 55968 20398 55996 20810
rect 56048 20800 56100 20806
rect 56048 20742 56100 20748
rect 55956 20392 56008 20398
rect 55956 20334 56008 20340
rect 55968 20058 55996 20334
rect 56060 20262 56088 20742
rect 56048 20256 56100 20262
rect 56048 20198 56100 20204
rect 55956 20052 56008 20058
rect 55956 19994 56008 20000
rect 55956 19712 56008 19718
rect 55956 19654 56008 19660
rect 55968 17814 55996 19654
rect 56060 18086 56088 20198
rect 56152 19922 56180 20946
rect 56704 20942 56732 21422
rect 56692 20936 56744 20942
rect 56692 20878 56744 20884
rect 56232 20800 56284 20806
rect 56232 20742 56284 20748
rect 56324 20800 56376 20806
rect 56324 20742 56376 20748
rect 56244 20482 56272 20742
rect 56336 20602 56364 20742
rect 56324 20596 56376 20602
rect 56324 20538 56376 20544
rect 56244 20466 56364 20482
rect 56244 20460 56376 20466
rect 56244 20454 56324 20460
rect 56324 20402 56376 20408
rect 56140 19916 56192 19922
rect 56140 19858 56192 19864
rect 56704 19854 56732 20878
rect 56692 19848 56744 19854
rect 56692 19790 56744 19796
rect 56796 19514 56824 24908
rect 57704 24608 57756 24614
rect 57704 24550 57756 24556
rect 57716 24342 57744 24550
rect 57704 24336 57756 24342
rect 57704 24278 57756 24284
rect 57428 24200 57480 24206
rect 57428 24142 57480 24148
rect 57440 23662 57468 24142
rect 58256 24064 58308 24070
rect 58256 24006 58308 24012
rect 58268 23730 58296 24006
rect 58256 23724 58308 23730
rect 58256 23666 58308 23672
rect 57428 23656 57480 23662
rect 57428 23598 57480 23604
rect 57440 23322 57468 23598
rect 58440 23520 58492 23526
rect 58440 23462 58492 23468
rect 57428 23316 57480 23322
rect 57428 23258 57480 23264
rect 58452 23225 58480 23462
rect 58438 23216 58494 23225
rect 58438 23151 58494 23160
rect 58256 22636 58308 22642
rect 58256 22578 58308 22584
rect 57520 21956 57572 21962
rect 57520 21898 57572 21904
rect 57532 21690 57560 21898
rect 58268 21894 58296 22578
rect 58438 22536 58494 22545
rect 58438 22471 58440 22480
rect 58492 22471 58494 22480
rect 58440 22442 58492 22448
rect 58256 21888 58308 21894
rect 58256 21830 58308 21836
rect 58440 21888 58492 21894
rect 58440 21830 58492 21836
rect 57520 21684 57572 21690
rect 57520 21626 57572 21632
rect 56968 21616 57020 21622
rect 56968 21558 57020 21564
rect 56876 21548 56928 21554
rect 56876 21490 56928 21496
rect 56888 20505 56916 21490
rect 56874 20496 56930 20505
rect 56874 20431 56930 20440
rect 56784 19508 56836 19514
rect 56784 19450 56836 19456
rect 56600 19372 56652 19378
rect 56600 19314 56652 19320
rect 56048 18080 56100 18086
rect 56048 18022 56100 18028
rect 56416 18080 56468 18086
rect 56416 18022 56468 18028
rect 55956 17808 56008 17814
rect 55956 17750 56008 17756
rect 55772 17604 55824 17610
rect 55772 17546 55824 17552
rect 55680 17536 55732 17542
rect 55680 17478 55732 17484
rect 55312 16652 55364 16658
rect 55312 16594 55364 16600
rect 55324 16522 55352 16594
rect 55312 16516 55364 16522
rect 55312 16458 55364 16464
rect 55324 16182 55352 16458
rect 55312 16176 55364 16182
rect 55312 16118 55364 16124
rect 55692 16114 55720 17478
rect 55784 17338 55812 17546
rect 55772 17332 55824 17338
rect 55772 17274 55824 17280
rect 55784 16658 55812 17274
rect 55772 16652 55824 16658
rect 55772 16594 55824 16600
rect 55968 16522 55996 17750
rect 56428 17678 56456 18022
rect 56612 17882 56640 19314
rect 56876 18760 56928 18766
rect 56876 18702 56928 18708
rect 56784 18284 56836 18290
rect 56784 18226 56836 18232
rect 56600 17876 56652 17882
rect 56600 17818 56652 17824
rect 56416 17672 56468 17678
rect 56416 17614 56468 17620
rect 56600 17672 56652 17678
rect 56796 17649 56824 18226
rect 56888 17678 56916 18702
rect 56980 18426 57008 21558
rect 58452 21554 58480 21830
rect 58440 21548 58492 21554
rect 58440 21490 58492 21496
rect 57796 20868 57848 20874
rect 57796 20810 57848 20816
rect 57808 20602 57836 20810
rect 57796 20596 57848 20602
rect 57796 20538 57848 20544
rect 58164 19848 58216 19854
rect 58164 19790 58216 19796
rect 58256 19848 58308 19854
rect 58256 19790 58308 19796
rect 58438 19816 58494 19825
rect 57888 19712 57940 19718
rect 57888 19654 57940 19660
rect 57060 19236 57112 19242
rect 57060 19178 57112 19184
rect 56968 18420 57020 18426
rect 56968 18362 57020 18368
rect 56968 18284 57020 18290
rect 57072 18272 57100 19178
rect 57428 19168 57480 19174
rect 57900 19145 57928 19654
rect 57428 19110 57480 19116
rect 57886 19136 57942 19145
rect 57440 18766 57468 19110
rect 57886 19071 57942 19080
rect 57428 18760 57480 18766
rect 57428 18702 57480 18708
rect 58176 18290 58204 19790
rect 58268 19310 58296 19790
rect 58438 19751 58494 19760
rect 58452 19718 58480 19751
rect 58440 19712 58492 19718
rect 58440 19654 58492 19660
rect 58256 19304 58308 19310
rect 58256 19246 58308 19252
rect 58268 18970 58296 19246
rect 58256 18964 58308 18970
rect 58256 18906 58308 18912
rect 57020 18244 57100 18272
rect 58164 18284 58216 18290
rect 56968 18226 57020 18232
rect 58164 18226 58216 18232
rect 56876 17672 56928 17678
rect 56600 17614 56652 17620
rect 56782 17640 56838 17649
rect 56232 17536 56284 17542
rect 56232 17478 56284 17484
rect 56244 17270 56272 17478
rect 56232 17264 56284 17270
rect 56232 17206 56284 17212
rect 56612 16794 56640 17614
rect 56692 17604 56744 17610
rect 56876 17614 56928 17620
rect 56782 17575 56838 17584
rect 56692 17546 56744 17552
rect 56704 17241 56732 17546
rect 56888 17338 56916 17614
rect 56876 17332 56928 17338
rect 56876 17274 56928 17280
rect 56784 17264 56836 17270
rect 56690 17232 56746 17241
rect 56980 17218 57008 18226
rect 57428 18080 57480 18086
rect 57428 18022 57480 18028
rect 57440 17678 57468 18022
rect 58176 17882 58204 18226
rect 58164 17876 58216 17882
rect 58164 17818 58216 17824
rect 57428 17672 57480 17678
rect 57428 17614 57480 17620
rect 56836 17212 57008 17218
rect 56784 17206 57008 17212
rect 56690 17167 56746 17176
rect 56796 17190 57008 17206
rect 56704 17134 56732 17167
rect 56692 17128 56744 17134
rect 56692 17070 56744 17076
rect 56600 16788 56652 16794
rect 56600 16730 56652 16736
rect 55956 16516 56008 16522
rect 55956 16458 56008 16464
rect 56796 16266 56824 17190
rect 57520 17128 57572 17134
rect 57520 17070 57572 17076
rect 57532 16590 57560 17070
rect 57520 16584 57572 16590
rect 57520 16526 57572 16532
rect 57244 16516 57296 16522
rect 57244 16458 57296 16464
rect 57336 16516 57388 16522
rect 57336 16458 57388 16464
rect 56968 16448 57020 16454
rect 56968 16390 57020 16396
rect 56048 16244 56100 16250
rect 56048 16186 56100 16192
rect 56704 16238 56824 16266
rect 55680 16108 55732 16114
rect 55680 16050 55732 16056
rect 55404 15972 55456 15978
rect 55404 15914 55456 15920
rect 55416 15434 55444 15914
rect 55956 15904 56008 15910
rect 55956 15846 56008 15852
rect 55968 15502 55996 15846
rect 56060 15570 56088 16186
rect 56704 16182 56732 16238
rect 56692 16176 56744 16182
rect 56692 16118 56744 16124
rect 56600 16040 56652 16046
rect 56600 15982 56652 15988
rect 56612 15706 56640 15982
rect 56232 15700 56284 15706
rect 56232 15642 56284 15648
rect 56600 15700 56652 15706
rect 56600 15642 56652 15648
rect 56048 15564 56100 15570
rect 56048 15506 56100 15512
rect 56244 15502 56272 15642
rect 55680 15496 55732 15502
rect 55680 15438 55732 15444
rect 55956 15496 56008 15502
rect 55956 15438 56008 15444
rect 56232 15496 56284 15502
rect 56324 15496 56376 15502
rect 56232 15438 56284 15444
rect 56322 15464 56324 15473
rect 56376 15464 56378 15473
rect 55404 15428 55456 15434
rect 55404 15370 55456 15376
rect 55220 15360 55272 15366
rect 55692 15337 55720 15438
rect 55220 15302 55272 15308
rect 55678 15328 55734 15337
rect 55678 15263 55734 15272
rect 55128 15156 55180 15162
rect 55128 15098 55180 15104
rect 55034 15056 55090 15065
rect 55034 14991 55090 15000
rect 55048 14958 55076 14991
rect 55036 14952 55088 14958
rect 55036 14894 55088 14900
rect 54944 13524 54996 13530
rect 54944 13466 54996 13472
rect 55140 13394 55168 15098
rect 55128 13388 55180 13394
rect 55128 13330 55180 13336
rect 55692 13258 55720 15263
rect 55968 14958 55996 15438
rect 56322 15399 56378 15408
rect 56508 15360 56560 15366
rect 56508 15302 56560 15308
rect 56520 15094 56548 15302
rect 56508 15088 56560 15094
rect 56508 15030 56560 15036
rect 55956 14952 56008 14958
rect 55956 14894 56008 14900
rect 56704 14822 56732 16118
rect 56980 15502 57008 16390
rect 57256 15910 57284 16458
rect 57244 15904 57296 15910
rect 57244 15846 57296 15852
rect 57348 15638 57376 16458
rect 57704 15904 57756 15910
rect 57704 15846 57756 15852
rect 57336 15632 57388 15638
rect 57336 15574 57388 15580
rect 57716 15502 57744 15846
rect 56968 15496 57020 15502
rect 56968 15438 57020 15444
rect 57704 15496 57756 15502
rect 57704 15438 57756 15444
rect 56692 14816 56744 14822
rect 56692 14758 56744 14764
rect 55680 13252 55732 13258
rect 56704 13240 56732 14758
rect 57612 13932 57664 13938
rect 57612 13874 57664 13880
rect 56784 13252 56836 13258
rect 56704 13212 56784 13240
rect 55680 13194 55732 13200
rect 56784 13194 56836 13200
rect 52276 13184 52328 13190
rect 52276 13126 52328 13132
rect 57428 13184 57480 13190
rect 57428 13126 57480 13132
rect 50528 12980 50580 12986
rect 50528 12922 50580 12928
rect 57440 12850 57468 13126
rect 57624 12986 57652 13874
rect 58440 13728 58492 13734
rect 58438 13696 58440 13705
rect 58492 13696 58494 13705
rect 58438 13631 58494 13640
rect 57612 12980 57664 12986
rect 57612 12922 57664 12928
rect 50160 12844 50212 12850
rect 50160 12786 50212 12792
rect 57428 12844 57480 12850
rect 57428 12786 57480 12792
rect 48136 12776 48188 12782
rect 48136 12718 48188 12724
rect 46204 12436 46256 12442
rect 46204 12378 46256 12384
rect 46756 12436 46808 12442
rect 46756 12378 46808 12384
rect 45928 12300 45980 12306
rect 45928 12242 45980 12248
rect 46216 12238 46244 12378
rect 46204 12232 46256 12238
rect 46204 12174 46256 12180
rect 44272 11892 44324 11898
rect 44272 11834 44324 11840
rect 42800 11824 42852 11830
rect 42800 11766 42852 11772
rect 41696 11076 41748 11082
rect 41696 11018 41748 11024
rect 41512 9988 41564 9994
rect 41512 9930 41564 9936
rect 41236 9580 41288 9586
rect 41236 9522 41288 9528
rect 41524 8634 41552 9930
rect 41512 8628 41564 8634
rect 41512 8570 41564 8576
rect 40316 8084 40368 8090
rect 40316 8026 40368 8032
rect 41052 8084 41104 8090
rect 41052 8026 41104 8032
rect 38016 7880 38068 7886
rect 38016 7822 38068 7828
rect 40040 7880 40092 7886
rect 40040 7822 40092 7828
rect 38028 7546 38056 7822
rect 38752 7744 38804 7750
rect 38752 7686 38804 7692
rect 38016 7540 38068 7546
rect 38016 7482 38068 7488
rect 37924 7472 37976 7478
rect 37924 7414 37976 7420
rect 37648 7336 37700 7342
rect 37648 7278 37700 7284
rect 37372 5908 37424 5914
rect 37372 5850 37424 5856
rect 37384 5370 37412 5850
rect 37936 5658 37964 7414
rect 38764 7410 38792 7686
rect 40052 7410 40080 7822
rect 38752 7404 38804 7410
rect 38752 7346 38804 7352
rect 40040 7404 40092 7410
rect 40040 7346 40092 7352
rect 37844 5642 37964 5658
rect 37832 5636 37964 5642
rect 37884 5630 37964 5636
rect 37832 5578 37884 5584
rect 37372 5364 37424 5370
rect 37372 5306 37424 5312
rect 37096 5228 37148 5234
rect 37096 5170 37148 5176
rect 34152 4820 34204 4826
rect 34152 4762 34204 4768
rect 34612 4820 34664 4826
rect 34612 4762 34664 4768
rect 34796 4820 34848 4826
rect 34796 4762 34848 4768
rect 36176 4820 36228 4826
rect 36176 4762 36228 4768
rect 34624 4554 34652 4762
rect 34612 4548 34664 4554
rect 34612 4490 34664 4496
rect 35594 4380 35902 4389
rect 35594 4378 35600 4380
rect 35656 4378 35680 4380
rect 35736 4378 35760 4380
rect 35816 4378 35840 4380
rect 35896 4378 35902 4380
rect 35656 4326 35658 4378
rect 35838 4326 35840 4378
rect 35594 4324 35600 4326
rect 35656 4324 35680 4326
rect 35736 4324 35760 4326
rect 35816 4324 35840 4326
rect 35896 4324 35902 4326
rect 35594 4315 35902 4324
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 35594 3292 35902 3301
rect 35594 3290 35600 3292
rect 35656 3290 35680 3292
rect 35736 3290 35760 3292
rect 35816 3290 35840 3292
rect 35896 3290 35902 3292
rect 35656 3238 35658 3290
rect 35838 3238 35840 3290
rect 35594 3236 35600 3238
rect 35656 3236 35680 3238
rect 35736 3236 35760 3238
rect 35816 3236 35840 3238
rect 35896 3236 35902 3238
rect 35594 3227 35902 3236
rect 33784 3188 33836 3194
rect 33784 3130 33836 3136
rect 32312 3120 32364 3126
rect 32312 3062 32364 3068
rect 32404 3120 32456 3126
rect 32404 3062 32456 3068
rect 32864 3120 32916 3126
rect 32864 3062 32916 3068
rect 35348 3052 35400 3058
rect 35348 2994 35400 3000
rect 37280 3052 37332 3058
rect 37280 2994 37332 3000
rect 42432 3052 42484 3058
rect 42432 2994 42484 3000
rect 43628 3052 43680 3058
rect 43628 2994 43680 3000
rect 31484 2984 31536 2990
rect 31484 2926 31536 2932
rect 34152 2848 34204 2854
rect 34152 2790 34204 2796
rect 34796 2848 34848 2854
rect 34796 2790 34848 2796
rect 30104 2440 30156 2446
rect 30104 2382 30156 2388
rect 30288 2440 30340 2446
rect 30288 2382 30340 2388
rect 30748 2440 30800 2446
rect 30748 2382 30800 2388
rect 29644 2372 29696 2378
rect 29644 2314 29696 2320
rect 29656 800 29684 2314
rect 30288 2304 30340 2310
rect 30288 2246 30340 2252
rect 30932 2304 30984 2310
rect 30932 2246 30984 2252
rect 30300 800 30328 2246
rect 30944 800 30972 2246
rect 34164 800 34192 2790
rect 34808 800 34836 2790
rect 34934 2748 35242 2757
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 35360 2514 35388 2994
rect 35440 2848 35492 2854
rect 35440 2790 35492 2796
rect 36084 2848 36136 2854
rect 36084 2790 36136 2796
rect 36728 2848 36780 2854
rect 36728 2790 36780 2796
rect 35348 2508 35400 2514
rect 35348 2450 35400 2456
rect 35452 800 35480 2790
rect 35594 2204 35902 2213
rect 35594 2202 35600 2204
rect 35656 2202 35680 2204
rect 35736 2202 35760 2204
rect 35816 2202 35840 2204
rect 35896 2202 35902 2204
rect 35656 2150 35658 2202
rect 35838 2150 35840 2202
rect 35594 2148 35600 2150
rect 35656 2148 35680 2150
rect 35736 2148 35760 2150
rect 35816 2148 35840 2150
rect 35896 2148 35902 2150
rect 35594 2139 35902 2148
rect 36096 800 36124 2790
rect 36740 800 36768 2790
rect 37292 2514 37320 2994
rect 37372 2848 37424 2854
rect 37372 2790 37424 2796
rect 38016 2848 38068 2854
rect 38016 2790 38068 2796
rect 38660 2848 38712 2854
rect 38660 2790 38712 2796
rect 39304 2848 39356 2854
rect 39304 2790 39356 2796
rect 39948 2848 40000 2854
rect 39948 2790 40000 2796
rect 40592 2848 40644 2854
rect 40592 2790 40644 2796
rect 41236 2848 41288 2854
rect 41236 2790 41288 2796
rect 41880 2848 41932 2854
rect 41880 2790 41932 2796
rect 37280 2508 37332 2514
rect 37280 2450 37332 2456
rect 37384 800 37412 2790
rect 38028 800 38056 2790
rect 38672 800 38700 2790
rect 39316 800 39344 2790
rect 39960 800 39988 2790
rect 40604 800 40632 2790
rect 41248 800 41276 2790
rect 41892 800 41920 2790
rect 42444 2514 42472 2994
rect 42524 2848 42576 2854
rect 42524 2790 42576 2796
rect 43168 2848 43220 2854
rect 43168 2790 43220 2796
rect 42432 2508 42484 2514
rect 42432 2450 42484 2456
rect 42536 800 42564 2790
rect 43180 800 43208 2790
rect 43640 2514 43668 2994
rect 43812 2848 43864 2854
rect 43812 2790 43864 2796
rect 44456 2848 44508 2854
rect 44456 2790 44508 2796
rect 45100 2848 45152 2854
rect 45100 2790 45152 2796
rect 43628 2508 43680 2514
rect 43628 2450 43680 2456
rect 43824 800 43852 2790
rect 44468 800 44496 2790
rect 45112 800 45140 2790
rect 18 0 74 800
rect 662 0 718 800
rect 1306 0 1362 800
rect 1950 0 2006 800
rect 2594 0 2650 800
rect 3238 0 3294 800
rect 3882 0 3938 800
rect 4526 0 4582 800
rect 5170 0 5226 800
rect 5814 0 5870 800
rect 6458 0 6514 800
rect 7102 0 7158 800
rect 7746 0 7802 800
rect 8390 0 8446 800
rect 9034 0 9090 800
rect 9678 0 9734 800
rect 10322 0 10378 800
rect 10966 0 11022 800
rect 11610 0 11666 800
rect 12254 0 12310 800
rect 12898 0 12954 800
rect 13542 0 13598 800
rect 14186 0 14242 800
rect 14830 0 14886 800
rect 15474 0 15530 800
rect 16118 0 16174 800
rect 16762 0 16818 800
rect 17406 0 17462 800
rect 18050 0 18106 800
rect 18694 0 18750 800
rect 19338 0 19394 800
rect 20626 0 20682 800
rect 21270 0 21326 800
rect 22558 0 22614 800
rect 23202 0 23258 800
rect 28998 0 29054 800
rect 29642 0 29698 800
rect 30286 0 30342 800
rect 30930 0 30986 800
rect 34150 0 34206 800
rect 34794 0 34850 800
rect 35438 0 35494 800
rect 36082 0 36138 800
rect 36726 0 36782 800
rect 37370 0 37426 800
rect 38014 0 38070 800
rect 38658 0 38714 800
rect 39302 0 39358 800
rect 39946 0 40002 800
rect 40590 0 40646 800
rect 41234 0 41290 800
rect 41878 0 41934 800
rect 42522 0 42578 800
rect 43166 0 43222 800
rect 43810 0 43866 800
rect 44454 0 44510 800
rect 45098 0 45154 800
<< via2 >>
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 4880 37018 4936 37020
rect 4960 37018 5016 37020
rect 5040 37018 5096 37020
rect 5120 37018 5176 37020
rect 4880 36966 4926 37018
rect 4926 36966 4936 37018
rect 4960 36966 4990 37018
rect 4990 36966 5002 37018
rect 5002 36966 5016 37018
rect 5040 36966 5054 37018
rect 5054 36966 5066 37018
rect 5066 36966 5096 37018
rect 5120 36966 5130 37018
rect 5130 36966 5176 37018
rect 4880 36964 4936 36966
rect 4960 36964 5016 36966
rect 5040 36964 5096 36966
rect 5120 36964 5176 36966
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4880 35930 4936 35932
rect 4960 35930 5016 35932
rect 5040 35930 5096 35932
rect 5120 35930 5176 35932
rect 4880 35878 4926 35930
rect 4926 35878 4936 35930
rect 4960 35878 4990 35930
rect 4990 35878 5002 35930
rect 5002 35878 5016 35930
rect 5040 35878 5054 35930
rect 5054 35878 5066 35930
rect 5066 35878 5096 35930
rect 5120 35878 5130 35930
rect 5130 35878 5176 35930
rect 4880 35876 4936 35878
rect 4960 35876 5016 35878
rect 5040 35876 5096 35878
rect 5120 35876 5176 35878
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4880 34842 4936 34844
rect 4960 34842 5016 34844
rect 5040 34842 5096 34844
rect 5120 34842 5176 34844
rect 4880 34790 4926 34842
rect 4926 34790 4936 34842
rect 4960 34790 4990 34842
rect 4990 34790 5002 34842
rect 5002 34790 5016 34842
rect 5040 34790 5054 34842
rect 5054 34790 5066 34842
rect 5066 34790 5096 34842
rect 5120 34790 5130 34842
rect 5130 34790 5176 34842
rect 4880 34788 4936 34790
rect 4960 34788 5016 34790
rect 5040 34788 5096 34790
rect 5120 34788 5176 34790
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4880 33754 4936 33756
rect 4960 33754 5016 33756
rect 5040 33754 5096 33756
rect 5120 33754 5176 33756
rect 4880 33702 4926 33754
rect 4926 33702 4936 33754
rect 4960 33702 4990 33754
rect 4990 33702 5002 33754
rect 5002 33702 5016 33754
rect 5040 33702 5054 33754
rect 5054 33702 5066 33754
rect 5066 33702 5096 33754
rect 5120 33702 5130 33754
rect 5130 33702 5176 33754
rect 4880 33700 4936 33702
rect 4960 33700 5016 33702
rect 5040 33700 5096 33702
rect 5120 33700 5176 33702
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4880 32666 4936 32668
rect 4960 32666 5016 32668
rect 5040 32666 5096 32668
rect 5120 32666 5176 32668
rect 4880 32614 4926 32666
rect 4926 32614 4936 32666
rect 4960 32614 4990 32666
rect 4990 32614 5002 32666
rect 5002 32614 5016 32666
rect 5040 32614 5054 32666
rect 5054 32614 5066 32666
rect 5066 32614 5096 32666
rect 5120 32614 5130 32666
rect 5130 32614 5176 32666
rect 4880 32612 4936 32614
rect 4960 32612 5016 32614
rect 5040 32612 5096 32614
rect 5120 32612 5176 32614
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4880 31578 4936 31580
rect 4960 31578 5016 31580
rect 5040 31578 5096 31580
rect 5120 31578 5176 31580
rect 4880 31526 4926 31578
rect 4926 31526 4936 31578
rect 4960 31526 4990 31578
rect 4990 31526 5002 31578
rect 5002 31526 5016 31578
rect 5040 31526 5054 31578
rect 5054 31526 5066 31578
rect 5066 31526 5096 31578
rect 5120 31526 5130 31578
rect 5130 31526 5176 31578
rect 4880 31524 4936 31526
rect 4960 31524 5016 31526
rect 5040 31524 5096 31526
rect 5120 31524 5176 31526
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4880 30490 4936 30492
rect 4960 30490 5016 30492
rect 5040 30490 5096 30492
rect 5120 30490 5176 30492
rect 4880 30438 4926 30490
rect 4926 30438 4936 30490
rect 4960 30438 4990 30490
rect 4990 30438 5002 30490
rect 5002 30438 5016 30490
rect 5040 30438 5054 30490
rect 5054 30438 5066 30490
rect 5066 30438 5096 30490
rect 5120 30438 5130 30490
rect 5130 30438 5176 30490
rect 4880 30436 4936 30438
rect 4960 30436 5016 30438
rect 5040 30436 5096 30438
rect 5120 30436 5176 30438
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4880 29402 4936 29404
rect 4960 29402 5016 29404
rect 5040 29402 5096 29404
rect 5120 29402 5176 29404
rect 4880 29350 4926 29402
rect 4926 29350 4936 29402
rect 4960 29350 4990 29402
rect 4990 29350 5002 29402
rect 5002 29350 5016 29402
rect 5040 29350 5054 29402
rect 5054 29350 5066 29402
rect 5066 29350 5096 29402
rect 5120 29350 5130 29402
rect 5130 29350 5176 29402
rect 4880 29348 4936 29350
rect 4960 29348 5016 29350
rect 5040 29348 5096 29350
rect 5120 29348 5176 29350
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4880 28314 4936 28316
rect 4960 28314 5016 28316
rect 5040 28314 5096 28316
rect 5120 28314 5176 28316
rect 4880 28262 4926 28314
rect 4926 28262 4936 28314
rect 4960 28262 4990 28314
rect 4990 28262 5002 28314
rect 5002 28262 5016 28314
rect 5040 28262 5054 28314
rect 5054 28262 5066 28314
rect 5066 28262 5096 28314
rect 5120 28262 5130 28314
rect 5130 28262 5176 28314
rect 4880 28260 4936 28262
rect 4960 28260 5016 28262
rect 5040 28260 5096 28262
rect 5120 28260 5176 28262
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4880 27226 4936 27228
rect 4960 27226 5016 27228
rect 5040 27226 5096 27228
rect 5120 27226 5176 27228
rect 4880 27174 4926 27226
rect 4926 27174 4936 27226
rect 4960 27174 4990 27226
rect 4990 27174 5002 27226
rect 5002 27174 5016 27226
rect 5040 27174 5054 27226
rect 5054 27174 5066 27226
rect 5066 27174 5096 27226
rect 5120 27174 5130 27226
rect 5130 27174 5176 27226
rect 4880 27172 4936 27174
rect 4960 27172 5016 27174
rect 5040 27172 5096 27174
rect 5120 27172 5176 27174
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4880 26138 4936 26140
rect 4960 26138 5016 26140
rect 5040 26138 5096 26140
rect 5120 26138 5176 26140
rect 4880 26086 4926 26138
rect 4926 26086 4936 26138
rect 4960 26086 4990 26138
rect 4990 26086 5002 26138
rect 5002 26086 5016 26138
rect 5040 26086 5054 26138
rect 5054 26086 5066 26138
rect 5066 26086 5096 26138
rect 5120 26086 5130 26138
rect 5130 26086 5176 26138
rect 4880 26084 4936 26086
rect 4960 26084 5016 26086
rect 5040 26084 5096 26086
rect 5120 26084 5176 26086
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4880 25050 4936 25052
rect 4960 25050 5016 25052
rect 5040 25050 5096 25052
rect 5120 25050 5176 25052
rect 4880 24998 4926 25050
rect 4926 24998 4936 25050
rect 4960 24998 4990 25050
rect 4990 24998 5002 25050
rect 5002 24998 5016 25050
rect 5040 24998 5054 25050
rect 5054 24998 5066 25050
rect 5066 24998 5096 25050
rect 5120 24998 5130 25050
rect 5130 24998 5176 25050
rect 4880 24996 4936 24998
rect 4960 24996 5016 24998
rect 5040 24996 5096 24998
rect 5120 24996 5176 24998
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4880 23962 4936 23964
rect 4960 23962 5016 23964
rect 5040 23962 5096 23964
rect 5120 23962 5176 23964
rect 4880 23910 4926 23962
rect 4926 23910 4936 23962
rect 4960 23910 4990 23962
rect 4990 23910 5002 23962
rect 5002 23910 5016 23962
rect 5040 23910 5054 23962
rect 5054 23910 5066 23962
rect 5066 23910 5096 23962
rect 5120 23910 5130 23962
rect 5130 23910 5176 23962
rect 4880 23908 4936 23910
rect 4960 23908 5016 23910
rect 5040 23908 5096 23910
rect 5120 23908 5176 23910
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4880 22874 4936 22876
rect 4960 22874 5016 22876
rect 5040 22874 5096 22876
rect 5120 22874 5176 22876
rect 4880 22822 4926 22874
rect 4926 22822 4936 22874
rect 4960 22822 4990 22874
rect 4990 22822 5002 22874
rect 5002 22822 5016 22874
rect 5040 22822 5054 22874
rect 5054 22822 5066 22874
rect 5066 22822 5096 22874
rect 5120 22822 5130 22874
rect 5130 22822 5176 22874
rect 4880 22820 4936 22822
rect 4960 22820 5016 22822
rect 5040 22820 5096 22822
rect 5120 22820 5176 22822
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4880 21786 4936 21788
rect 4960 21786 5016 21788
rect 5040 21786 5096 21788
rect 5120 21786 5176 21788
rect 4880 21734 4926 21786
rect 4926 21734 4936 21786
rect 4960 21734 4990 21786
rect 4990 21734 5002 21786
rect 5002 21734 5016 21786
rect 5040 21734 5054 21786
rect 5054 21734 5066 21786
rect 5066 21734 5096 21786
rect 5120 21734 5130 21786
rect 5130 21734 5176 21786
rect 4880 21732 4936 21734
rect 4960 21732 5016 21734
rect 5040 21732 5096 21734
rect 5120 21732 5176 21734
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4880 20698 4936 20700
rect 4960 20698 5016 20700
rect 5040 20698 5096 20700
rect 5120 20698 5176 20700
rect 4880 20646 4926 20698
rect 4926 20646 4936 20698
rect 4960 20646 4990 20698
rect 4990 20646 5002 20698
rect 5002 20646 5016 20698
rect 5040 20646 5054 20698
rect 5054 20646 5066 20698
rect 5066 20646 5096 20698
rect 5120 20646 5130 20698
rect 5130 20646 5176 20698
rect 4880 20644 4936 20646
rect 4960 20644 5016 20646
rect 5040 20644 5096 20646
rect 5120 20644 5176 20646
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 846 19660 848 19680
rect 848 19660 900 19680
rect 900 19660 902 19680
rect 846 19624 902 19660
rect 4880 19610 4936 19612
rect 4960 19610 5016 19612
rect 5040 19610 5096 19612
rect 5120 19610 5176 19612
rect 4880 19558 4926 19610
rect 4926 19558 4936 19610
rect 4960 19558 4990 19610
rect 4990 19558 5002 19610
rect 5002 19558 5016 19610
rect 5040 19558 5054 19610
rect 5054 19558 5066 19610
rect 5066 19558 5096 19610
rect 5120 19558 5130 19610
rect 5130 19558 5176 19610
rect 4880 19556 4936 19558
rect 4960 19556 5016 19558
rect 5040 19556 5096 19558
rect 5120 19556 5176 19558
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4880 18522 4936 18524
rect 4960 18522 5016 18524
rect 5040 18522 5096 18524
rect 5120 18522 5176 18524
rect 4880 18470 4926 18522
rect 4926 18470 4936 18522
rect 4960 18470 4990 18522
rect 4990 18470 5002 18522
rect 5002 18470 5016 18522
rect 5040 18470 5054 18522
rect 5054 18470 5066 18522
rect 5066 18470 5096 18522
rect 5120 18470 5130 18522
rect 5130 18470 5176 18522
rect 4880 18468 4936 18470
rect 4960 18468 5016 18470
rect 5040 18468 5096 18470
rect 5120 18468 5176 18470
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4880 17434 4936 17436
rect 4960 17434 5016 17436
rect 5040 17434 5096 17436
rect 5120 17434 5176 17436
rect 4880 17382 4926 17434
rect 4926 17382 4936 17434
rect 4960 17382 4990 17434
rect 4990 17382 5002 17434
rect 5002 17382 5016 17434
rect 5040 17382 5054 17434
rect 5054 17382 5066 17434
rect 5066 17382 5096 17434
rect 5120 17382 5130 17434
rect 5130 17382 5176 17434
rect 4880 17380 4936 17382
rect 4960 17380 5016 17382
rect 5040 17380 5096 17382
rect 5120 17380 5176 17382
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4880 16346 4936 16348
rect 4960 16346 5016 16348
rect 5040 16346 5096 16348
rect 5120 16346 5176 16348
rect 4880 16294 4926 16346
rect 4926 16294 4936 16346
rect 4960 16294 4990 16346
rect 4990 16294 5002 16346
rect 5002 16294 5016 16346
rect 5040 16294 5054 16346
rect 5054 16294 5066 16346
rect 5066 16294 5096 16346
rect 5120 16294 5130 16346
rect 5130 16294 5176 16346
rect 4880 16292 4936 16294
rect 4960 16292 5016 16294
rect 5040 16292 5096 16294
rect 5120 16292 5176 16294
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4880 15258 4936 15260
rect 4960 15258 5016 15260
rect 5040 15258 5096 15260
rect 5120 15258 5176 15260
rect 4880 15206 4926 15258
rect 4926 15206 4936 15258
rect 4960 15206 4990 15258
rect 4990 15206 5002 15258
rect 5002 15206 5016 15258
rect 5040 15206 5054 15258
rect 5054 15206 5066 15258
rect 5066 15206 5096 15258
rect 5120 15206 5130 15258
rect 5130 15206 5176 15258
rect 4880 15204 4936 15206
rect 4960 15204 5016 15206
rect 5040 15204 5096 15206
rect 5120 15204 5176 15206
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 1214 14356 1216 14376
rect 1216 14356 1268 14376
rect 1268 14356 1270 14376
rect 1214 14320 1270 14356
rect 4880 14170 4936 14172
rect 4960 14170 5016 14172
rect 5040 14170 5096 14172
rect 5120 14170 5176 14172
rect 4880 14118 4926 14170
rect 4926 14118 4936 14170
rect 4960 14118 4990 14170
rect 4990 14118 5002 14170
rect 5002 14118 5016 14170
rect 5040 14118 5054 14170
rect 5054 14118 5066 14170
rect 5066 14118 5096 14170
rect 5120 14118 5130 14170
rect 5130 14118 5176 14170
rect 4880 14116 4936 14118
rect 4960 14116 5016 14118
rect 5040 14116 5096 14118
rect 5120 14116 5176 14118
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4880 13082 4936 13084
rect 4960 13082 5016 13084
rect 5040 13082 5096 13084
rect 5120 13082 5176 13084
rect 4880 13030 4926 13082
rect 4926 13030 4936 13082
rect 4960 13030 4990 13082
rect 4990 13030 5002 13082
rect 5002 13030 5016 13082
rect 5040 13030 5054 13082
rect 5054 13030 5066 13082
rect 5066 13030 5096 13082
rect 5120 13030 5130 13082
rect 5130 13030 5176 13082
rect 4880 13028 4936 13030
rect 4960 13028 5016 13030
rect 5040 13028 5096 13030
rect 5120 13028 5176 13030
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4880 11994 4936 11996
rect 4960 11994 5016 11996
rect 5040 11994 5096 11996
rect 5120 11994 5176 11996
rect 4880 11942 4926 11994
rect 4926 11942 4936 11994
rect 4960 11942 4990 11994
rect 4990 11942 5002 11994
rect 5002 11942 5016 11994
rect 5040 11942 5054 11994
rect 5054 11942 5066 11994
rect 5066 11942 5096 11994
rect 5120 11942 5130 11994
rect 5130 11942 5176 11994
rect 4880 11940 4936 11942
rect 4960 11940 5016 11942
rect 5040 11940 5096 11942
rect 5120 11940 5176 11942
rect 19706 31456 19762 31512
rect 19430 25064 19486 25120
rect 19890 21972 19892 21992
rect 19892 21972 19944 21992
rect 19944 21972 19946 21992
rect 19890 21936 19946 21972
rect 19798 20460 19854 20496
rect 19798 20440 19800 20460
rect 19800 20440 19852 20460
rect 19852 20440 19854 20460
rect 21730 25200 21786 25256
rect 20994 23860 21050 23896
rect 20994 23840 20996 23860
rect 20996 23840 21048 23860
rect 21048 23840 21050 23860
rect 20074 22344 20130 22400
rect 20442 22480 20498 22536
rect 22374 24248 22430 24304
rect 19982 20712 20038 20768
rect 20442 21684 20498 21720
rect 20442 21664 20444 21684
rect 20444 21664 20496 21684
rect 20496 21664 20498 21684
rect 22098 23976 22154 24032
rect 22558 23840 22614 23896
rect 20994 20748 20996 20768
rect 20996 20748 21048 20768
rect 21048 20748 21050 20768
rect 20994 20712 21050 20748
rect 22558 20476 22560 20496
rect 22560 20476 22612 20496
rect 22612 20476 22614 20496
rect 22558 20440 22614 20476
rect 19798 18672 19854 18728
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4880 10906 4936 10908
rect 4960 10906 5016 10908
rect 5040 10906 5096 10908
rect 5120 10906 5176 10908
rect 4880 10854 4926 10906
rect 4926 10854 4936 10906
rect 4960 10854 4990 10906
rect 4990 10854 5002 10906
rect 5002 10854 5016 10906
rect 5040 10854 5054 10906
rect 5054 10854 5066 10906
rect 5066 10854 5096 10906
rect 5120 10854 5130 10906
rect 5130 10854 5176 10906
rect 4880 10852 4936 10854
rect 4960 10852 5016 10854
rect 5040 10852 5096 10854
rect 5120 10852 5176 10854
rect 23386 31456 23442 31512
rect 23018 25064 23074 25120
rect 23294 25236 23296 25256
rect 23296 25236 23348 25256
rect 23348 25236 23350 25256
rect 23294 25200 23350 25236
rect 22834 24520 22890 24576
rect 22926 24248 22982 24304
rect 23846 23976 23902 24032
rect 23202 20440 23258 20496
rect 23846 21664 23902 21720
rect 25042 26288 25098 26344
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 35600 37018 35656 37020
rect 35680 37018 35736 37020
rect 35760 37018 35816 37020
rect 35840 37018 35896 37020
rect 35600 36966 35646 37018
rect 35646 36966 35656 37018
rect 35680 36966 35710 37018
rect 35710 36966 35722 37018
rect 35722 36966 35736 37018
rect 35760 36966 35774 37018
rect 35774 36966 35786 37018
rect 35786 36966 35816 37018
rect 35840 36966 35850 37018
rect 35850 36966 35896 37018
rect 35600 36964 35656 36966
rect 35680 36964 35736 36966
rect 35760 36964 35816 36966
rect 35840 36964 35896 36966
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 28078 29028 28134 29064
rect 28078 29008 28080 29028
rect 28080 29008 28132 29028
rect 28132 29008 28134 29028
rect 25962 26324 25964 26344
rect 25964 26324 26016 26344
rect 26016 26324 26018 26344
rect 25962 26288 26018 26324
rect 25318 24812 25374 24848
rect 25318 24792 25320 24812
rect 25320 24792 25372 24812
rect 25372 24792 25374 24812
rect 20074 18844 20076 18864
rect 20076 18844 20128 18864
rect 20128 18844 20130 18864
rect 20074 18808 20130 18844
rect 20534 18284 20590 18320
rect 20534 18264 20536 18284
rect 20536 18264 20588 18284
rect 20588 18264 20590 18284
rect 20350 15020 20406 15056
rect 22926 18808 22982 18864
rect 22466 18284 22522 18320
rect 22466 18264 22468 18284
rect 22468 18264 22520 18284
rect 22520 18264 22522 18284
rect 20350 15000 20352 15020
rect 20352 15000 20404 15020
rect 20404 15000 20406 15020
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4880 9818 4936 9820
rect 4960 9818 5016 9820
rect 5040 9818 5096 9820
rect 5120 9818 5176 9820
rect 4880 9766 4926 9818
rect 4926 9766 4936 9818
rect 4960 9766 4990 9818
rect 4990 9766 5002 9818
rect 5002 9766 5016 9818
rect 5040 9766 5054 9818
rect 5054 9766 5066 9818
rect 5066 9766 5096 9818
rect 5120 9766 5130 9818
rect 5130 9766 5176 9818
rect 4880 9764 4936 9766
rect 4960 9764 5016 9766
rect 5040 9764 5096 9766
rect 5120 9764 5176 9766
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4880 8730 4936 8732
rect 4960 8730 5016 8732
rect 5040 8730 5096 8732
rect 5120 8730 5176 8732
rect 4880 8678 4926 8730
rect 4926 8678 4936 8730
rect 4960 8678 4990 8730
rect 4990 8678 5002 8730
rect 5002 8678 5016 8730
rect 5040 8678 5054 8730
rect 5054 8678 5066 8730
rect 5066 8678 5096 8730
rect 5120 8678 5130 8730
rect 5130 8678 5176 8730
rect 4880 8676 4936 8678
rect 4960 8676 5016 8678
rect 5040 8676 5096 8678
rect 5120 8676 5176 8678
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4880 7642 4936 7644
rect 4960 7642 5016 7644
rect 5040 7642 5096 7644
rect 5120 7642 5176 7644
rect 4880 7590 4926 7642
rect 4926 7590 4936 7642
rect 4960 7590 4990 7642
rect 4990 7590 5002 7642
rect 5002 7590 5016 7642
rect 5040 7590 5054 7642
rect 5054 7590 5066 7642
rect 5066 7590 5096 7642
rect 5120 7590 5130 7642
rect 5130 7590 5176 7642
rect 4880 7588 4936 7590
rect 4960 7588 5016 7590
rect 5040 7588 5096 7590
rect 5120 7588 5176 7590
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4880 6554 4936 6556
rect 4960 6554 5016 6556
rect 5040 6554 5096 6556
rect 5120 6554 5176 6556
rect 4880 6502 4926 6554
rect 4926 6502 4936 6554
rect 4960 6502 4990 6554
rect 4990 6502 5002 6554
rect 5002 6502 5016 6554
rect 5040 6502 5054 6554
rect 5054 6502 5066 6554
rect 5066 6502 5096 6554
rect 5120 6502 5130 6554
rect 5130 6502 5176 6554
rect 4880 6500 4936 6502
rect 4960 6500 5016 6502
rect 5040 6500 5096 6502
rect 5120 6500 5176 6502
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4880 5466 4936 5468
rect 4960 5466 5016 5468
rect 5040 5466 5096 5468
rect 5120 5466 5176 5468
rect 4880 5414 4926 5466
rect 4926 5414 4936 5466
rect 4960 5414 4990 5466
rect 4990 5414 5002 5466
rect 5002 5414 5016 5466
rect 5040 5414 5054 5466
rect 5054 5414 5066 5466
rect 5066 5414 5096 5466
rect 5120 5414 5130 5466
rect 5130 5414 5176 5466
rect 4880 5412 4936 5414
rect 4960 5412 5016 5414
rect 5040 5412 5096 5414
rect 5120 5412 5176 5414
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4880 4378 4936 4380
rect 4960 4378 5016 4380
rect 5040 4378 5096 4380
rect 5120 4378 5176 4380
rect 4880 4326 4926 4378
rect 4926 4326 4936 4378
rect 4960 4326 4990 4378
rect 4990 4326 5002 4378
rect 5002 4326 5016 4378
rect 5040 4326 5054 4378
rect 5054 4326 5066 4378
rect 5066 4326 5096 4378
rect 5120 4326 5130 4378
rect 5130 4326 5176 4378
rect 4880 4324 4936 4326
rect 4960 4324 5016 4326
rect 5040 4324 5096 4326
rect 5120 4324 5176 4326
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4880 3290 4936 3292
rect 4960 3290 5016 3292
rect 5040 3290 5096 3292
rect 5120 3290 5176 3292
rect 4880 3238 4926 3290
rect 4926 3238 4936 3290
rect 4960 3238 4990 3290
rect 4990 3238 5002 3290
rect 5002 3238 5016 3290
rect 5040 3238 5054 3290
rect 5054 3238 5066 3290
rect 5066 3238 5096 3290
rect 5120 3238 5130 3290
rect 5130 3238 5176 3290
rect 4880 3236 4936 3238
rect 4960 3236 5016 3238
rect 5040 3236 5096 3238
rect 5120 3236 5176 3238
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 20258 13776 20314 13832
rect 22834 15020 22890 15056
rect 22834 15000 22836 15020
rect 22836 15000 22888 15020
rect 22888 15000 22890 15020
rect 24858 20712 24914 20768
rect 24582 19080 24638 19136
rect 24858 19080 24914 19136
rect 23294 15544 23350 15600
rect 24674 16904 24730 16960
rect 25778 24384 25834 24440
rect 25410 23976 25466 24032
rect 25134 18944 25190 19000
rect 25594 23840 25650 23896
rect 25410 18536 25466 18592
rect 25042 16632 25098 16688
rect 25042 16532 25044 16552
rect 25044 16532 25096 16552
rect 25096 16532 25098 16552
rect 25042 16496 25098 16532
rect 25318 16788 25374 16824
rect 25318 16768 25320 16788
rect 25320 16768 25372 16788
rect 25372 16768 25374 16788
rect 25870 23568 25926 23624
rect 27710 26324 27712 26344
rect 27712 26324 27764 26344
rect 27764 26324 27766 26344
rect 27710 26288 27766 26324
rect 26514 24404 26570 24440
rect 26514 24384 26516 24404
rect 26516 24384 26568 24404
rect 26568 24384 26570 24404
rect 26330 24248 26386 24304
rect 26330 24132 26386 24168
rect 26330 24112 26332 24132
rect 26332 24112 26384 24132
rect 26384 24112 26386 24132
rect 28446 26288 28502 26344
rect 25594 19216 25650 19272
rect 27066 23740 27068 23760
rect 27068 23740 27120 23760
rect 27120 23740 27122 23760
rect 27066 23704 27122 23740
rect 26146 20460 26202 20496
rect 26146 20440 26148 20460
rect 26148 20440 26200 20460
rect 26200 20440 26202 20460
rect 25870 19080 25926 19136
rect 26146 18672 26202 18728
rect 26514 19080 26570 19136
rect 26422 18808 26478 18864
rect 26606 18944 26662 19000
rect 26330 17076 26332 17096
rect 26332 17076 26384 17096
rect 26384 17076 26386 17096
rect 26330 17040 26386 17076
rect 26422 16652 26478 16688
rect 27526 24520 27582 24576
rect 27342 23160 27398 23216
rect 26790 18572 26792 18592
rect 26792 18572 26844 18592
rect 26844 18572 26846 18592
rect 26790 18536 26846 18572
rect 26974 19216 27030 19272
rect 26974 18964 27030 19000
rect 26974 18944 26976 18964
rect 26976 18944 27028 18964
rect 27028 18944 27030 18964
rect 26974 18672 27030 18728
rect 26422 16632 26424 16652
rect 26424 16632 26476 16652
rect 26476 16632 26478 16652
rect 27802 23568 27858 23624
rect 27434 21956 27490 21992
rect 27434 21936 27436 21956
rect 27436 21936 27488 21956
rect 27488 21936 27490 21956
rect 27250 18944 27306 19000
rect 27342 18808 27398 18864
rect 28446 24384 28502 24440
rect 28998 25200 29054 25256
rect 28814 24384 28870 24440
rect 27802 16904 27858 16960
rect 27710 15544 27766 15600
rect 27986 15544 28042 15600
rect 26238 12960 26294 13016
rect 27618 12980 27674 13016
rect 27618 12960 27620 12980
rect 27620 12960 27672 12980
rect 27672 12960 27674 12980
rect 26698 11056 26754 11112
rect 4880 2202 4936 2204
rect 4960 2202 5016 2204
rect 5040 2202 5096 2204
rect 5120 2202 5176 2204
rect 4880 2150 4926 2202
rect 4926 2150 4936 2202
rect 4960 2150 4990 2202
rect 4990 2150 5002 2202
rect 5002 2150 5016 2202
rect 5040 2150 5054 2202
rect 5054 2150 5066 2202
rect 5066 2150 5096 2202
rect 5120 2150 5130 2202
rect 5130 2150 5176 2202
rect 4880 2148 4936 2150
rect 4960 2148 5016 2150
rect 5040 2148 5096 2150
rect 5120 2148 5176 2150
rect 33046 32544 33102 32600
rect 35600 35930 35656 35932
rect 35680 35930 35736 35932
rect 35760 35930 35816 35932
rect 35840 35930 35896 35932
rect 35600 35878 35646 35930
rect 35646 35878 35656 35930
rect 35680 35878 35710 35930
rect 35710 35878 35722 35930
rect 35722 35878 35736 35930
rect 35760 35878 35774 35930
rect 35774 35878 35786 35930
rect 35786 35878 35816 35930
rect 35840 35878 35850 35930
rect 35850 35878 35896 35930
rect 35600 35876 35656 35878
rect 35680 35876 35736 35878
rect 35760 35876 35816 35878
rect 35840 35876 35896 35878
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 35600 34842 35656 34844
rect 35680 34842 35736 34844
rect 35760 34842 35816 34844
rect 35840 34842 35896 34844
rect 35600 34790 35646 34842
rect 35646 34790 35656 34842
rect 35680 34790 35710 34842
rect 35710 34790 35722 34842
rect 35722 34790 35736 34842
rect 35760 34790 35774 34842
rect 35774 34790 35786 34842
rect 35786 34790 35816 34842
rect 35840 34790 35850 34842
rect 35850 34790 35896 34842
rect 35600 34788 35656 34790
rect 35680 34788 35736 34790
rect 35760 34788 35816 34790
rect 35840 34788 35896 34790
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 35600 33754 35656 33756
rect 35680 33754 35736 33756
rect 35760 33754 35816 33756
rect 35840 33754 35896 33756
rect 35600 33702 35646 33754
rect 35646 33702 35656 33754
rect 35680 33702 35710 33754
rect 35710 33702 35722 33754
rect 35722 33702 35736 33754
rect 35760 33702 35774 33754
rect 35774 33702 35786 33754
rect 35786 33702 35816 33754
rect 35840 33702 35850 33754
rect 35850 33702 35896 33754
rect 35600 33700 35656 33702
rect 35680 33700 35736 33702
rect 35760 33700 35816 33702
rect 35840 33700 35896 33702
rect 33322 32272 33378 32328
rect 33506 32544 33562 32600
rect 33598 32272 33654 32328
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 35600 32666 35656 32668
rect 35680 32666 35736 32668
rect 35760 32666 35816 32668
rect 35840 32666 35896 32668
rect 35600 32614 35646 32666
rect 35646 32614 35656 32666
rect 35680 32614 35710 32666
rect 35710 32614 35722 32666
rect 35722 32614 35736 32666
rect 35760 32614 35774 32666
rect 35774 32614 35786 32666
rect 35786 32614 35816 32666
rect 35840 32614 35850 32666
rect 35850 32614 35896 32666
rect 35600 32612 35656 32614
rect 35680 32612 35736 32614
rect 35760 32612 35816 32614
rect 35840 32612 35896 32614
rect 34886 32272 34942 32328
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 35600 31578 35656 31580
rect 35680 31578 35736 31580
rect 35760 31578 35816 31580
rect 35840 31578 35896 31580
rect 35600 31526 35646 31578
rect 35646 31526 35656 31578
rect 35680 31526 35710 31578
rect 35710 31526 35722 31578
rect 35722 31526 35736 31578
rect 35760 31526 35774 31578
rect 35774 31526 35786 31578
rect 35786 31526 35816 31578
rect 35840 31526 35850 31578
rect 35850 31526 35896 31578
rect 35600 31524 35656 31526
rect 35680 31524 35736 31526
rect 35760 31524 35816 31526
rect 35840 31524 35896 31526
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 33782 30540 33784 30560
rect 33784 30540 33836 30560
rect 33836 30540 33838 30560
rect 33782 30504 33838 30540
rect 34610 30504 34666 30560
rect 29182 24384 29238 24440
rect 28906 20576 28962 20632
rect 28906 16632 28962 16688
rect 31666 24656 31722 24712
rect 32310 23160 32366 23216
rect 32586 23160 32642 23216
rect 35600 30490 35656 30492
rect 35680 30490 35736 30492
rect 35760 30490 35816 30492
rect 35840 30490 35896 30492
rect 35600 30438 35646 30490
rect 35646 30438 35656 30490
rect 35680 30438 35710 30490
rect 35710 30438 35722 30490
rect 35722 30438 35736 30490
rect 35760 30438 35774 30490
rect 35774 30438 35786 30490
rect 35786 30438 35816 30490
rect 35840 30438 35850 30490
rect 35850 30438 35896 30490
rect 35600 30436 35656 30438
rect 35680 30436 35736 30438
rect 35760 30436 35816 30438
rect 35840 30436 35896 30438
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 35600 29402 35656 29404
rect 35680 29402 35736 29404
rect 35760 29402 35816 29404
rect 35840 29402 35896 29404
rect 35600 29350 35646 29402
rect 35646 29350 35656 29402
rect 35680 29350 35710 29402
rect 35710 29350 35722 29402
rect 35722 29350 35736 29402
rect 35760 29350 35774 29402
rect 35774 29350 35786 29402
rect 35786 29350 35816 29402
rect 35840 29350 35850 29402
rect 35850 29350 35896 29402
rect 35600 29348 35656 29350
rect 35680 29348 35736 29350
rect 35760 29348 35816 29350
rect 35840 29348 35896 29350
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 35600 28314 35656 28316
rect 35680 28314 35736 28316
rect 35760 28314 35816 28316
rect 35840 28314 35896 28316
rect 35600 28262 35646 28314
rect 35646 28262 35656 28314
rect 35680 28262 35710 28314
rect 35710 28262 35722 28314
rect 35722 28262 35736 28314
rect 35760 28262 35774 28314
rect 35774 28262 35786 28314
rect 35786 28262 35816 28314
rect 35840 28262 35850 28314
rect 35850 28262 35896 28314
rect 35600 28260 35656 28262
rect 35680 28260 35736 28262
rect 35760 28260 35816 28262
rect 35840 28260 35896 28262
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 34058 24404 34114 24440
rect 34058 24384 34060 24404
rect 34060 24384 34112 24404
rect 34112 24384 34114 24404
rect 33966 24248 34022 24304
rect 34334 24248 34390 24304
rect 33598 23568 33654 23624
rect 33322 23160 33378 23216
rect 35600 27226 35656 27228
rect 35680 27226 35736 27228
rect 35760 27226 35816 27228
rect 35840 27226 35896 27228
rect 35600 27174 35646 27226
rect 35646 27174 35656 27226
rect 35680 27174 35710 27226
rect 35710 27174 35722 27226
rect 35722 27174 35736 27226
rect 35760 27174 35774 27226
rect 35774 27174 35786 27226
rect 35786 27174 35816 27226
rect 35840 27174 35850 27226
rect 35850 27174 35896 27226
rect 35600 27172 35656 27174
rect 35680 27172 35736 27174
rect 35760 27172 35816 27174
rect 35840 27172 35896 27174
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 35070 26324 35072 26344
rect 35072 26324 35124 26344
rect 35124 26324 35126 26344
rect 35070 26288 35126 26324
rect 35898 26460 35900 26480
rect 35900 26460 35952 26480
rect 35952 26460 35954 26480
rect 35898 26424 35954 26460
rect 35600 26138 35656 26140
rect 35680 26138 35736 26140
rect 35760 26138 35816 26140
rect 35840 26138 35896 26140
rect 35600 26086 35646 26138
rect 35646 26086 35656 26138
rect 35680 26086 35710 26138
rect 35710 26086 35722 26138
rect 35722 26086 35736 26138
rect 35760 26086 35774 26138
rect 35774 26086 35786 26138
rect 35786 26086 35816 26138
rect 35840 26086 35850 26138
rect 35850 26086 35896 26138
rect 35600 26084 35656 26086
rect 35680 26084 35736 26086
rect 35760 26084 35816 26086
rect 35840 26084 35896 26086
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 36450 26424 36506 26480
rect 36358 26324 36360 26344
rect 36360 26324 36412 26344
rect 36412 26324 36414 26344
rect 36358 26288 36414 26324
rect 35600 25050 35656 25052
rect 35680 25050 35736 25052
rect 35760 25050 35816 25052
rect 35840 25050 35896 25052
rect 35600 24998 35646 25050
rect 35646 24998 35656 25050
rect 35680 24998 35710 25050
rect 35710 24998 35722 25050
rect 35722 24998 35736 25050
rect 35760 24998 35774 25050
rect 35774 24998 35786 25050
rect 35786 24998 35816 25050
rect 35840 24998 35850 25050
rect 35850 24998 35896 25050
rect 35600 24996 35656 24998
rect 35680 24996 35736 24998
rect 35760 24996 35816 24998
rect 35840 24996 35896 24998
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 35162 24112 35218 24168
rect 35622 24248 35678 24304
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 36082 25064 36138 25120
rect 35990 23976 36046 24032
rect 35600 23962 35656 23964
rect 35680 23962 35736 23964
rect 35760 23962 35816 23964
rect 35840 23962 35896 23964
rect 35600 23910 35646 23962
rect 35646 23910 35656 23962
rect 35680 23910 35710 23962
rect 35710 23910 35722 23962
rect 35722 23910 35736 23962
rect 35760 23910 35774 23962
rect 35774 23910 35786 23962
rect 35786 23910 35816 23962
rect 35840 23910 35850 23962
rect 35850 23910 35896 23962
rect 35600 23908 35656 23910
rect 35680 23908 35736 23910
rect 35760 23908 35816 23910
rect 35840 23908 35896 23910
rect 35438 23724 35494 23760
rect 35438 23704 35440 23724
rect 35440 23704 35492 23724
rect 35492 23704 35494 23724
rect 35346 23024 35402 23080
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 31758 20440 31814 20496
rect 29458 16496 29514 16552
rect 29826 19216 29882 19272
rect 29918 17196 29974 17232
rect 29918 17176 29920 17196
rect 29920 17176 29972 17196
rect 29972 17176 29974 17196
rect 30746 16904 30802 16960
rect 31022 17312 31078 17368
rect 31850 18264 31906 18320
rect 31022 16632 31078 16688
rect 31390 16668 31392 16688
rect 31392 16668 31444 16688
rect 31444 16668 31446 16688
rect 31390 16632 31446 16668
rect 31022 16496 31078 16552
rect 34702 20848 34758 20904
rect 34702 20576 34758 20632
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 35622 23044 35678 23080
rect 35622 23024 35624 23044
rect 35624 23024 35676 23044
rect 35676 23024 35678 23044
rect 36174 23160 36230 23216
rect 36174 23024 36230 23080
rect 35600 22874 35656 22876
rect 35680 22874 35736 22876
rect 35760 22874 35816 22876
rect 35840 22874 35896 22876
rect 35600 22822 35646 22874
rect 35646 22822 35656 22874
rect 35680 22822 35710 22874
rect 35710 22822 35722 22874
rect 35722 22822 35736 22874
rect 35760 22822 35774 22874
rect 35774 22822 35786 22874
rect 35786 22822 35816 22874
rect 35840 22822 35850 22874
rect 35850 22822 35896 22874
rect 35600 22820 35656 22822
rect 35680 22820 35736 22822
rect 35760 22820 35816 22822
rect 35840 22820 35896 22822
rect 35622 22344 35678 22400
rect 35898 22516 35900 22536
rect 35900 22516 35952 22536
rect 35952 22516 35954 22536
rect 35898 22480 35954 22516
rect 35600 21786 35656 21788
rect 35680 21786 35736 21788
rect 35760 21786 35816 21788
rect 35840 21786 35896 21788
rect 35600 21734 35646 21786
rect 35646 21734 35656 21786
rect 35680 21734 35710 21786
rect 35710 21734 35722 21786
rect 35722 21734 35736 21786
rect 35760 21734 35774 21786
rect 35774 21734 35786 21786
rect 35786 21734 35816 21786
rect 35840 21734 35850 21786
rect 35850 21734 35896 21786
rect 35600 21732 35656 21734
rect 35680 21732 35736 21734
rect 35760 21732 35816 21734
rect 35840 21732 35896 21734
rect 36634 24384 36690 24440
rect 36818 24656 36874 24712
rect 36818 24268 36874 24304
rect 36818 24248 36820 24268
rect 36820 24248 36872 24268
rect 36872 24248 36874 24268
rect 37002 25236 37004 25256
rect 37004 25236 37056 25256
rect 37056 25236 37058 25256
rect 37002 25200 37058 25236
rect 36818 24112 36874 24168
rect 37738 24384 37794 24440
rect 36818 23840 36874 23896
rect 36358 22344 36414 22400
rect 35600 20698 35656 20700
rect 35680 20698 35736 20700
rect 35760 20698 35816 20700
rect 35840 20698 35896 20700
rect 35600 20646 35646 20698
rect 35646 20646 35656 20698
rect 35680 20646 35710 20698
rect 35710 20646 35722 20698
rect 35722 20646 35736 20698
rect 35760 20646 35774 20698
rect 35774 20646 35786 20698
rect 35786 20646 35816 20698
rect 35840 20646 35850 20698
rect 35850 20646 35896 20698
rect 35600 20644 35656 20646
rect 35680 20644 35736 20646
rect 35760 20644 35816 20646
rect 35840 20644 35896 20646
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 34518 19796 34520 19816
rect 34520 19796 34572 19816
rect 34572 19796 34574 19816
rect 34518 19760 34574 19796
rect 31850 16940 31852 16960
rect 31852 16940 31904 16960
rect 31904 16940 31906 16960
rect 31850 16904 31906 16940
rect 29274 11636 29276 11656
rect 29276 11636 29328 11656
rect 29328 11636 29330 11656
rect 29274 11600 29330 11636
rect 29090 11192 29146 11248
rect 28998 10920 29054 10976
rect 29642 11872 29698 11928
rect 29734 11756 29790 11792
rect 29734 11736 29736 11756
rect 29736 11736 29788 11756
rect 29788 11736 29790 11756
rect 32402 17332 32458 17368
rect 32402 17312 32404 17332
rect 32404 17312 32456 17332
rect 32456 17312 32458 17332
rect 34794 19080 34850 19136
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 35622 19780 35678 19816
rect 35622 19760 35624 19780
rect 35624 19760 35676 19780
rect 35676 19760 35678 19780
rect 35600 19610 35656 19612
rect 35680 19610 35736 19612
rect 35760 19610 35816 19612
rect 35840 19610 35896 19612
rect 35600 19558 35646 19610
rect 35646 19558 35656 19610
rect 35680 19558 35710 19610
rect 35710 19558 35722 19610
rect 35722 19558 35736 19610
rect 35760 19558 35774 19610
rect 35774 19558 35786 19610
rect 35786 19558 35816 19610
rect 35840 19558 35850 19610
rect 35850 19558 35896 19610
rect 35600 19556 35656 19558
rect 35680 19556 35736 19558
rect 35760 19556 35816 19558
rect 35840 19556 35896 19558
rect 36358 20848 36414 20904
rect 36726 22480 36782 22536
rect 36818 20868 36874 20904
rect 36818 20848 36820 20868
rect 36820 20848 36872 20868
rect 36872 20848 36874 20868
rect 35600 18522 35656 18524
rect 35680 18522 35736 18524
rect 35760 18522 35816 18524
rect 35840 18522 35896 18524
rect 35600 18470 35646 18522
rect 35646 18470 35656 18522
rect 35680 18470 35710 18522
rect 35710 18470 35722 18522
rect 35722 18470 35736 18522
rect 35760 18470 35774 18522
rect 35774 18470 35786 18522
rect 35786 18470 35816 18522
rect 35840 18470 35850 18522
rect 35850 18470 35896 18522
rect 35600 18468 35656 18470
rect 35680 18468 35736 18470
rect 35760 18468 35816 18470
rect 35840 18468 35896 18470
rect 35600 17434 35656 17436
rect 35680 17434 35736 17436
rect 35760 17434 35816 17436
rect 35840 17434 35896 17436
rect 35600 17382 35646 17434
rect 35646 17382 35656 17434
rect 35680 17382 35710 17434
rect 35710 17382 35722 17434
rect 35722 17382 35736 17434
rect 35760 17382 35774 17434
rect 35774 17382 35786 17434
rect 35786 17382 35816 17434
rect 35840 17382 35850 17434
rect 35850 17382 35896 17434
rect 35600 17380 35656 17382
rect 35680 17380 35736 17382
rect 35760 17380 35816 17382
rect 35840 17380 35896 17382
rect 35806 16632 35862 16688
rect 36082 16632 36138 16688
rect 35438 16532 35440 16552
rect 35440 16532 35492 16552
rect 35492 16532 35494 16552
rect 35438 16496 35494 16532
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 32586 12280 32642 12336
rect 30930 11192 30986 11248
rect 31022 10920 31078 10976
rect 32218 12144 32274 12200
rect 32402 10648 32458 10704
rect 32310 10512 32366 10568
rect 31850 10104 31906 10160
rect 32310 10124 32366 10160
rect 32310 10104 32312 10124
rect 32312 10104 32364 10124
rect 32364 10104 32366 10124
rect 32494 10104 32550 10160
rect 33046 11872 33102 11928
rect 33322 11892 33378 11928
rect 33322 11872 33324 11892
rect 33324 11872 33376 11892
rect 33376 11872 33378 11892
rect 33690 12280 33746 12336
rect 34242 12300 34298 12336
rect 34242 12280 34244 12300
rect 34244 12280 34296 12300
rect 34296 12280 34298 12300
rect 33782 12180 33784 12200
rect 33784 12180 33836 12200
rect 33836 12180 33838 12200
rect 33598 10104 33654 10160
rect 33782 12144 33838 12180
rect 34610 11600 34666 11656
rect 35600 16346 35656 16348
rect 35680 16346 35736 16348
rect 35760 16346 35816 16348
rect 35840 16346 35896 16348
rect 35600 16294 35646 16346
rect 35646 16294 35656 16346
rect 35680 16294 35710 16346
rect 35710 16294 35722 16346
rect 35722 16294 35736 16346
rect 35760 16294 35774 16346
rect 35774 16294 35786 16346
rect 35786 16294 35816 16346
rect 35840 16294 35850 16346
rect 35850 16294 35896 16346
rect 35600 16292 35656 16294
rect 35680 16292 35736 16294
rect 35760 16292 35816 16294
rect 35840 16292 35896 16294
rect 35600 15258 35656 15260
rect 35680 15258 35736 15260
rect 35760 15258 35816 15260
rect 35840 15258 35896 15260
rect 35600 15206 35646 15258
rect 35646 15206 35656 15258
rect 35680 15206 35710 15258
rect 35710 15206 35722 15258
rect 35722 15206 35736 15258
rect 35760 15206 35774 15258
rect 35774 15206 35786 15258
rect 35786 15206 35816 15258
rect 35840 15206 35850 15258
rect 35850 15206 35896 15258
rect 35600 15204 35656 15206
rect 35680 15204 35736 15206
rect 35760 15204 35816 15206
rect 35840 15204 35896 15206
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 35600 14170 35656 14172
rect 35680 14170 35736 14172
rect 35760 14170 35816 14172
rect 35840 14170 35896 14172
rect 35600 14118 35646 14170
rect 35646 14118 35656 14170
rect 35680 14118 35710 14170
rect 35710 14118 35722 14170
rect 35722 14118 35736 14170
rect 35760 14118 35774 14170
rect 35774 14118 35786 14170
rect 35786 14118 35816 14170
rect 35840 14118 35850 14170
rect 35850 14118 35896 14170
rect 35600 14116 35656 14118
rect 35680 14116 35736 14118
rect 35760 14116 35816 14118
rect 35840 14116 35896 14118
rect 36818 18572 36820 18592
rect 36820 18572 36872 18592
rect 36872 18572 36874 18592
rect 36818 18536 36874 18572
rect 36818 16668 36820 16688
rect 36820 16668 36872 16688
rect 36872 16668 36874 16688
rect 36818 16632 36874 16668
rect 36634 13776 36690 13832
rect 35600 13082 35656 13084
rect 35680 13082 35736 13084
rect 35760 13082 35816 13084
rect 35840 13082 35896 13084
rect 35600 13030 35646 13082
rect 35646 13030 35656 13082
rect 35680 13030 35710 13082
rect 35710 13030 35722 13082
rect 35722 13030 35736 13082
rect 35760 13030 35774 13082
rect 35774 13030 35786 13082
rect 35786 13030 35816 13082
rect 35840 13030 35850 13082
rect 35850 13030 35896 13082
rect 35600 13028 35656 13030
rect 35680 13028 35736 13030
rect 35760 13028 35816 13030
rect 35840 13028 35896 13030
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 35346 12144 35402 12200
rect 35070 11600 35126 11656
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 35600 11994 35656 11996
rect 35680 11994 35736 11996
rect 35760 11994 35816 11996
rect 35840 11994 35896 11996
rect 35600 11942 35646 11994
rect 35646 11942 35656 11994
rect 35680 11942 35710 11994
rect 35710 11942 35722 11994
rect 35722 11942 35736 11994
rect 35760 11942 35774 11994
rect 35774 11942 35786 11994
rect 35786 11942 35816 11994
rect 35840 11942 35850 11994
rect 35850 11942 35896 11994
rect 35600 11940 35656 11942
rect 35680 11940 35736 11942
rect 35760 11940 35816 11942
rect 35840 11940 35896 11942
rect 35070 11192 35126 11248
rect 35346 11076 35402 11112
rect 35346 11056 35348 11076
rect 35348 11056 35400 11076
rect 35400 11056 35402 11076
rect 35600 10906 35656 10908
rect 35680 10906 35736 10908
rect 35760 10906 35816 10908
rect 35840 10906 35896 10908
rect 35600 10854 35646 10906
rect 35646 10854 35656 10906
rect 35680 10854 35710 10906
rect 35710 10854 35722 10906
rect 35722 10854 35736 10906
rect 35760 10854 35774 10906
rect 35774 10854 35786 10906
rect 35786 10854 35816 10906
rect 35840 10854 35850 10906
rect 35850 10854 35896 10906
rect 35600 10852 35656 10854
rect 35680 10852 35736 10854
rect 35760 10852 35816 10854
rect 35840 10852 35896 10854
rect 35070 10684 35072 10704
rect 35072 10684 35124 10704
rect 35124 10684 35126 10704
rect 35070 10648 35126 10684
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 35898 10512 35954 10568
rect 36358 10512 36414 10568
rect 35600 9818 35656 9820
rect 35680 9818 35736 9820
rect 35760 9818 35816 9820
rect 35840 9818 35896 9820
rect 35600 9766 35646 9818
rect 35646 9766 35656 9818
rect 35680 9766 35710 9818
rect 35710 9766 35722 9818
rect 35722 9766 35736 9818
rect 35760 9766 35774 9818
rect 35774 9766 35786 9818
rect 35786 9766 35816 9818
rect 35840 9766 35850 9818
rect 35850 9766 35896 9818
rect 35600 9764 35656 9766
rect 35680 9764 35736 9766
rect 35760 9764 35816 9766
rect 35840 9764 35896 9766
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 35600 8730 35656 8732
rect 35680 8730 35736 8732
rect 35760 8730 35816 8732
rect 35840 8730 35896 8732
rect 35600 8678 35646 8730
rect 35646 8678 35656 8730
rect 35680 8678 35710 8730
rect 35710 8678 35722 8730
rect 35722 8678 35736 8730
rect 35760 8678 35774 8730
rect 35774 8678 35786 8730
rect 35786 8678 35816 8730
rect 35840 8678 35850 8730
rect 35850 8678 35896 8730
rect 35600 8676 35656 8678
rect 35680 8676 35736 8678
rect 35760 8676 35816 8678
rect 35840 8676 35896 8678
rect 37094 18708 37096 18728
rect 37096 18708 37148 18728
rect 37148 18708 37150 18728
rect 37094 18672 37150 18708
rect 37094 17604 37150 17640
rect 37094 17584 37096 17604
rect 37096 17584 37148 17604
rect 37148 17584 37150 17604
rect 37002 16496 37058 16552
rect 37278 16360 37334 16416
rect 38934 28192 38990 28248
rect 40038 28092 40040 28112
rect 40040 28092 40092 28112
rect 40092 28092 40094 28112
rect 40038 28056 40094 28092
rect 38566 23976 38622 24032
rect 38106 23568 38162 23624
rect 38842 25064 38898 25120
rect 38842 24792 38898 24848
rect 38750 24520 38806 24576
rect 39118 25336 39174 25392
rect 37830 20440 37886 20496
rect 39670 23740 39672 23760
rect 39672 23740 39724 23760
rect 39724 23740 39726 23760
rect 39670 23704 39726 23740
rect 38014 18264 38070 18320
rect 37462 15988 37464 16008
rect 37464 15988 37516 16008
rect 37516 15988 37518 16008
rect 37462 15952 37518 15988
rect 38934 18128 38990 18184
rect 38750 17196 38806 17232
rect 38750 17176 38752 17196
rect 38752 17176 38804 17196
rect 38804 17176 38806 17196
rect 38750 16516 38806 16552
rect 38750 16496 38752 16516
rect 38752 16496 38804 16516
rect 38804 16496 38806 16516
rect 39210 18284 39266 18320
rect 39210 18264 39212 18284
rect 39212 18264 39264 18284
rect 39264 18264 39266 18284
rect 39118 18128 39174 18184
rect 40498 24248 40554 24304
rect 40498 23740 40500 23760
rect 40500 23740 40552 23760
rect 40552 23740 40554 23760
rect 40498 23704 40554 23740
rect 39762 22380 39764 22400
rect 39764 22380 39816 22400
rect 39816 22380 39818 22400
rect 39762 22344 39818 22380
rect 39210 16632 39266 16688
rect 40774 24132 40830 24168
rect 40774 24112 40776 24132
rect 40776 24112 40828 24132
rect 40828 24112 40830 24132
rect 40682 23976 40738 24032
rect 39762 17196 39818 17232
rect 39762 17176 39764 17196
rect 39764 17176 39816 17196
rect 39816 17176 39818 17196
rect 41970 25356 42026 25392
rect 41970 25336 41972 25356
rect 41972 25336 42024 25356
rect 42024 25336 42026 25356
rect 42062 25200 42118 25256
rect 40866 23976 40922 24032
rect 41602 23196 41604 23216
rect 41604 23196 41656 23216
rect 41656 23196 41658 23216
rect 41602 23160 41658 23196
rect 42798 28076 42854 28112
rect 42798 28056 42800 28076
rect 42800 28056 42852 28076
rect 42852 28056 42854 28076
rect 43258 28500 43260 28520
rect 43260 28500 43312 28520
rect 43312 28500 43314 28520
rect 43258 28464 43314 28500
rect 42706 25336 42762 25392
rect 42246 23160 42302 23216
rect 42982 24384 43038 24440
rect 43350 24520 43406 24576
rect 45282 28500 45284 28520
rect 45284 28500 45336 28520
rect 45336 28500 45338 28520
rect 45282 28464 45338 28500
rect 43810 25916 43812 25936
rect 43812 25916 43864 25936
rect 43864 25916 43866 25936
rect 43810 25880 43866 25916
rect 43810 24692 43812 24712
rect 43812 24692 43864 24712
rect 43864 24692 43866 24712
rect 43810 24656 43866 24692
rect 42982 23976 43038 24032
rect 43166 23840 43222 23896
rect 42154 23044 42210 23080
rect 42154 23024 42156 23044
rect 42156 23024 42208 23044
rect 42208 23024 42210 23044
rect 40222 16768 40278 16824
rect 39946 15544 40002 15600
rect 39854 15428 39910 15464
rect 39854 15408 39856 15428
rect 39856 15408 39908 15428
rect 39908 15408 39910 15428
rect 39670 15156 39726 15192
rect 39670 15136 39672 15156
rect 39672 15136 39724 15156
rect 39724 15136 39726 15156
rect 40314 14864 40370 14920
rect 37646 12688 37702 12744
rect 38934 12688 38990 12744
rect 38382 11736 38438 11792
rect 37462 11192 37518 11248
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 35600 7642 35656 7644
rect 35680 7642 35736 7644
rect 35760 7642 35816 7644
rect 35840 7642 35896 7644
rect 35600 7590 35646 7642
rect 35646 7590 35656 7642
rect 35680 7590 35710 7642
rect 35710 7590 35722 7642
rect 35722 7590 35736 7642
rect 35760 7590 35774 7642
rect 35774 7590 35786 7642
rect 35786 7590 35816 7642
rect 35840 7590 35850 7642
rect 35850 7590 35896 7642
rect 35600 7588 35656 7590
rect 35680 7588 35736 7590
rect 35760 7588 35816 7590
rect 35840 7588 35896 7590
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 35600 6554 35656 6556
rect 35680 6554 35736 6556
rect 35760 6554 35816 6556
rect 35840 6554 35896 6556
rect 35600 6502 35646 6554
rect 35646 6502 35656 6554
rect 35680 6502 35710 6554
rect 35710 6502 35722 6554
rect 35722 6502 35736 6554
rect 35760 6502 35774 6554
rect 35774 6502 35786 6554
rect 35786 6502 35816 6554
rect 35840 6502 35850 6554
rect 35850 6502 35896 6554
rect 35600 6500 35656 6502
rect 35680 6500 35736 6502
rect 35760 6500 35816 6502
rect 35840 6500 35896 6502
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 35600 5466 35656 5468
rect 35680 5466 35736 5468
rect 35760 5466 35816 5468
rect 35840 5466 35896 5468
rect 35600 5414 35646 5466
rect 35646 5414 35656 5466
rect 35680 5414 35710 5466
rect 35710 5414 35722 5466
rect 35722 5414 35736 5466
rect 35760 5414 35774 5466
rect 35774 5414 35786 5466
rect 35786 5414 35816 5466
rect 35840 5414 35850 5466
rect 35850 5414 35896 5466
rect 35600 5412 35656 5414
rect 35680 5412 35736 5414
rect 35760 5412 35816 5414
rect 35840 5412 35896 5414
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 38198 11056 38254 11112
rect 38750 11756 38806 11792
rect 38750 11736 38752 11756
rect 38752 11736 38804 11756
rect 38804 11736 38806 11756
rect 38842 11192 38898 11248
rect 39210 11192 39266 11248
rect 40958 18128 41014 18184
rect 40866 17856 40922 17912
rect 40866 17312 40922 17368
rect 41142 17992 41198 18048
rect 41142 17584 41198 17640
rect 41142 16496 41198 16552
rect 41602 18284 41658 18320
rect 41602 18264 41604 18284
rect 41604 18264 41656 18284
rect 41656 18264 41658 18284
rect 41510 16668 41512 16688
rect 41512 16668 41564 16688
rect 41564 16668 41566 16688
rect 41510 16632 41566 16668
rect 40682 15544 40738 15600
rect 40958 15428 41014 15464
rect 40958 15408 40960 15428
rect 40960 15408 41012 15428
rect 41012 15408 41014 15428
rect 41142 14864 41198 14920
rect 41050 13524 41106 13560
rect 41050 13504 41052 13524
rect 41052 13504 41104 13524
rect 41104 13504 41106 13524
rect 39946 11192 40002 11248
rect 41602 12280 41658 12336
rect 42154 21528 42210 21584
rect 42982 20576 43038 20632
rect 42890 20460 42946 20496
rect 42890 20440 42892 20460
rect 42892 20440 42944 20460
rect 42944 20440 42946 20460
rect 43442 24248 43498 24304
rect 43442 23976 43498 24032
rect 43626 22344 43682 22400
rect 43810 21936 43866 21992
rect 42706 17856 42762 17912
rect 43166 16768 43222 16824
rect 42062 14592 42118 14648
rect 44086 22344 44142 22400
rect 46938 24792 46994 24848
rect 46386 23432 46442 23488
rect 45466 21528 45522 21584
rect 44914 20576 44970 20632
rect 43810 14612 43866 14648
rect 43810 14592 43812 14612
rect 43812 14592 43864 14612
rect 43864 14592 43866 14612
rect 44086 14864 44142 14920
rect 45558 18672 45614 18728
rect 49514 26460 49516 26480
rect 49516 26460 49568 26480
rect 49568 26460 49570 26480
rect 49514 26424 49570 26460
rect 47214 23840 47270 23896
rect 47122 21936 47178 21992
rect 46846 20884 46848 20904
rect 46848 20884 46900 20904
rect 46900 20884 46902 20904
rect 46846 20848 46902 20884
rect 47306 21936 47362 21992
rect 47214 21800 47270 21856
rect 46110 15952 46166 16008
rect 42890 12144 42946 12200
rect 46662 19216 46718 19272
rect 46938 19352 46994 19408
rect 47582 23840 47638 23896
rect 48318 24112 48374 24168
rect 48042 23840 48098 23896
rect 47950 21140 48006 21176
rect 47950 21120 47952 21140
rect 47952 21120 48004 21140
rect 48004 21120 48006 21140
rect 47858 20596 47914 20632
rect 47858 20576 47860 20596
rect 47860 20576 47912 20596
rect 47912 20576 47914 20596
rect 48502 21528 48558 21584
rect 48962 24556 48964 24576
rect 48964 24556 49016 24576
rect 49016 24556 49018 24576
rect 48962 24520 49018 24556
rect 48594 20984 48650 21040
rect 49238 24692 49240 24712
rect 49240 24692 49292 24712
rect 49292 24692 49294 24712
rect 49238 24656 49294 24692
rect 49146 23976 49202 24032
rect 48962 22888 49018 22944
rect 49054 21528 49110 21584
rect 49606 25200 49662 25256
rect 49330 21664 49386 21720
rect 49238 21528 49294 21584
rect 49238 21256 49294 21312
rect 49238 20984 49294 21040
rect 48778 20712 48834 20768
rect 48594 20440 48650 20496
rect 48318 19488 48374 19544
rect 48410 17856 48466 17912
rect 47214 15136 47270 15192
rect 48226 17720 48282 17776
rect 48778 20168 48834 20224
rect 48686 20032 48742 20088
rect 48594 19896 48650 19952
rect 48594 19760 48650 19816
rect 48502 17040 48558 17096
rect 48226 16496 48282 16552
rect 48042 15580 48044 15600
rect 48044 15580 48096 15600
rect 48096 15580 48098 15600
rect 48042 15544 48098 15580
rect 48962 20032 49018 20088
rect 49146 20712 49202 20768
rect 49514 20440 49570 20496
rect 49238 20168 49294 20224
rect 49054 19624 49110 19680
rect 49238 19216 49294 19272
rect 48778 17856 48834 17912
rect 48778 17176 48834 17232
rect 48594 16224 48650 16280
rect 49054 16904 49110 16960
rect 49790 21936 49846 21992
rect 49790 21256 49846 21312
rect 50434 26444 50490 26480
rect 50434 26424 50436 26444
rect 50436 26424 50488 26444
rect 50488 26424 50490 26444
rect 50158 25236 50160 25256
rect 50160 25236 50212 25256
rect 50212 25236 50214 25256
rect 50158 25200 50214 25236
rect 50066 23432 50122 23488
rect 50434 25764 50490 25800
rect 50434 25744 50436 25764
rect 50436 25744 50488 25764
rect 50488 25744 50490 25764
rect 50802 25200 50858 25256
rect 50710 24828 50712 24848
rect 50712 24828 50764 24848
rect 50764 24828 50766 24848
rect 50710 24792 50766 24828
rect 49790 19760 49846 19816
rect 49790 19660 49792 19680
rect 49792 19660 49844 19680
rect 49844 19660 49846 19680
rect 49790 19624 49846 19660
rect 50158 20984 50214 21040
rect 50158 20576 50214 20632
rect 49974 17176 50030 17232
rect 48502 15000 48558 15056
rect 48410 14864 48466 14920
rect 48686 14864 48742 14920
rect 48502 14728 48558 14784
rect 48778 14356 48780 14376
rect 48780 14356 48832 14376
rect 48832 14356 48834 14376
rect 48778 14320 48834 14356
rect 49698 16244 49754 16280
rect 49698 16224 49700 16244
rect 49700 16224 49752 16244
rect 49752 16224 49754 16244
rect 49054 13932 49110 13968
rect 49054 13912 49056 13932
rect 49056 13912 49108 13932
rect 49108 13912 49110 13932
rect 50710 21256 50766 21312
rect 51262 21140 51318 21176
rect 51262 21120 51264 21140
rect 51264 21120 51316 21140
rect 51316 21120 51318 21140
rect 50802 20984 50858 21040
rect 56690 25900 56746 25936
rect 56690 25880 56692 25900
rect 56692 25880 56744 25900
rect 56744 25880 56746 25900
rect 57886 25880 57942 25936
rect 51262 20712 51318 20768
rect 50434 17040 50490 17096
rect 50618 15272 50674 15328
rect 50802 17040 50858 17096
rect 50802 15408 50858 15464
rect 50434 14340 50490 14376
rect 50434 14320 50436 14340
rect 50436 14320 50488 14340
rect 50488 14320 50490 14340
rect 52550 21528 52606 21584
rect 52182 20884 52184 20904
rect 52184 20884 52236 20904
rect 52236 20884 52238 20904
rect 52182 20848 52238 20884
rect 51170 17720 51226 17776
rect 53838 23432 53894 23488
rect 56874 25744 56930 25800
rect 56690 23024 56746 23080
rect 53378 20032 53434 20088
rect 51630 15408 51686 15464
rect 51630 13932 51686 13968
rect 51630 13912 51632 13932
rect 51632 13912 51684 13932
rect 51684 13912 51686 13932
rect 52366 15136 52422 15192
rect 53010 16904 53066 16960
rect 53378 17448 53434 17504
rect 54942 21256 54998 21312
rect 55402 21800 55458 21856
rect 54574 19896 54630 19952
rect 53746 17196 53802 17232
rect 53746 17176 53748 17196
rect 53748 17176 53800 17196
rect 53800 17176 53802 17196
rect 54206 17484 54208 17504
rect 54208 17484 54260 17504
rect 54260 17484 54262 17504
rect 54206 17448 54262 17484
rect 53562 15444 53564 15464
rect 53564 15444 53616 15464
rect 53616 15444 53618 15464
rect 53562 15408 53618 15444
rect 53194 15272 53250 15328
rect 52826 15000 52882 15056
rect 54758 16108 54814 16144
rect 54758 16088 54760 16108
rect 54760 16088 54812 16108
rect 54812 16088 54814 16108
rect 56690 21564 56692 21584
rect 56692 21564 56744 21584
rect 56744 21564 56746 21584
rect 56690 21528 56746 21564
rect 58438 23160 58494 23216
rect 58438 22500 58494 22536
rect 58438 22480 58440 22500
rect 58440 22480 58492 22500
rect 58492 22480 58494 22500
rect 56874 20440 56930 20496
rect 57886 19080 57942 19136
rect 58438 19760 58494 19816
rect 56782 17584 56838 17640
rect 56690 17176 56746 17232
rect 56322 15444 56324 15464
rect 56324 15444 56376 15464
rect 56376 15444 56378 15464
rect 55678 15272 55734 15328
rect 55034 15000 55090 15056
rect 56322 15408 56378 15444
rect 58438 13676 58440 13696
rect 58440 13676 58492 13696
rect 58492 13676 58494 13696
rect 58438 13640 58494 13676
rect 35600 4378 35656 4380
rect 35680 4378 35736 4380
rect 35760 4378 35816 4380
rect 35840 4378 35896 4380
rect 35600 4326 35646 4378
rect 35646 4326 35656 4378
rect 35680 4326 35710 4378
rect 35710 4326 35722 4378
rect 35722 4326 35736 4378
rect 35760 4326 35774 4378
rect 35774 4326 35786 4378
rect 35786 4326 35816 4378
rect 35840 4326 35850 4378
rect 35850 4326 35896 4378
rect 35600 4324 35656 4326
rect 35680 4324 35736 4326
rect 35760 4324 35816 4326
rect 35840 4324 35896 4326
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 35600 3290 35656 3292
rect 35680 3290 35736 3292
rect 35760 3290 35816 3292
rect 35840 3290 35896 3292
rect 35600 3238 35646 3290
rect 35646 3238 35656 3290
rect 35680 3238 35710 3290
rect 35710 3238 35722 3290
rect 35722 3238 35736 3290
rect 35760 3238 35774 3290
rect 35774 3238 35786 3290
rect 35786 3238 35816 3290
rect 35840 3238 35850 3290
rect 35850 3238 35896 3290
rect 35600 3236 35656 3238
rect 35680 3236 35736 3238
rect 35760 3236 35816 3238
rect 35840 3236 35896 3238
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 35600 2202 35656 2204
rect 35680 2202 35736 2204
rect 35760 2202 35816 2204
rect 35840 2202 35896 2204
rect 35600 2150 35646 2202
rect 35646 2150 35656 2202
rect 35680 2150 35710 2202
rect 35710 2150 35722 2202
rect 35722 2150 35736 2202
rect 35760 2150 35774 2202
rect 35774 2150 35786 2202
rect 35786 2150 35816 2202
rect 35840 2150 35850 2202
rect 35850 2150 35896 2202
rect 35600 2148 35656 2150
rect 35680 2148 35736 2150
rect 35760 2148 35816 2150
rect 35840 2148 35896 2150
<< metal3 >>
rect 4210 37568 4526 37569
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 34930 37568 35246 37569
rect 34930 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35246 37568
rect 34930 37503 35246 37504
rect 4870 37024 5186 37025
rect 4870 36960 4876 37024
rect 4940 36960 4956 37024
rect 5020 36960 5036 37024
rect 5100 36960 5116 37024
rect 5180 36960 5186 37024
rect 4870 36959 5186 36960
rect 35590 37024 35906 37025
rect 35590 36960 35596 37024
rect 35660 36960 35676 37024
rect 35740 36960 35756 37024
rect 35820 36960 35836 37024
rect 35900 36960 35906 37024
rect 35590 36959 35906 36960
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 34930 36480 35246 36481
rect 34930 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35246 36480
rect 34930 36415 35246 36416
rect 4870 35936 5186 35937
rect 4870 35872 4876 35936
rect 4940 35872 4956 35936
rect 5020 35872 5036 35936
rect 5100 35872 5116 35936
rect 5180 35872 5186 35936
rect 4870 35871 5186 35872
rect 35590 35936 35906 35937
rect 35590 35872 35596 35936
rect 35660 35872 35676 35936
rect 35740 35872 35756 35936
rect 35820 35872 35836 35936
rect 35900 35872 35906 35936
rect 35590 35871 35906 35872
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 34930 35392 35246 35393
rect 34930 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35246 35392
rect 34930 35327 35246 35328
rect 4870 34848 5186 34849
rect 4870 34784 4876 34848
rect 4940 34784 4956 34848
rect 5020 34784 5036 34848
rect 5100 34784 5116 34848
rect 5180 34784 5186 34848
rect 4870 34783 5186 34784
rect 35590 34848 35906 34849
rect 35590 34784 35596 34848
rect 35660 34784 35676 34848
rect 35740 34784 35756 34848
rect 35820 34784 35836 34848
rect 35900 34784 35906 34848
rect 35590 34783 35906 34784
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 34930 34304 35246 34305
rect 34930 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35246 34304
rect 34930 34239 35246 34240
rect 4870 33760 5186 33761
rect 4870 33696 4876 33760
rect 4940 33696 4956 33760
rect 5020 33696 5036 33760
rect 5100 33696 5116 33760
rect 5180 33696 5186 33760
rect 4870 33695 5186 33696
rect 35590 33760 35906 33761
rect 35590 33696 35596 33760
rect 35660 33696 35676 33760
rect 35740 33696 35756 33760
rect 35820 33696 35836 33760
rect 35900 33696 35906 33760
rect 35590 33695 35906 33696
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 34930 33216 35246 33217
rect 34930 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35246 33216
rect 34930 33151 35246 33152
rect 4870 32672 5186 32673
rect 4870 32608 4876 32672
rect 4940 32608 4956 32672
rect 5020 32608 5036 32672
rect 5100 32608 5116 32672
rect 5180 32608 5186 32672
rect 4870 32607 5186 32608
rect 35590 32672 35906 32673
rect 35590 32608 35596 32672
rect 35660 32608 35676 32672
rect 35740 32608 35756 32672
rect 35820 32608 35836 32672
rect 35900 32608 35906 32672
rect 35590 32607 35906 32608
rect 33041 32602 33107 32605
rect 33501 32602 33567 32605
rect 33041 32600 33567 32602
rect 33041 32544 33046 32600
rect 33102 32544 33506 32600
rect 33562 32544 33567 32600
rect 33041 32542 33567 32544
rect 33041 32539 33107 32542
rect 33501 32539 33567 32542
rect 33317 32330 33383 32333
rect 33593 32330 33659 32333
rect 34881 32330 34947 32333
rect 33317 32328 34947 32330
rect 33317 32272 33322 32328
rect 33378 32272 33598 32328
rect 33654 32272 34886 32328
rect 34942 32272 34947 32328
rect 33317 32270 34947 32272
rect 33317 32267 33383 32270
rect 33593 32267 33659 32270
rect 34881 32267 34947 32270
rect 4210 32128 4526 32129
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 34930 32128 35246 32129
rect 34930 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35246 32128
rect 34930 32063 35246 32064
rect 4870 31584 5186 31585
rect 4870 31520 4876 31584
rect 4940 31520 4956 31584
rect 5020 31520 5036 31584
rect 5100 31520 5116 31584
rect 5180 31520 5186 31584
rect 4870 31519 5186 31520
rect 35590 31584 35906 31585
rect 35590 31520 35596 31584
rect 35660 31520 35676 31584
rect 35740 31520 35756 31584
rect 35820 31520 35836 31584
rect 35900 31520 35906 31584
rect 35590 31519 35906 31520
rect 19701 31514 19767 31517
rect 23381 31514 23447 31517
rect 19701 31512 23447 31514
rect 19701 31456 19706 31512
rect 19762 31456 23386 31512
rect 23442 31456 23447 31512
rect 19701 31454 23447 31456
rect 19701 31451 19767 31454
rect 23381 31451 23447 31454
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 34930 31040 35246 31041
rect 34930 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35246 31040
rect 34930 30975 35246 30976
rect 33777 30562 33843 30565
rect 34605 30562 34671 30565
rect 33777 30560 34671 30562
rect 33777 30504 33782 30560
rect 33838 30504 34610 30560
rect 34666 30504 34671 30560
rect 33777 30502 34671 30504
rect 33777 30499 33843 30502
rect 34605 30499 34671 30502
rect 4870 30496 5186 30497
rect 4870 30432 4876 30496
rect 4940 30432 4956 30496
rect 5020 30432 5036 30496
rect 5100 30432 5116 30496
rect 5180 30432 5186 30496
rect 4870 30431 5186 30432
rect 35590 30496 35906 30497
rect 35590 30432 35596 30496
rect 35660 30432 35676 30496
rect 35740 30432 35756 30496
rect 35820 30432 35836 30496
rect 35900 30432 35906 30496
rect 35590 30431 35906 30432
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 34930 29952 35246 29953
rect 34930 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35246 29952
rect 34930 29887 35246 29888
rect 4870 29408 5186 29409
rect 4870 29344 4876 29408
rect 4940 29344 4956 29408
rect 5020 29344 5036 29408
rect 5100 29344 5116 29408
rect 5180 29344 5186 29408
rect 4870 29343 5186 29344
rect 35590 29408 35906 29409
rect 35590 29344 35596 29408
rect 35660 29344 35676 29408
rect 35740 29344 35756 29408
rect 35820 29344 35836 29408
rect 35900 29344 35906 29408
rect 35590 29343 35906 29344
rect 28073 29068 28139 29069
rect 28022 29004 28028 29068
rect 28092 29066 28139 29068
rect 28092 29064 28184 29066
rect 28134 29008 28184 29064
rect 28092 29006 28184 29008
rect 28092 29004 28139 29006
rect 28073 29003 28139 29004
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 34930 28864 35246 28865
rect 34930 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35246 28864
rect 34930 28799 35246 28800
rect 43253 28522 43319 28525
rect 45277 28522 45343 28525
rect 43253 28520 45343 28522
rect 43253 28464 43258 28520
rect 43314 28464 45282 28520
rect 45338 28464 45343 28520
rect 43253 28462 45343 28464
rect 43253 28459 43319 28462
rect 45277 28459 45343 28462
rect 4870 28320 5186 28321
rect 4870 28256 4876 28320
rect 4940 28256 4956 28320
rect 5020 28256 5036 28320
rect 5100 28256 5116 28320
rect 5180 28256 5186 28320
rect 4870 28255 5186 28256
rect 35590 28320 35906 28321
rect 35590 28256 35596 28320
rect 35660 28256 35676 28320
rect 35740 28256 35756 28320
rect 35820 28256 35836 28320
rect 35900 28256 35906 28320
rect 35590 28255 35906 28256
rect 38929 28250 38995 28253
rect 39982 28250 39988 28252
rect 38929 28248 39988 28250
rect 38929 28192 38934 28248
rect 38990 28192 39988 28248
rect 38929 28190 39988 28192
rect 38929 28187 38995 28190
rect 39982 28188 39988 28190
rect 40052 28188 40058 28252
rect 40033 28114 40099 28117
rect 42793 28114 42859 28117
rect 40033 28112 42859 28114
rect 40033 28056 40038 28112
rect 40094 28056 42798 28112
rect 42854 28056 42859 28112
rect 40033 28054 42859 28056
rect 40033 28051 40099 28054
rect 42793 28051 42859 28054
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 34930 27776 35246 27777
rect 34930 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35246 27776
rect 34930 27711 35246 27712
rect 4870 27232 5186 27233
rect 4870 27168 4876 27232
rect 4940 27168 4956 27232
rect 5020 27168 5036 27232
rect 5100 27168 5116 27232
rect 5180 27168 5186 27232
rect 4870 27167 5186 27168
rect 35590 27232 35906 27233
rect 35590 27168 35596 27232
rect 35660 27168 35676 27232
rect 35740 27168 35756 27232
rect 35820 27168 35836 27232
rect 35900 27168 35906 27232
rect 35590 27167 35906 27168
rect 4210 26688 4526 26689
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 34930 26688 35246 26689
rect 34930 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35246 26688
rect 34930 26623 35246 26624
rect 35893 26482 35959 26485
rect 36445 26482 36511 26485
rect 35893 26480 36511 26482
rect 35893 26424 35898 26480
rect 35954 26424 36450 26480
rect 36506 26424 36511 26480
rect 35893 26422 36511 26424
rect 35893 26419 35959 26422
rect 36445 26419 36511 26422
rect 49509 26482 49575 26485
rect 50429 26482 50495 26485
rect 49509 26480 50495 26482
rect 49509 26424 49514 26480
rect 49570 26424 50434 26480
rect 50490 26424 50495 26480
rect 49509 26422 50495 26424
rect 49509 26419 49575 26422
rect 50429 26419 50495 26422
rect 25037 26346 25103 26349
rect 25957 26346 26023 26349
rect 27705 26346 27771 26349
rect 28441 26346 28507 26349
rect 25037 26344 28507 26346
rect 25037 26288 25042 26344
rect 25098 26288 25962 26344
rect 26018 26288 27710 26344
rect 27766 26288 28446 26344
rect 28502 26288 28507 26344
rect 25037 26286 28507 26288
rect 25037 26283 25103 26286
rect 25957 26283 26023 26286
rect 27705 26283 27771 26286
rect 28441 26283 28507 26286
rect 35065 26346 35131 26349
rect 36353 26346 36419 26349
rect 35065 26344 36419 26346
rect 35065 26288 35070 26344
rect 35126 26288 36358 26344
rect 36414 26288 36419 26344
rect 35065 26286 36419 26288
rect 35065 26283 35131 26286
rect 36353 26283 36419 26286
rect 4870 26144 5186 26145
rect 4870 26080 4876 26144
rect 4940 26080 4956 26144
rect 5020 26080 5036 26144
rect 5100 26080 5116 26144
rect 5180 26080 5186 26144
rect 4870 26079 5186 26080
rect 35590 26144 35906 26145
rect 35590 26080 35596 26144
rect 35660 26080 35676 26144
rect 35740 26080 35756 26144
rect 35820 26080 35836 26144
rect 35900 26080 35906 26144
rect 35590 26079 35906 26080
rect 43805 25938 43871 25941
rect 56685 25938 56751 25941
rect 43805 25936 56751 25938
rect 43805 25880 43810 25936
rect 43866 25880 56690 25936
rect 56746 25880 56751 25936
rect 43805 25878 56751 25880
rect 43805 25875 43871 25878
rect 56685 25875 56751 25878
rect 57881 25938 57947 25941
rect 59200 25938 60000 25968
rect 57881 25936 60000 25938
rect 57881 25880 57886 25936
rect 57942 25880 60000 25936
rect 57881 25878 60000 25880
rect 57881 25875 57947 25878
rect 59200 25848 60000 25878
rect 50429 25802 50495 25805
rect 56869 25802 56935 25805
rect 50429 25800 56935 25802
rect 50429 25744 50434 25800
rect 50490 25744 56874 25800
rect 56930 25744 56935 25800
rect 50429 25742 56935 25744
rect 50429 25739 50495 25742
rect 56869 25739 56935 25742
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 34930 25600 35246 25601
rect 34930 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35246 25600
rect 34930 25535 35246 25536
rect 39113 25394 39179 25397
rect 41965 25394 42031 25397
rect 42701 25394 42767 25397
rect 39113 25392 42031 25394
rect 39113 25336 39118 25392
rect 39174 25336 41970 25392
rect 42026 25336 42031 25392
rect 39113 25334 42031 25336
rect 39113 25331 39179 25334
rect 41965 25331 42031 25334
rect 42198 25392 42767 25394
rect 42198 25336 42706 25392
rect 42762 25336 42767 25392
rect 42198 25334 42767 25336
rect 21725 25258 21791 25261
rect 23289 25258 23355 25261
rect 21725 25256 23355 25258
rect 21725 25200 21730 25256
rect 21786 25200 23294 25256
rect 23350 25200 23355 25256
rect 21725 25198 23355 25200
rect 21725 25195 21791 25198
rect 23289 25195 23355 25198
rect 28993 25258 29059 25261
rect 36997 25258 37063 25261
rect 42057 25258 42123 25261
rect 42198 25258 42258 25334
rect 42701 25331 42767 25334
rect 28993 25256 37063 25258
rect 28993 25200 28998 25256
rect 29054 25200 37002 25256
rect 37058 25200 37063 25256
rect 28993 25198 37063 25200
rect 28993 25195 29059 25198
rect 36997 25195 37063 25198
rect 41370 25256 42258 25258
rect 41370 25200 42062 25256
rect 42118 25200 42258 25256
rect 41370 25198 42258 25200
rect 49601 25258 49667 25261
rect 49734 25258 49740 25260
rect 49601 25256 49740 25258
rect 49601 25200 49606 25256
rect 49662 25200 49740 25256
rect 49601 25198 49740 25200
rect 19425 25122 19491 25125
rect 23013 25122 23079 25125
rect 36077 25124 36143 25125
rect 36077 25122 36124 25124
rect 19425 25120 23079 25122
rect 19425 25064 19430 25120
rect 19486 25064 23018 25120
rect 23074 25064 23079 25120
rect 19425 25062 23079 25064
rect 36032 25120 36124 25122
rect 36032 25064 36082 25120
rect 36032 25062 36124 25064
rect 19425 25059 19491 25062
rect 23013 25059 23079 25062
rect 36077 25060 36124 25062
rect 36188 25060 36194 25124
rect 38837 25122 38903 25125
rect 41370 25122 41430 25198
rect 42057 25195 42123 25198
rect 49601 25195 49667 25198
rect 49734 25196 49740 25198
rect 49804 25258 49810 25260
rect 50153 25258 50219 25261
rect 50797 25258 50863 25261
rect 49804 25256 50863 25258
rect 49804 25200 50158 25256
rect 50214 25200 50802 25256
rect 50858 25200 50863 25256
rect 49804 25198 50863 25200
rect 49804 25196 49810 25198
rect 50153 25195 50219 25198
rect 50797 25195 50863 25198
rect 38837 25120 41430 25122
rect 38837 25064 38842 25120
rect 38898 25064 41430 25120
rect 38837 25062 41430 25064
rect 36077 25059 36143 25060
rect 38837 25059 38903 25062
rect 4870 25056 5186 25057
rect 4870 24992 4876 25056
rect 4940 24992 4956 25056
rect 5020 24992 5036 25056
rect 5100 24992 5116 25056
rect 5180 24992 5186 25056
rect 4870 24991 5186 24992
rect 35590 25056 35906 25057
rect 35590 24992 35596 25056
rect 35660 24992 35676 25056
rect 35740 24992 35756 25056
rect 35820 24992 35836 25056
rect 35900 24992 35906 25056
rect 35590 24991 35906 24992
rect 25313 24852 25379 24853
rect 25262 24850 25268 24852
rect 25186 24790 25268 24850
rect 25332 24850 25379 24852
rect 38837 24850 38903 24853
rect 25332 24848 38903 24850
rect 25374 24792 38842 24848
rect 38898 24792 38903 24848
rect 25262 24788 25268 24790
rect 25332 24790 38903 24792
rect 25332 24788 25379 24790
rect 25313 24787 25379 24788
rect 38837 24787 38903 24790
rect 46933 24850 46999 24853
rect 48446 24850 48452 24852
rect 46933 24848 48452 24850
rect 46933 24792 46938 24848
rect 46994 24792 48452 24848
rect 46933 24790 48452 24792
rect 46933 24787 46999 24790
rect 48446 24788 48452 24790
rect 48516 24850 48522 24852
rect 50705 24850 50771 24853
rect 48516 24848 50771 24850
rect 48516 24792 50710 24848
rect 50766 24792 50771 24848
rect 48516 24790 50771 24792
rect 48516 24788 48522 24790
rect 50705 24787 50771 24790
rect 31661 24714 31727 24717
rect 36813 24714 36879 24717
rect 31661 24712 36879 24714
rect 31661 24656 31666 24712
rect 31722 24656 36818 24712
rect 36874 24656 36879 24712
rect 31661 24654 36879 24656
rect 31661 24651 31727 24654
rect 36813 24651 36879 24654
rect 43805 24714 43871 24717
rect 49233 24714 49299 24717
rect 43805 24712 49299 24714
rect 43805 24656 43810 24712
rect 43866 24656 49238 24712
rect 49294 24656 49299 24712
rect 43805 24654 49299 24656
rect 43805 24651 43871 24654
rect 49233 24651 49299 24654
rect 22829 24578 22895 24581
rect 27521 24578 27587 24581
rect 22829 24576 27587 24578
rect 22829 24520 22834 24576
rect 22890 24520 27526 24576
rect 27582 24520 27587 24576
rect 22829 24518 27587 24520
rect 22829 24515 22895 24518
rect 27521 24515 27587 24518
rect 38745 24578 38811 24581
rect 43345 24578 43411 24581
rect 48957 24578 49023 24581
rect 38745 24576 49023 24578
rect 38745 24520 38750 24576
rect 38806 24520 43350 24576
rect 43406 24520 48962 24576
rect 49018 24520 49023 24576
rect 38745 24518 49023 24520
rect 38745 24515 38811 24518
rect 43345 24515 43411 24518
rect 48957 24515 49023 24518
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 34930 24512 35246 24513
rect 34930 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35246 24512
rect 34930 24447 35246 24448
rect 25773 24442 25839 24445
rect 26509 24442 26575 24445
rect 25773 24440 26575 24442
rect 25773 24384 25778 24440
rect 25834 24384 26514 24440
rect 26570 24384 26575 24440
rect 25773 24382 26575 24384
rect 25773 24379 25839 24382
rect 26509 24379 26575 24382
rect 28441 24442 28507 24445
rect 28809 24442 28875 24445
rect 28441 24440 28875 24442
rect 28441 24384 28446 24440
rect 28502 24384 28814 24440
rect 28870 24384 28875 24440
rect 28441 24382 28875 24384
rect 28441 24379 28507 24382
rect 28809 24379 28875 24382
rect 29177 24442 29243 24445
rect 34053 24442 34119 24445
rect 36629 24442 36695 24445
rect 37733 24442 37799 24445
rect 42977 24442 43043 24445
rect 29177 24440 34119 24442
rect 29177 24384 29182 24440
rect 29238 24384 34058 24440
rect 34114 24384 34119 24440
rect 29177 24382 34119 24384
rect 29177 24379 29243 24382
rect 34053 24379 34119 24382
rect 35390 24440 43043 24442
rect 35390 24384 36634 24440
rect 36690 24384 37738 24440
rect 37794 24384 42982 24440
rect 43038 24384 43043 24440
rect 35390 24382 43043 24384
rect 22369 24306 22435 24309
rect 22921 24306 22987 24309
rect 26325 24306 26391 24309
rect 33961 24306 34027 24309
rect 22369 24304 22987 24306
rect 22369 24248 22374 24304
rect 22430 24248 22926 24304
rect 22982 24248 22987 24304
rect 22369 24246 22987 24248
rect 22369 24243 22435 24246
rect 22921 24243 22987 24246
rect 25454 24304 34027 24306
rect 25454 24248 26330 24304
rect 26386 24248 33966 24304
rect 34022 24248 34027 24304
rect 25454 24246 34027 24248
rect 25454 24037 25514 24246
rect 26325 24243 26391 24246
rect 33961 24243 34027 24246
rect 34329 24306 34395 24309
rect 35390 24306 35450 24382
rect 36629 24379 36695 24382
rect 37733 24379 37799 24382
rect 42977 24379 43043 24382
rect 34329 24304 35450 24306
rect 34329 24248 34334 24304
rect 34390 24248 35450 24304
rect 34329 24246 35450 24248
rect 35617 24306 35683 24309
rect 36813 24306 36879 24309
rect 35617 24304 36879 24306
rect 35617 24248 35622 24304
rect 35678 24248 36818 24304
rect 36874 24248 36879 24304
rect 35617 24246 36879 24248
rect 34329 24243 34395 24246
rect 35617 24243 35683 24246
rect 36813 24243 36879 24246
rect 40493 24306 40559 24309
rect 43437 24306 43503 24309
rect 40493 24304 43503 24306
rect 40493 24248 40498 24304
rect 40554 24248 43442 24304
rect 43498 24248 43503 24304
rect 40493 24246 43503 24248
rect 40493 24243 40559 24246
rect 43437 24243 43503 24246
rect 26325 24170 26391 24173
rect 35157 24170 35223 24173
rect 36813 24170 36879 24173
rect 26325 24168 36879 24170
rect 26325 24112 26330 24168
rect 26386 24112 35162 24168
rect 35218 24112 36818 24168
rect 36874 24112 36879 24168
rect 26325 24110 36879 24112
rect 26325 24107 26391 24110
rect 35157 24107 35223 24110
rect 36813 24107 36879 24110
rect 40769 24170 40835 24173
rect 48313 24170 48379 24173
rect 40769 24168 48379 24170
rect 40769 24112 40774 24168
rect 40830 24112 48318 24168
rect 48374 24112 48379 24168
rect 40769 24110 48379 24112
rect 40769 24107 40835 24110
rect 48313 24107 48379 24110
rect 22093 24034 22159 24037
rect 23841 24034 23907 24037
rect 22093 24032 23907 24034
rect 22093 23976 22098 24032
rect 22154 23976 23846 24032
rect 23902 23976 23907 24032
rect 22093 23974 23907 23976
rect 22093 23971 22159 23974
rect 23841 23971 23907 23974
rect 25405 24032 25514 24037
rect 25405 23976 25410 24032
rect 25466 23976 25514 24032
rect 25405 23974 25514 23976
rect 35985 24034 36051 24037
rect 38561 24034 38627 24037
rect 40677 24034 40743 24037
rect 35985 24032 40743 24034
rect 35985 23976 35990 24032
rect 36046 23976 38566 24032
rect 38622 23976 40682 24032
rect 40738 23976 40743 24032
rect 35985 23974 40743 23976
rect 25405 23971 25471 23974
rect 35985 23971 36051 23974
rect 38561 23971 38627 23974
rect 40677 23971 40743 23974
rect 40861 24034 40927 24037
rect 42977 24034 43043 24037
rect 40861 24032 43043 24034
rect 40861 23976 40866 24032
rect 40922 23976 42982 24032
rect 43038 23976 43043 24032
rect 40861 23974 43043 23976
rect 40861 23971 40927 23974
rect 42977 23971 43043 23974
rect 43437 24034 43503 24037
rect 49141 24034 49207 24037
rect 43437 24032 49207 24034
rect 43437 23976 43442 24032
rect 43498 23976 49146 24032
rect 49202 23976 49207 24032
rect 43437 23974 49207 23976
rect 43437 23971 43503 23974
rect 49141 23971 49207 23974
rect 4870 23968 5186 23969
rect 4870 23904 4876 23968
rect 4940 23904 4956 23968
rect 5020 23904 5036 23968
rect 5100 23904 5116 23968
rect 5180 23904 5186 23968
rect 4870 23903 5186 23904
rect 35590 23968 35906 23969
rect 35590 23904 35596 23968
rect 35660 23904 35676 23968
rect 35740 23904 35756 23968
rect 35820 23904 35836 23968
rect 35900 23904 35906 23968
rect 35590 23903 35906 23904
rect 20989 23898 21055 23901
rect 22553 23898 22619 23901
rect 25589 23898 25655 23901
rect 20989 23896 25655 23898
rect 20989 23840 20994 23896
rect 21050 23840 22558 23896
rect 22614 23840 25594 23896
rect 25650 23840 25655 23896
rect 20989 23838 25655 23840
rect 20989 23835 21055 23838
rect 22553 23835 22619 23838
rect 25589 23835 25655 23838
rect 36813 23898 36879 23901
rect 40718 23898 40724 23900
rect 36813 23896 40724 23898
rect 36813 23840 36818 23896
rect 36874 23840 40724 23896
rect 36813 23838 40724 23840
rect 36813 23835 36879 23838
rect 40718 23836 40724 23838
rect 40788 23898 40794 23900
rect 43161 23898 43227 23901
rect 47209 23898 47275 23901
rect 47577 23898 47643 23901
rect 48037 23898 48103 23901
rect 40788 23896 48103 23898
rect 40788 23840 43166 23896
rect 43222 23840 47214 23896
rect 47270 23840 47582 23896
rect 47638 23840 48042 23896
rect 48098 23840 48103 23896
rect 40788 23838 48103 23840
rect 40788 23836 40794 23838
rect 43161 23835 43227 23838
rect 47209 23835 47275 23838
rect 47577 23835 47643 23838
rect 48037 23835 48103 23838
rect 27061 23762 27127 23765
rect 35433 23762 35499 23765
rect 27061 23760 35499 23762
rect 27061 23704 27066 23760
rect 27122 23704 35438 23760
rect 35494 23704 35499 23760
rect 27061 23702 35499 23704
rect 27061 23699 27127 23702
rect 35433 23699 35499 23702
rect 39665 23762 39731 23765
rect 40493 23762 40559 23765
rect 39665 23760 40559 23762
rect 39665 23704 39670 23760
rect 39726 23704 40498 23760
rect 40554 23704 40559 23760
rect 39665 23702 40559 23704
rect 39665 23699 39731 23702
rect 40493 23699 40559 23702
rect 25865 23626 25931 23629
rect 27654 23626 27660 23628
rect 25865 23624 27660 23626
rect 25865 23568 25870 23624
rect 25926 23568 27660 23624
rect 25865 23566 27660 23568
rect 25865 23563 25931 23566
rect 27654 23564 27660 23566
rect 27724 23626 27730 23628
rect 27797 23626 27863 23629
rect 27724 23624 27863 23626
rect 27724 23568 27802 23624
rect 27858 23568 27863 23624
rect 27724 23566 27863 23568
rect 27724 23564 27730 23566
rect 27797 23563 27863 23566
rect 33593 23626 33659 23629
rect 38101 23626 38167 23629
rect 33593 23624 38167 23626
rect 33593 23568 33598 23624
rect 33654 23568 38106 23624
rect 38162 23568 38167 23624
rect 33593 23566 38167 23568
rect 33593 23563 33659 23566
rect 38101 23563 38167 23566
rect 46381 23490 46447 23493
rect 50061 23490 50127 23493
rect 53833 23490 53899 23493
rect 46381 23488 53899 23490
rect 46381 23432 46386 23488
rect 46442 23432 50066 23488
rect 50122 23432 53838 23488
rect 53894 23432 53899 23488
rect 46381 23430 53899 23432
rect 46381 23427 46447 23430
rect 50061 23427 50127 23430
rect 53833 23427 53899 23430
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 34930 23424 35246 23425
rect 34930 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35246 23424
rect 34930 23359 35246 23360
rect 27337 23218 27403 23221
rect 32305 23218 32371 23221
rect 27337 23216 32371 23218
rect 27337 23160 27342 23216
rect 27398 23160 32310 23216
rect 32366 23160 32371 23216
rect 27337 23158 32371 23160
rect 27337 23155 27403 23158
rect 32305 23155 32371 23158
rect 32581 23218 32647 23221
rect 33317 23218 33383 23221
rect 36169 23218 36235 23221
rect 32581 23216 36235 23218
rect 32581 23160 32586 23216
rect 32642 23160 33322 23216
rect 33378 23160 36174 23216
rect 36230 23160 36235 23216
rect 32581 23158 36235 23160
rect 32581 23155 32647 23158
rect 33317 23155 33383 23158
rect 36169 23155 36235 23158
rect 41597 23218 41663 23221
rect 42241 23218 42307 23221
rect 41597 23216 42307 23218
rect 41597 23160 41602 23216
rect 41658 23160 42246 23216
rect 42302 23160 42307 23216
rect 41597 23158 42307 23160
rect 41597 23155 41663 23158
rect 42241 23155 42307 23158
rect 58433 23218 58499 23221
rect 59200 23218 60000 23248
rect 58433 23216 60000 23218
rect 58433 23160 58438 23216
rect 58494 23160 60000 23216
rect 58433 23158 60000 23160
rect 58433 23155 58499 23158
rect 59200 23128 60000 23158
rect 35341 23082 35407 23085
rect 35617 23082 35683 23085
rect 36169 23084 36235 23085
rect 36118 23082 36124 23084
rect 35341 23080 36124 23082
rect 36188 23080 36235 23084
rect 35341 23024 35346 23080
rect 35402 23024 35622 23080
rect 35678 23024 36124 23080
rect 36230 23024 36235 23080
rect 35341 23022 36124 23024
rect 35341 23019 35407 23022
rect 35617 23019 35683 23022
rect 36118 23020 36124 23022
rect 36188 23020 36235 23024
rect 36169 23019 36235 23020
rect 42149 23082 42215 23085
rect 56685 23082 56751 23085
rect 42149 23080 56751 23082
rect 42149 23024 42154 23080
rect 42210 23024 56690 23080
rect 56746 23024 56751 23080
rect 42149 23022 56751 23024
rect 42149 23019 42215 23022
rect 56685 23019 56751 23022
rect 48957 22948 49023 22949
rect 48957 22946 49004 22948
rect 48912 22944 49004 22946
rect 48912 22888 48962 22944
rect 48912 22886 49004 22888
rect 48957 22884 49004 22886
rect 49068 22884 49074 22948
rect 48957 22883 49023 22884
rect 4870 22880 5186 22881
rect 4870 22816 4876 22880
rect 4940 22816 4956 22880
rect 5020 22816 5036 22880
rect 5100 22816 5116 22880
rect 5180 22816 5186 22880
rect 4870 22815 5186 22816
rect 35590 22880 35906 22881
rect 35590 22816 35596 22880
rect 35660 22816 35676 22880
rect 35740 22816 35756 22880
rect 35820 22816 35836 22880
rect 35900 22816 35906 22880
rect 35590 22815 35906 22816
rect 20437 22538 20503 22541
rect 20118 22536 20503 22538
rect 20118 22480 20442 22536
rect 20498 22480 20503 22536
rect 20118 22478 20503 22480
rect 20118 22405 20178 22478
rect 20437 22475 20503 22478
rect 35893 22538 35959 22541
rect 36721 22538 36787 22541
rect 35893 22536 36787 22538
rect 35893 22480 35898 22536
rect 35954 22480 36726 22536
rect 36782 22480 36787 22536
rect 35893 22478 36787 22480
rect 35893 22475 35959 22478
rect 36721 22475 36787 22478
rect 58433 22538 58499 22541
rect 59200 22538 60000 22568
rect 58433 22536 60000 22538
rect 58433 22480 58438 22536
rect 58494 22480 60000 22536
rect 58433 22478 60000 22480
rect 58433 22475 58499 22478
rect 59200 22448 60000 22478
rect 20069 22400 20178 22405
rect 20069 22344 20074 22400
rect 20130 22344 20178 22400
rect 20069 22342 20178 22344
rect 35617 22402 35683 22405
rect 36353 22402 36419 22405
rect 35617 22400 36419 22402
rect 35617 22344 35622 22400
rect 35678 22344 36358 22400
rect 36414 22344 36419 22400
rect 35617 22342 36419 22344
rect 20069 22339 20135 22342
rect 35617 22339 35683 22342
rect 36353 22339 36419 22342
rect 39614 22340 39620 22404
rect 39684 22402 39690 22404
rect 39757 22402 39823 22405
rect 39684 22400 39823 22402
rect 39684 22344 39762 22400
rect 39818 22344 39823 22400
rect 39684 22342 39823 22344
rect 39684 22340 39690 22342
rect 39757 22339 39823 22342
rect 43621 22402 43687 22405
rect 44081 22402 44147 22405
rect 43621 22400 44147 22402
rect 43621 22344 43626 22400
rect 43682 22344 44086 22400
rect 44142 22344 44147 22400
rect 43621 22342 44147 22344
rect 43621 22339 43687 22342
rect 44081 22339 44147 22342
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 34930 22336 35246 22337
rect 34930 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35246 22336
rect 34930 22271 35246 22272
rect 19885 21994 19951 21997
rect 27429 21994 27495 21997
rect 28022 21994 28028 21996
rect 19885 21992 28028 21994
rect 19885 21936 19890 21992
rect 19946 21936 27434 21992
rect 27490 21936 28028 21992
rect 19885 21934 28028 21936
rect 19885 21931 19951 21934
rect 27429 21931 27495 21934
rect 28022 21932 28028 21934
rect 28092 21932 28098 21996
rect 43805 21994 43871 21997
rect 47117 21994 47183 21997
rect 43805 21992 47183 21994
rect 43805 21936 43810 21992
rect 43866 21936 47122 21992
rect 47178 21936 47183 21992
rect 43805 21934 47183 21936
rect 43805 21931 43871 21934
rect 47117 21931 47183 21934
rect 47301 21994 47367 21997
rect 49785 21994 49851 21997
rect 47301 21992 49851 21994
rect 47301 21936 47306 21992
rect 47362 21936 49790 21992
rect 49846 21936 49851 21992
rect 47301 21934 49851 21936
rect 47301 21931 47367 21934
rect 49785 21931 49851 21934
rect 47209 21858 47275 21861
rect 55397 21858 55463 21861
rect 47209 21856 55463 21858
rect 47209 21800 47214 21856
rect 47270 21800 55402 21856
rect 55458 21800 55463 21856
rect 47209 21798 55463 21800
rect 47209 21795 47275 21798
rect 55397 21795 55463 21798
rect 4870 21792 5186 21793
rect 4870 21728 4876 21792
rect 4940 21728 4956 21792
rect 5020 21728 5036 21792
rect 5100 21728 5116 21792
rect 5180 21728 5186 21792
rect 4870 21727 5186 21728
rect 35590 21792 35906 21793
rect 35590 21728 35596 21792
rect 35660 21728 35676 21792
rect 35740 21728 35756 21792
rect 35820 21728 35836 21792
rect 35900 21728 35906 21792
rect 35590 21727 35906 21728
rect 20437 21722 20503 21725
rect 23841 21722 23907 21725
rect 20437 21720 23907 21722
rect 20437 21664 20442 21720
rect 20498 21664 23846 21720
rect 23902 21664 23907 21720
rect 20437 21662 23907 21664
rect 20437 21659 20503 21662
rect 23841 21659 23907 21662
rect 49182 21660 49188 21724
rect 49252 21722 49258 21724
rect 49325 21722 49391 21725
rect 49252 21720 49391 21722
rect 49252 21664 49330 21720
rect 49386 21664 49391 21720
rect 49252 21662 49391 21664
rect 49252 21660 49258 21662
rect 49325 21659 49391 21662
rect 42149 21586 42215 21589
rect 45461 21586 45527 21589
rect 42149 21584 45527 21586
rect 42149 21528 42154 21584
rect 42210 21528 45466 21584
rect 45522 21528 45527 21584
rect 42149 21526 45527 21528
rect 42149 21523 42215 21526
rect 45461 21523 45527 21526
rect 48497 21586 48563 21589
rect 49049 21586 49115 21589
rect 48497 21584 49115 21586
rect 48497 21528 48502 21584
rect 48558 21528 49054 21584
rect 49110 21528 49115 21584
rect 48497 21526 49115 21528
rect 48497 21523 48563 21526
rect 49049 21523 49115 21526
rect 49233 21586 49299 21589
rect 52545 21586 52611 21589
rect 56685 21586 56751 21589
rect 49233 21584 52611 21586
rect 49233 21528 49238 21584
rect 49294 21528 52550 21584
rect 52606 21528 52611 21584
rect 49233 21526 52611 21528
rect 49233 21523 49299 21526
rect 52545 21523 52611 21526
rect 55630 21584 56751 21586
rect 55630 21528 56690 21584
rect 56746 21528 56751 21584
rect 55630 21526 56751 21528
rect 39982 21388 39988 21452
rect 40052 21450 40058 21452
rect 55630 21450 55690 21526
rect 56685 21523 56751 21526
rect 40052 21390 55690 21450
rect 40052 21388 40058 21390
rect 41270 21252 41276 21316
rect 41340 21314 41346 21316
rect 49233 21314 49299 21317
rect 41340 21312 49299 21314
rect 41340 21256 49238 21312
rect 49294 21256 49299 21312
rect 41340 21254 49299 21256
rect 41340 21252 41346 21254
rect 49233 21251 49299 21254
rect 49785 21314 49851 21317
rect 50705 21314 50771 21317
rect 54937 21314 55003 21317
rect 49785 21312 55003 21314
rect 49785 21256 49790 21312
rect 49846 21256 50710 21312
rect 50766 21256 54942 21312
rect 54998 21256 55003 21312
rect 49785 21254 55003 21256
rect 49785 21251 49851 21254
rect 50705 21251 50771 21254
rect 54937 21251 55003 21254
rect 4210 21248 4526 21249
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 34930 21248 35246 21249
rect 34930 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35246 21248
rect 34930 21183 35246 21184
rect 47945 21178 48011 21181
rect 51257 21178 51323 21181
rect 47945 21176 51323 21178
rect 47945 21120 47950 21176
rect 48006 21120 51262 21176
rect 51318 21120 51323 21176
rect 47945 21118 51323 21120
rect 47945 21115 48011 21118
rect 51257 21115 51323 21118
rect 48589 21042 48655 21045
rect 48998 21042 49004 21044
rect 48589 21040 49004 21042
rect 48589 20984 48594 21040
rect 48650 20984 49004 21040
rect 48589 20982 49004 20984
rect 48589 20979 48655 20982
rect 48998 20980 49004 20982
rect 49068 21042 49074 21044
rect 49233 21042 49299 21045
rect 49068 21040 49299 21042
rect 49068 20984 49238 21040
rect 49294 20984 49299 21040
rect 49068 20982 49299 20984
rect 49068 20980 49074 20982
rect 49233 20979 49299 20982
rect 50153 21042 50219 21045
rect 50797 21042 50863 21045
rect 50153 21040 50863 21042
rect 50153 20984 50158 21040
rect 50214 20984 50802 21040
rect 50858 20984 50863 21040
rect 50153 20982 50863 20984
rect 50153 20979 50219 20982
rect 50797 20979 50863 20982
rect 34697 20906 34763 20909
rect 36353 20906 36419 20909
rect 34697 20904 36419 20906
rect 34697 20848 34702 20904
rect 34758 20848 36358 20904
rect 36414 20848 36419 20904
rect 34697 20846 36419 20848
rect 34697 20843 34763 20846
rect 36353 20843 36419 20846
rect 36813 20906 36879 20909
rect 41270 20906 41276 20908
rect 36813 20904 41276 20906
rect 36813 20848 36818 20904
rect 36874 20848 41276 20904
rect 36813 20846 41276 20848
rect 36813 20843 36879 20846
rect 41270 20844 41276 20846
rect 41340 20844 41346 20908
rect 46841 20906 46907 20909
rect 52177 20906 52243 20909
rect 46841 20904 52243 20906
rect 46841 20848 46846 20904
rect 46902 20848 52182 20904
rect 52238 20848 52243 20904
rect 46841 20846 52243 20848
rect 46841 20843 46907 20846
rect 52177 20843 52243 20846
rect 19977 20770 20043 20773
rect 20989 20770 21055 20773
rect 24853 20770 24919 20773
rect 19977 20768 24919 20770
rect 19977 20712 19982 20768
rect 20038 20712 20994 20768
rect 21050 20712 24858 20768
rect 24914 20712 24919 20768
rect 19977 20710 24919 20712
rect 19977 20707 20043 20710
rect 20989 20707 21055 20710
rect 24853 20707 24919 20710
rect 48773 20772 48839 20773
rect 48773 20768 48820 20772
rect 48884 20770 48890 20772
rect 49141 20770 49207 20773
rect 51257 20770 51323 20773
rect 48773 20712 48778 20768
rect 48773 20708 48820 20712
rect 48884 20710 48930 20770
rect 49141 20768 51323 20770
rect 49141 20712 49146 20768
rect 49202 20712 51262 20768
rect 51318 20712 51323 20768
rect 49141 20710 51323 20712
rect 48884 20708 48890 20710
rect 48773 20707 48839 20708
rect 49141 20707 49207 20710
rect 51257 20707 51323 20710
rect 4870 20704 5186 20705
rect 4870 20640 4876 20704
rect 4940 20640 4956 20704
rect 5020 20640 5036 20704
rect 5100 20640 5116 20704
rect 5180 20640 5186 20704
rect 4870 20639 5186 20640
rect 35590 20704 35906 20705
rect 35590 20640 35596 20704
rect 35660 20640 35676 20704
rect 35740 20640 35756 20704
rect 35820 20640 35836 20704
rect 35900 20640 35906 20704
rect 35590 20639 35906 20640
rect 28901 20634 28967 20637
rect 34697 20634 34763 20637
rect 28901 20632 34763 20634
rect 28901 20576 28906 20632
rect 28962 20576 34702 20632
rect 34758 20576 34763 20632
rect 28901 20574 34763 20576
rect 28901 20571 28967 20574
rect 34697 20571 34763 20574
rect 42977 20634 43043 20637
rect 44909 20634 44975 20637
rect 42977 20632 44975 20634
rect 42977 20576 42982 20632
rect 43038 20576 44914 20632
rect 44970 20576 44975 20632
rect 42977 20574 44975 20576
rect 42977 20571 43043 20574
rect 44909 20571 44975 20574
rect 47853 20634 47919 20637
rect 48446 20634 48452 20636
rect 47853 20632 48452 20634
rect 47853 20576 47858 20632
rect 47914 20576 48452 20632
rect 47853 20574 48452 20576
rect 47853 20571 47919 20574
rect 48446 20572 48452 20574
rect 48516 20634 48522 20636
rect 50153 20634 50219 20637
rect 48516 20632 50219 20634
rect 48516 20576 50158 20632
rect 50214 20576 50219 20632
rect 48516 20574 50219 20576
rect 48516 20572 48522 20574
rect 50153 20571 50219 20574
rect 19793 20498 19859 20501
rect 22553 20498 22619 20501
rect 23197 20498 23263 20501
rect 19793 20496 23263 20498
rect 19793 20440 19798 20496
rect 19854 20440 22558 20496
rect 22614 20440 23202 20496
rect 23258 20440 23263 20496
rect 19793 20438 23263 20440
rect 19793 20435 19859 20438
rect 22553 20435 22619 20438
rect 23197 20435 23263 20438
rect 25262 20436 25268 20500
rect 25332 20498 25338 20500
rect 26141 20498 26207 20501
rect 25332 20496 26207 20498
rect 25332 20440 26146 20496
rect 26202 20440 26207 20496
rect 25332 20438 26207 20440
rect 25332 20436 25338 20438
rect 26141 20435 26207 20438
rect 31753 20498 31819 20501
rect 37825 20498 37891 20501
rect 31753 20496 37891 20498
rect 31753 20440 31758 20496
rect 31814 20440 37830 20496
rect 37886 20440 37891 20496
rect 31753 20438 37891 20440
rect 31753 20435 31819 20438
rect 37825 20435 37891 20438
rect 42885 20498 42951 20501
rect 48589 20498 48655 20501
rect 42885 20496 48655 20498
rect 42885 20440 42890 20496
rect 42946 20440 48594 20496
rect 48650 20440 48655 20496
rect 42885 20438 48655 20440
rect 42885 20435 42951 20438
rect 48589 20435 48655 20438
rect 49509 20498 49575 20501
rect 56869 20498 56935 20501
rect 49509 20496 56935 20498
rect 49509 20440 49514 20496
rect 49570 20440 56874 20496
rect 56930 20440 56935 20496
rect 49509 20438 56935 20440
rect 49509 20435 49575 20438
rect 56869 20435 56935 20438
rect 48773 20226 48839 20229
rect 49233 20226 49299 20229
rect 48773 20224 49299 20226
rect 48773 20168 48778 20224
rect 48834 20168 49238 20224
rect 49294 20168 49299 20224
rect 48773 20166 49299 20168
rect 48773 20163 48839 20166
rect 49233 20163 49299 20166
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 34930 20160 35246 20161
rect 34930 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35246 20160
rect 34930 20095 35246 20096
rect 48681 20090 48747 20093
rect 48814 20090 48820 20092
rect 48681 20088 48820 20090
rect 48681 20032 48686 20088
rect 48742 20032 48820 20088
rect 48681 20030 48820 20032
rect 48681 20027 48747 20030
rect 48814 20028 48820 20030
rect 48884 20028 48890 20092
rect 48957 20090 49023 20093
rect 53373 20090 53439 20093
rect 48957 20088 53439 20090
rect 48957 20032 48962 20088
rect 49018 20032 53378 20088
rect 53434 20032 53439 20088
rect 48957 20030 53439 20032
rect 48957 20027 49023 20030
rect 53373 20027 53439 20030
rect 48589 19954 48655 19957
rect 54569 19954 54635 19957
rect 48589 19952 54635 19954
rect 48589 19896 48594 19952
rect 48650 19896 54574 19952
rect 54630 19896 54635 19952
rect 48589 19894 54635 19896
rect 48589 19891 48655 19894
rect 54569 19891 54635 19894
rect 0 19818 800 19848
rect 34513 19818 34579 19821
rect 35617 19818 35683 19821
rect 0 19728 858 19818
rect 34513 19816 35683 19818
rect 34513 19760 34518 19816
rect 34574 19760 35622 19816
rect 35678 19760 35683 19816
rect 34513 19758 35683 19760
rect 34513 19755 34579 19758
rect 35617 19755 35683 19758
rect 48589 19818 48655 19821
rect 49785 19818 49851 19821
rect 48589 19816 49851 19818
rect 48589 19760 48594 19816
rect 48650 19760 49790 19816
rect 49846 19760 49851 19816
rect 48589 19758 49851 19760
rect 48589 19755 48655 19758
rect 49785 19755 49851 19758
rect 58433 19818 58499 19821
rect 59200 19818 60000 19848
rect 58433 19816 60000 19818
rect 58433 19760 58438 19816
rect 58494 19760 60000 19816
rect 58433 19758 60000 19760
rect 58433 19755 58499 19758
rect 59200 19728 60000 19758
rect 798 19685 858 19728
rect 798 19680 907 19685
rect 798 19624 846 19680
rect 902 19624 907 19680
rect 798 19622 907 19624
rect 841 19619 907 19622
rect 49049 19682 49115 19685
rect 49785 19684 49851 19685
rect 49734 19682 49740 19684
rect 49049 19680 49740 19682
rect 49804 19682 49851 19684
rect 49804 19680 49896 19682
rect 49049 19624 49054 19680
rect 49110 19624 49740 19680
rect 49846 19624 49896 19680
rect 49049 19622 49740 19624
rect 49049 19619 49115 19622
rect 49734 19620 49740 19622
rect 49804 19622 49896 19624
rect 49804 19620 49851 19622
rect 49785 19619 49851 19620
rect 4870 19616 5186 19617
rect 4870 19552 4876 19616
rect 4940 19552 4956 19616
rect 5020 19552 5036 19616
rect 5100 19552 5116 19616
rect 5180 19552 5186 19616
rect 4870 19551 5186 19552
rect 35590 19616 35906 19617
rect 35590 19552 35596 19616
rect 35660 19552 35676 19616
rect 35740 19552 35756 19616
rect 35820 19552 35836 19616
rect 35900 19552 35906 19616
rect 35590 19551 35906 19552
rect 48313 19546 48379 19549
rect 49182 19546 49188 19548
rect 48313 19544 49188 19546
rect 48313 19488 48318 19544
rect 48374 19488 49188 19544
rect 48313 19486 49188 19488
rect 48313 19483 48379 19486
rect 49182 19484 49188 19486
rect 49252 19484 49258 19548
rect 46933 19410 46999 19413
rect 46798 19408 46999 19410
rect 46798 19352 46938 19408
rect 46994 19352 46999 19408
rect 46798 19350 46999 19352
rect 25446 19212 25452 19276
rect 25516 19274 25522 19276
rect 25589 19274 25655 19277
rect 25516 19272 25655 19274
rect 25516 19216 25594 19272
rect 25650 19216 25655 19272
rect 25516 19214 25655 19216
rect 25516 19212 25522 19214
rect 25589 19211 25655 19214
rect 26969 19274 27035 19277
rect 29821 19274 29887 19277
rect 26969 19272 29887 19274
rect 26969 19216 26974 19272
rect 27030 19216 29826 19272
rect 29882 19216 29887 19272
rect 26969 19214 29887 19216
rect 26969 19211 27035 19214
rect 29821 19211 29887 19214
rect 46657 19274 46723 19277
rect 46798 19274 46858 19350
rect 46933 19347 46999 19350
rect 46657 19272 46858 19274
rect 46657 19216 46662 19272
rect 46718 19216 46858 19272
rect 46657 19214 46858 19216
rect 46657 19211 46723 19214
rect 48630 19212 48636 19276
rect 48700 19274 48706 19276
rect 49233 19274 49299 19277
rect 48700 19272 49299 19274
rect 48700 19216 49238 19272
rect 49294 19216 49299 19272
rect 48700 19214 49299 19216
rect 48700 19212 48706 19214
rect 49233 19211 49299 19214
rect 24577 19138 24643 19141
rect 24853 19138 24919 19141
rect 25865 19138 25931 19141
rect 24577 19136 25931 19138
rect 24577 19080 24582 19136
rect 24638 19080 24858 19136
rect 24914 19080 25870 19136
rect 25926 19080 25931 19136
rect 24577 19078 25931 19080
rect 24577 19075 24643 19078
rect 24853 19075 24919 19078
rect 25865 19075 25931 19078
rect 26509 19138 26575 19141
rect 34789 19138 34855 19141
rect 26509 19136 34855 19138
rect 26509 19080 26514 19136
rect 26570 19080 34794 19136
rect 34850 19080 34855 19136
rect 26509 19078 34855 19080
rect 26509 19075 26575 19078
rect 34789 19075 34855 19078
rect 57881 19138 57947 19141
rect 59200 19138 60000 19168
rect 57881 19136 60000 19138
rect 57881 19080 57886 19136
rect 57942 19080 60000 19136
rect 57881 19078 60000 19080
rect 57881 19075 57947 19078
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 34930 19072 35246 19073
rect 34930 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35246 19072
rect 59200 19048 60000 19078
rect 34930 19007 35246 19008
rect 25129 19002 25195 19005
rect 26601 19002 26667 19005
rect 25129 19000 26667 19002
rect 25129 18944 25134 19000
rect 25190 18944 26606 19000
rect 26662 18944 26667 19000
rect 25129 18942 26667 18944
rect 25129 18939 25195 18942
rect 26601 18939 26667 18942
rect 26969 19002 27035 19005
rect 27245 19002 27311 19005
rect 26969 19000 27311 19002
rect 26969 18944 26974 19000
rect 27030 18944 27250 19000
rect 27306 18944 27311 19000
rect 26969 18942 27311 18944
rect 26969 18939 27035 18942
rect 27245 18939 27311 18942
rect 20069 18866 20135 18869
rect 22921 18866 22987 18869
rect 26417 18866 26483 18869
rect 27337 18866 27403 18869
rect 20069 18864 27403 18866
rect 20069 18808 20074 18864
rect 20130 18808 22926 18864
rect 22982 18808 26422 18864
rect 26478 18808 27342 18864
rect 27398 18808 27403 18864
rect 20069 18806 27403 18808
rect 20069 18803 20135 18806
rect 22921 18803 22987 18806
rect 26417 18803 26483 18806
rect 27337 18803 27403 18806
rect 19793 18730 19859 18733
rect 26141 18730 26207 18733
rect 26969 18730 27035 18733
rect 19793 18728 27035 18730
rect 19793 18672 19798 18728
rect 19854 18672 26146 18728
rect 26202 18672 26974 18728
rect 27030 18672 27035 18728
rect 19793 18670 27035 18672
rect 19793 18667 19859 18670
rect 26141 18667 26207 18670
rect 26969 18667 27035 18670
rect 37089 18730 37155 18733
rect 45553 18730 45619 18733
rect 37089 18728 45619 18730
rect 37089 18672 37094 18728
rect 37150 18672 45558 18728
rect 45614 18672 45619 18728
rect 37089 18670 45619 18672
rect 37089 18667 37155 18670
rect 45553 18667 45619 18670
rect 25405 18594 25471 18597
rect 26785 18594 26851 18597
rect 36813 18596 36879 18597
rect 36813 18594 36860 18596
rect 25405 18592 26851 18594
rect 25405 18536 25410 18592
rect 25466 18536 26790 18592
rect 26846 18536 26851 18592
rect 25405 18534 26851 18536
rect 36768 18592 36860 18594
rect 36768 18536 36818 18592
rect 36768 18534 36860 18536
rect 25405 18531 25471 18534
rect 26785 18531 26851 18534
rect 36813 18532 36860 18534
rect 36924 18532 36930 18596
rect 36813 18531 36879 18532
rect 4870 18528 5186 18529
rect 4870 18464 4876 18528
rect 4940 18464 4956 18528
rect 5020 18464 5036 18528
rect 5100 18464 5116 18528
rect 5180 18464 5186 18528
rect 4870 18463 5186 18464
rect 35590 18528 35906 18529
rect 35590 18464 35596 18528
rect 35660 18464 35676 18528
rect 35740 18464 35756 18528
rect 35820 18464 35836 18528
rect 35900 18464 35906 18528
rect 35590 18463 35906 18464
rect 20529 18322 20595 18325
rect 22461 18322 22527 18325
rect 20529 18320 22527 18322
rect 20529 18264 20534 18320
rect 20590 18264 22466 18320
rect 22522 18264 22527 18320
rect 20529 18262 22527 18264
rect 20529 18259 20595 18262
rect 22461 18259 22527 18262
rect 31845 18322 31911 18325
rect 38009 18322 38075 18325
rect 31845 18320 38075 18322
rect 31845 18264 31850 18320
rect 31906 18264 38014 18320
rect 38070 18264 38075 18320
rect 31845 18262 38075 18264
rect 31845 18259 31911 18262
rect 38009 18259 38075 18262
rect 39205 18322 39271 18325
rect 41597 18322 41663 18325
rect 39205 18320 41663 18322
rect 39205 18264 39210 18320
rect 39266 18264 41602 18320
rect 41658 18264 41663 18320
rect 39205 18262 41663 18264
rect 39205 18259 39271 18262
rect 41597 18259 41663 18262
rect 38929 18186 38995 18189
rect 39113 18186 39179 18189
rect 40953 18186 41019 18189
rect 38929 18184 41019 18186
rect 38929 18128 38934 18184
rect 38990 18128 39118 18184
rect 39174 18128 40958 18184
rect 41014 18128 41019 18184
rect 38929 18126 41019 18128
rect 38929 18123 38995 18126
rect 39113 18123 39179 18126
rect 40953 18123 41019 18126
rect 41137 18052 41203 18053
rect 41086 18050 41092 18052
rect 41046 17990 41092 18050
rect 41156 18048 41203 18052
rect 41198 17992 41203 18048
rect 41086 17988 41092 17990
rect 41156 17988 41203 17992
rect 41137 17987 41203 17988
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 34930 17984 35246 17985
rect 34930 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35246 17984
rect 34930 17919 35246 17920
rect 40861 17914 40927 17917
rect 42701 17914 42767 17917
rect 40861 17912 42767 17914
rect 40861 17856 40866 17912
rect 40922 17856 42706 17912
rect 42762 17856 42767 17912
rect 40861 17854 42767 17856
rect 40861 17851 40927 17854
rect 42701 17851 42767 17854
rect 48405 17914 48471 17917
rect 48773 17914 48839 17917
rect 48405 17912 48839 17914
rect 48405 17856 48410 17912
rect 48466 17856 48778 17912
rect 48834 17856 48839 17912
rect 48405 17854 48839 17856
rect 48405 17851 48471 17854
rect 48773 17851 48839 17854
rect 48221 17778 48287 17781
rect 51165 17778 51231 17781
rect 48221 17776 51231 17778
rect 48221 17720 48226 17776
rect 48282 17720 51170 17776
rect 51226 17720 51231 17776
rect 48221 17718 51231 17720
rect 48221 17715 48287 17718
rect 51165 17715 51231 17718
rect 37089 17642 37155 17645
rect 35390 17640 37155 17642
rect 35390 17584 37094 17640
rect 37150 17584 37155 17640
rect 35390 17582 37155 17584
rect 4870 17440 5186 17441
rect 4870 17376 4876 17440
rect 4940 17376 4956 17440
rect 5020 17376 5036 17440
rect 5100 17376 5116 17440
rect 5180 17376 5186 17440
rect 4870 17375 5186 17376
rect 31017 17370 31083 17373
rect 32397 17370 32463 17373
rect 35390 17370 35450 17582
rect 37089 17579 37155 17582
rect 41137 17642 41203 17645
rect 56777 17642 56843 17645
rect 41137 17640 56843 17642
rect 41137 17584 41142 17640
rect 41198 17584 56782 17640
rect 56838 17584 56843 17640
rect 41137 17582 56843 17584
rect 41137 17579 41203 17582
rect 56777 17579 56843 17582
rect 53373 17506 53439 17509
rect 54201 17506 54267 17509
rect 53373 17504 54267 17506
rect 53373 17448 53378 17504
rect 53434 17448 54206 17504
rect 54262 17448 54267 17504
rect 53373 17446 54267 17448
rect 53373 17443 53439 17446
rect 54201 17443 54267 17446
rect 35590 17440 35906 17441
rect 35590 17376 35596 17440
rect 35660 17376 35676 17440
rect 35740 17376 35756 17440
rect 35820 17376 35836 17440
rect 35900 17376 35906 17440
rect 35590 17375 35906 17376
rect 31017 17368 35450 17370
rect 31017 17312 31022 17368
rect 31078 17312 32402 17368
rect 32458 17312 35450 17368
rect 31017 17310 35450 17312
rect 31017 17307 31083 17310
rect 32397 17307 32463 17310
rect 40718 17308 40724 17372
rect 40788 17370 40794 17372
rect 40861 17370 40927 17373
rect 40788 17368 40927 17370
rect 40788 17312 40866 17368
rect 40922 17312 40927 17368
rect 40788 17310 40927 17312
rect 40788 17308 40794 17310
rect 40861 17307 40927 17310
rect 29913 17234 29979 17237
rect 38745 17234 38811 17237
rect 29913 17232 38811 17234
rect 29913 17176 29918 17232
rect 29974 17176 38750 17232
rect 38806 17176 38811 17232
rect 29913 17174 38811 17176
rect 29913 17171 29979 17174
rect 38745 17171 38811 17174
rect 39757 17234 39823 17237
rect 48773 17234 48839 17237
rect 49969 17234 50035 17237
rect 39757 17232 50035 17234
rect 39757 17176 39762 17232
rect 39818 17176 48778 17232
rect 48834 17176 49974 17232
rect 50030 17176 50035 17232
rect 39757 17174 50035 17176
rect 39757 17171 39823 17174
rect 48773 17171 48839 17174
rect 49969 17171 50035 17174
rect 53741 17234 53807 17237
rect 56685 17234 56751 17237
rect 53741 17232 56751 17234
rect 53741 17176 53746 17232
rect 53802 17176 56690 17232
rect 56746 17176 56751 17232
rect 53741 17174 56751 17176
rect 53741 17171 53807 17174
rect 56685 17171 56751 17174
rect 26325 17098 26391 17101
rect 39614 17098 39620 17100
rect 26325 17096 39620 17098
rect 26325 17040 26330 17096
rect 26386 17040 39620 17096
rect 26325 17038 39620 17040
rect 26325 17035 26391 17038
rect 39614 17036 39620 17038
rect 39684 17036 39690 17100
rect 48497 17098 48563 17101
rect 50429 17098 50495 17101
rect 50797 17098 50863 17101
rect 48497 17096 50863 17098
rect 48497 17040 48502 17096
rect 48558 17040 50434 17096
rect 50490 17040 50802 17096
rect 50858 17040 50863 17096
rect 48497 17038 50863 17040
rect 48497 17035 48563 17038
rect 50429 17035 50495 17038
rect 50797 17035 50863 17038
rect 24669 16962 24735 16965
rect 27797 16962 27863 16965
rect 24669 16960 27863 16962
rect 24669 16904 24674 16960
rect 24730 16904 27802 16960
rect 27858 16904 27863 16960
rect 24669 16902 27863 16904
rect 24669 16899 24735 16902
rect 27797 16899 27863 16902
rect 30741 16962 30807 16965
rect 31845 16962 31911 16965
rect 30741 16960 31911 16962
rect 30741 16904 30746 16960
rect 30802 16904 31850 16960
rect 31906 16904 31911 16960
rect 30741 16902 31911 16904
rect 30741 16899 30807 16902
rect 31845 16899 31911 16902
rect 49049 16962 49115 16965
rect 53005 16962 53071 16965
rect 49049 16960 53071 16962
rect 49049 16904 49054 16960
rect 49110 16904 53010 16960
rect 53066 16904 53071 16960
rect 49049 16902 53071 16904
rect 49049 16899 49115 16902
rect 53005 16899 53071 16902
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 34930 16896 35246 16897
rect 34930 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35246 16896
rect 34930 16831 35246 16832
rect 25313 16826 25379 16829
rect 25446 16826 25452 16828
rect 25313 16824 25452 16826
rect 25313 16768 25318 16824
rect 25374 16768 25452 16824
rect 25313 16766 25452 16768
rect 25313 16763 25379 16766
rect 25446 16764 25452 16766
rect 25516 16764 25522 16828
rect 40217 16826 40283 16829
rect 43161 16826 43227 16829
rect 40217 16824 43227 16826
rect 40217 16768 40222 16824
rect 40278 16768 43166 16824
rect 43222 16768 43227 16824
rect 40217 16766 43227 16768
rect 40217 16763 40283 16766
rect 43161 16763 43227 16766
rect 25037 16690 25103 16693
rect 26417 16690 26483 16693
rect 25037 16688 26483 16690
rect 25037 16632 25042 16688
rect 25098 16632 26422 16688
rect 26478 16632 26483 16688
rect 25037 16630 26483 16632
rect 25037 16627 25103 16630
rect 26417 16627 26483 16630
rect 28901 16690 28967 16693
rect 31017 16690 31083 16693
rect 28901 16688 31083 16690
rect 28901 16632 28906 16688
rect 28962 16632 31022 16688
rect 31078 16632 31083 16688
rect 28901 16630 31083 16632
rect 28901 16627 28967 16630
rect 31017 16627 31083 16630
rect 31385 16690 31451 16693
rect 35801 16690 35867 16693
rect 36077 16690 36143 16693
rect 36813 16690 36879 16693
rect 31385 16688 36879 16690
rect 31385 16632 31390 16688
rect 31446 16632 35806 16688
rect 35862 16632 36082 16688
rect 36138 16632 36818 16688
rect 36874 16632 36879 16688
rect 31385 16630 36879 16632
rect 31385 16627 31451 16630
rect 35801 16627 35867 16630
rect 36077 16627 36143 16630
rect 36813 16627 36879 16630
rect 39205 16690 39271 16693
rect 41505 16690 41571 16693
rect 39205 16688 41571 16690
rect 39205 16632 39210 16688
rect 39266 16632 41510 16688
rect 41566 16632 41571 16688
rect 39205 16630 41571 16632
rect 39205 16627 39271 16630
rect 41505 16627 41571 16630
rect 25037 16554 25103 16557
rect 25262 16554 25268 16556
rect 25037 16552 25268 16554
rect 25037 16496 25042 16552
rect 25098 16496 25268 16552
rect 25037 16494 25268 16496
rect 25037 16491 25103 16494
rect 25262 16492 25268 16494
rect 25332 16492 25338 16556
rect 29453 16554 29519 16557
rect 31017 16554 31083 16557
rect 29453 16552 31083 16554
rect 29453 16496 29458 16552
rect 29514 16496 31022 16552
rect 31078 16496 31083 16552
rect 29453 16494 31083 16496
rect 29453 16491 29519 16494
rect 31017 16491 31083 16494
rect 35433 16554 35499 16557
rect 36997 16554 37063 16557
rect 35433 16552 37063 16554
rect 35433 16496 35438 16552
rect 35494 16496 37002 16552
rect 37058 16496 37063 16552
rect 35433 16494 37063 16496
rect 35433 16491 35499 16494
rect 36997 16491 37063 16494
rect 38745 16554 38811 16557
rect 41137 16554 41203 16557
rect 48221 16554 48287 16557
rect 38745 16552 48287 16554
rect 38745 16496 38750 16552
rect 38806 16496 41142 16552
rect 41198 16496 48226 16552
rect 48282 16496 48287 16552
rect 38745 16494 48287 16496
rect 38745 16491 38811 16494
rect 41137 16491 41203 16494
rect 48221 16491 48287 16494
rect 37273 16418 37339 16421
rect 37273 16416 41430 16418
rect 37273 16360 37278 16416
rect 37334 16360 41430 16416
rect 37273 16358 41430 16360
rect 37273 16355 37339 16358
rect 4870 16352 5186 16353
rect 4870 16288 4876 16352
rect 4940 16288 4956 16352
rect 5020 16288 5036 16352
rect 5100 16288 5116 16352
rect 5180 16288 5186 16352
rect 4870 16287 5186 16288
rect 35590 16352 35906 16353
rect 35590 16288 35596 16352
rect 35660 16288 35676 16352
rect 35740 16288 35756 16352
rect 35820 16288 35836 16352
rect 35900 16288 35906 16352
rect 35590 16287 35906 16288
rect 41370 16146 41430 16358
rect 48589 16284 48655 16285
rect 49693 16284 49759 16285
rect 48589 16282 48636 16284
rect 48544 16280 48636 16282
rect 48544 16224 48594 16280
rect 48544 16222 48636 16224
rect 48589 16220 48636 16222
rect 48700 16220 48706 16284
rect 49693 16282 49740 16284
rect 49648 16280 49740 16282
rect 49648 16224 49698 16280
rect 49648 16222 49740 16224
rect 49693 16220 49740 16222
rect 49804 16220 49810 16284
rect 48589 16219 48655 16220
rect 49693 16219 49759 16220
rect 54753 16146 54819 16149
rect 41370 16144 54819 16146
rect 41370 16088 54758 16144
rect 54814 16088 54819 16144
rect 41370 16086 54819 16088
rect 54753 16083 54819 16086
rect 37457 16010 37523 16013
rect 41270 16010 41276 16012
rect 37457 16008 41276 16010
rect 37457 15952 37462 16008
rect 37518 15952 41276 16008
rect 37457 15950 41276 15952
rect 37457 15947 37523 15950
rect 41270 15948 41276 15950
rect 41340 16010 41346 16012
rect 46105 16010 46171 16013
rect 41340 16008 46171 16010
rect 41340 15952 46110 16008
rect 46166 15952 46171 16008
rect 41340 15950 46171 15952
rect 41340 15948 41346 15950
rect 46105 15947 46171 15950
rect 4210 15808 4526 15809
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 34930 15808 35246 15809
rect 34930 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35246 15808
rect 34930 15743 35246 15744
rect 23289 15602 23355 15605
rect 27705 15602 27771 15605
rect 27981 15602 28047 15605
rect 23289 15600 28047 15602
rect 23289 15544 23294 15600
rect 23350 15544 27710 15600
rect 27766 15544 27986 15600
rect 28042 15544 28047 15600
rect 23289 15542 28047 15544
rect 23289 15539 23355 15542
rect 27705 15539 27771 15542
rect 27981 15539 28047 15542
rect 39941 15602 40007 15605
rect 40677 15602 40743 15605
rect 48037 15602 48103 15605
rect 39941 15600 48103 15602
rect 39941 15544 39946 15600
rect 40002 15544 40682 15600
rect 40738 15544 48042 15600
rect 48098 15544 48103 15600
rect 39941 15542 48103 15544
rect 39941 15539 40007 15542
rect 40677 15539 40743 15542
rect 48037 15539 48103 15542
rect 39849 15466 39915 15469
rect 40953 15466 41019 15469
rect 39849 15464 41019 15466
rect 39849 15408 39854 15464
rect 39910 15408 40958 15464
rect 41014 15408 41019 15464
rect 39849 15406 41019 15408
rect 39849 15403 39915 15406
rect 40953 15403 41019 15406
rect 50797 15466 50863 15469
rect 51625 15466 51691 15469
rect 53557 15466 53623 15469
rect 56317 15466 56383 15469
rect 50797 15464 56383 15466
rect 50797 15408 50802 15464
rect 50858 15408 51630 15464
rect 51686 15408 53562 15464
rect 53618 15408 56322 15464
rect 56378 15408 56383 15464
rect 50797 15406 56383 15408
rect 50797 15403 50863 15406
rect 51625 15403 51691 15406
rect 53557 15403 53623 15406
rect 56317 15403 56383 15406
rect 50613 15330 50679 15333
rect 53189 15330 53255 15333
rect 55673 15330 55739 15333
rect 50613 15328 55739 15330
rect 50613 15272 50618 15328
rect 50674 15272 53194 15328
rect 53250 15272 55678 15328
rect 55734 15272 55739 15328
rect 50613 15270 55739 15272
rect 50613 15267 50679 15270
rect 53189 15267 53255 15270
rect 55673 15267 55739 15270
rect 4870 15264 5186 15265
rect 4870 15200 4876 15264
rect 4940 15200 4956 15264
rect 5020 15200 5036 15264
rect 5100 15200 5116 15264
rect 5180 15200 5186 15264
rect 4870 15199 5186 15200
rect 35590 15264 35906 15265
rect 35590 15200 35596 15264
rect 35660 15200 35676 15264
rect 35740 15200 35756 15264
rect 35820 15200 35836 15264
rect 35900 15200 35906 15264
rect 35590 15199 35906 15200
rect 39665 15194 39731 15197
rect 47209 15194 47275 15197
rect 52361 15194 52427 15197
rect 39665 15192 52427 15194
rect 39665 15136 39670 15192
rect 39726 15136 47214 15192
rect 47270 15136 52366 15192
rect 52422 15136 52427 15192
rect 39665 15134 52427 15136
rect 39665 15131 39731 15134
rect 47209 15131 47275 15134
rect 52361 15131 52427 15134
rect 20345 15058 20411 15061
rect 22829 15058 22895 15061
rect 48497 15058 48563 15061
rect 20345 15056 22895 15058
rect 20345 15000 20350 15056
rect 20406 15000 22834 15056
rect 22890 15000 22895 15056
rect 20345 14998 22895 15000
rect 20345 14995 20411 14998
rect 22829 14995 22895 14998
rect 48270 15056 48563 15058
rect 48270 15000 48502 15056
rect 48558 15000 48563 15056
rect 48270 14998 48563 15000
rect 40309 14922 40375 14925
rect 41137 14922 41203 14925
rect 44081 14922 44147 14925
rect 40309 14920 44147 14922
rect 40309 14864 40314 14920
rect 40370 14864 41142 14920
rect 41198 14864 44086 14920
rect 44142 14864 44147 14920
rect 40309 14862 44147 14864
rect 40309 14859 40375 14862
rect 41137 14859 41203 14862
rect 44081 14859 44147 14862
rect 48270 14786 48330 14998
rect 48497 14995 48563 14998
rect 52821 15058 52887 15061
rect 55029 15058 55095 15061
rect 52821 15056 55095 15058
rect 52821 15000 52826 15056
rect 52882 15000 55034 15056
rect 55090 15000 55095 15056
rect 52821 14998 55095 15000
rect 52821 14995 52887 14998
rect 55029 14995 55095 14998
rect 48405 14922 48471 14925
rect 48681 14922 48747 14925
rect 48405 14920 48747 14922
rect 48405 14864 48410 14920
rect 48466 14864 48686 14920
rect 48742 14864 48747 14920
rect 48405 14862 48747 14864
rect 48405 14859 48471 14862
rect 48681 14859 48747 14862
rect 48497 14786 48563 14789
rect 48270 14784 48563 14786
rect 48270 14728 48502 14784
rect 48558 14728 48563 14784
rect 48270 14726 48563 14728
rect 48497 14723 48563 14726
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 34930 14720 35246 14721
rect 34930 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35246 14720
rect 34930 14655 35246 14656
rect 42057 14650 42123 14653
rect 43805 14650 43871 14653
rect 42057 14648 43871 14650
rect 42057 14592 42062 14648
rect 42118 14592 43810 14648
rect 43866 14592 43871 14648
rect 42057 14590 43871 14592
rect 42057 14587 42123 14590
rect 43805 14587 43871 14590
rect 0 14378 800 14408
rect 1209 14378 1275 14381
rect 0 14376 1275 14378
rect 0 14320 1214 14376
rect 1270 14320 1275 14376
rect 0 14318 1275 14320
rect 0 14288 800 14318
rect 1209 14315 1275 14318
rect 48773 14378 48839 14381
rect 50429 14378 50495 14381
rect 48773 14376 50495 14378
rect 48773 14320 48778 14376
rect 48834 14320 50434 14376
rect 50490 14320 50495 14376
rect 48773 14318 50495 14320
rect 48773 14315 48839 14318
rect 50429 14315 50495 14318
rect 4870 14176 5186 14177
rect 4870 14112 4876 14176
rect 4940 14112 4956 14176
rect 5020 14112 5036 14176
rect 5100 14112 5116 14176
rect 5180 14112 5186 14176
rect 4870 14111 5186 14112
rect 35590 14176 35906 14177
rect 35590 14112 35596 14176
rect 35660 14112 35676 14176
rect 35740 14112 35756 14176
rect 35820 14112 35836 14176
rect 35900 14112 35906 14176
rect 35590 14111 35906 14112
rect 49049 13970 49115 13973
rect 51625 13970 51691 13973
rect 49049 13968 51691 13970
rect 49049 13912 49054 13968
rect 49110 13912 51630 13968
rect 51686 13912 51691 13968
rect 49049 13910 51691 13912
rect 49049 13907 49115 13910
rect 51625 13907 51691 13910
rect 20253 13834 20319 13837
rect 36629 13834 36695 13837
rect 20253 13832 36695 13834
rect 20253 13776 20258 13832
rect 20314 13776 36634 13832
rect 36690 13776 36695 13832
rect 20253 13774 36695 13776
rect 20253 13771 20319 13774
rect 36629 13771 36695 13774
rect 58433 13698 58499 13701
rect 59200 13698 60000 13728
rect 58433 13696 60000 13698
rect 58433 13640 58438 13696
rect 58494 13640 60000 13696
rect 58433 13638 60000 13640
rect 58433 13635 58499 13638
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 34930 13632 35246 13633
rect 34930 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35246 13632
rect 59200 13608 60000 13638
rect 34930 13567 35246 13568
rect 41045 13564 41111 13565
rect 41045 13562 41092 13564
rect 41000 13560 41092 13562
rect 41000 13504 41050 13560
rect 41000 13502 41092 13504
rect 41045 13500 41092 13502
rect 41156 13500 41162 13564
rect 41045 13499 41111 13500
rect 4870 13088 5186 13089
rect 4870 13024 4876 13088
rect 4940 13024 4956 13088
rect 5020 13024 5036 13088
rect 5100 13024 5116 13088
rect 5180 13024 5186 13088
rect 4870 13023 5186 13024
rect 35590 13088 35906 13089
rect 35590 13024 35596 13088
rect 35660 13024 35676 13088
rect 35740 13024 35756 13088
rect 35820 13024 35836 13088
rect 35900 13024 35906 13088
rect 35590 13023 35906 13024
rect 26233 13018 26299 13021
rect 27613 13020 27679 13021
rect 27613 13018 27660 13020
rect 26233 13016 27660 13018
rect 26233 12960 26238 13016
rect 26294 12960 27618 13016
rect 26233 12958 27660 12960
rect 26233 12955 26299 12958
rect 27613 12956 27660 12958
rect 27724 12956 27730 13020
rect 27613 12955 27679 12956
rect 37641 12746 37707 12749
rect 38929 12746 38995 12749
rect 37641 12744 38995 12746
rect 37641 12688 37646 12744
rect 37702 12688 38934 12744
rect 38990 12688 38995 12744
rect 37641 12686 38995 12688
rect 37641 12683 37707 12686
rect 38929 12683 38995 12686
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 34930 12544 35246 12545
rect 34930 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35246 12544
rect 34930 12479 35246 12480
rect 32581 12338 32647 12341
rect 33685 12338 33751 12341
rect 32581 12336 33751 12338
rect 32581 12280 32586 12336
rect 32642 12280 33690 12336
rect 33746 12280 33751 12336
rect 32581 12278 33751 12280
rect 32581 12275 32647 12278
rect 33685 12275 33751 12278
rect 34237 12338 34303 12341
rect 41597 12338 41663 12341
rect 34237 12336 41663 12338
rect 34237 12280 34242 12336
rect 34298 12280 41602 12336
rect 41658 12280 41663 12336
rect 34237 12278 41663 12280
rect 34237 12275 34303 12278
rect 41597 12275 41663 12278
rect 32213 12202 32279 12205
rect 33777 12202 33843 12205
rect 32213 12200 33843 12202
rect 32213 12144 32218 12200
rect 32274 12144 33782 12200
rect 33838 12144 33843 12200
rect 32213 12142 33843 12144
rect 32213 12139 32279 12142
rect 33777 12139 33843 12142
rect 35341 12202 35407 12205
rect 42885 12202 42951 12205
rect 35341 12200 42951 12202
rect 35341 12144 35346 12200
rect 35402 12144 42890 12200
rect 42946 12144 42951 12200
rect 35341 12142 42951 12144
rect 35341 12139 35407 12142
rect 42885 12139 42951 12142
rect 4870 12000 5186 12001
rect 4870 11936 4876 12000
rect 4940 11936 4956 12000
rect 5020 11936 5036 12000
rect 5100 11936 5116 12000
rect 5180 11936 5186 12000
rect 4870 11935 5186 11936
rect 35590 12000 35906 12001
rect 35590 11936 35596 12000
rect 35660 11936 35676 12000
rect 35740 11936 35756 12000
rect 35820 11936 35836 12000
rect 35900 11936 35906 12000
rect 35590 11935 35906 11936
rect 29637 11930 29703 11933
rect 33041 11930 33107 11933
rect 33317 11930 33383 11933
rect 29637 11928 33383 11930
rect 29637 11872 29642 11928
rect 29698 11872 33046 11928
rect 33102 11872 33322 11928
rect 33378 11872 33383 11928
rect 29637 11870 33383 11872
rect 29637 11867 29703 11870
rect 33041 11867 33107 11870
rect 33317 11867 33383 11870
rect 29729 11794 29795 11797
rect 38377 11794 38443 11797
rect 38745 11794 38811 11797
rect 29729 11792 38811 11794
rect 29729 11736 29734 11792
rect 29790 11736 38382 11792
rect 38438 11736 38750 11792
rect 38806 11736 38811 11792
rect 29729 11734 38811 11736
rect 29729 11731 29795 11734
rect 38377 11731 38443 11734
rect 38745 11731 38811 11734
rect 29269 11658 29335 11661
rect 34605 11658 34671 11661
rect 29269 11656 34671 11658
rect 29269 11600 29274 11656
rect 29330 11600 34610 11656
rect 34666 11600 34671 11656
rect 29269 11598 34671 11600
rect 29269 11595 29335 11598
rect 34605 11595 34671 11598
rect 35065 11658 35131 11661
rect 35065 11656 35404 11658
rect 35065 11600 35070 11656
rect 35126 11600 35404 11656
rect 35065 11598 35404 11600
rect 35065 11595 35131 11598
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 34930 11456 35246 11457
rect 34930 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35246 11456
rect 34930 11391 35246 11392
rect 29085 11250 29151 11253
rect 30925 11250 30991 11253
rect 29085 11248 30991 11250
rect 29085 11192 29090 11248
rect 29146 11192 30930 11248
rect 30986 11192 30991 11248
rect 29085 11190 30991 11192
rect 29085 11187 29151 11190
rect 30925 11187 30991 11190
rect 35065 11250 35131 11253
rect 35344 11250 35404 11598
rect 35065 11248 35404 11250
rect 35065 11192 35070 11248
rect 35126 11192 35404 11248
rect 35065 11190 35404 11192
rect 37457 11250 37523 11253
rect 38837 11250 38903 11253
rect 39205 11250 39271 11253
rect 39941 11250 40007 11253
rect 37457 11248 40007 11250
rect 37457 11192 37462 11248
rect 37518 11192 38842 11248
rect 38898 11192 39210 11248
rect 39266 11192 39946 11248
rect 40002 11192 40007 11248
rect 37457 11190 40007 11192
rect 35065 11187 35131 11190
rect 37457 11187 37523 11190
rect 38837 11187 38903 11190
rect 39205 11187 39271 11190
rect 39941 11187 40007 11190
rect 26693 11114 26759 11117
rect 35341 11114 35407 11117
rect 38193 11114 38259 11117
rect 26693 11112 38259 11114
rect 26693 11056 26698 11112
rect 26754 11056 35346 11112
rect 35402 11056 38198 11112
rect 38254 11056 38259 11112
rect 26693 11054 38259 11056
rect 26693 11051 26759 11054
rect 35341 11051 35407 11054
rect 38193 11051 38259 11054
rect 28993 10978 29059 10981
rect 31017 10978 31083 10981
rect 28993 10976 31083 10978
rect 28993 10920 28998 10976
rect 29054 10920 31022 10976
rect 31078 10920 31083 10976
rect 28993 10918 31083 10920
rect 28993 10915 29059 10918
rect 31017 10915 31083 10918
rect 4870 10912 5186 10913
rect 4870 10848 4876 10912
rect 4940 10848 4956 10912
rect 5020 10848 5036 10912
rect 5100 10848 5116 10912
rect 5180 10848 5186 10912
rect 4870 10847 5186 10848
rect 35590 10912 35906 10913
rect 35590 10848 35596 10912
rect 35660 10848 35676 10912
rect 35740 10848 35756 10912
rect 35820 10848 35836 10912
rect 35900 10848 35906 10912
rect 35590 10847 35906 10848
rect 32397 10706 32463 10709
rect 35065 10706 35131 10709
rect 32397 10704 35131 10706
rect 32397 10648 32402 10704
rect 32458 10648 35070 10704
rect 35126 10648 35131 10704
rect 32397 10646 35131 10648
rect 32397 10643 32463 10646
rect 35065 10643 35131 10646
rect 32305 10570 32371 10573
rect 35893 10570 35959 10573
rect 36353 10570 36419 10573
rect 32305 10568 36419 10570
rect 32305 10512 32310 10568
rect 32366 10512 35898 10568
rect 35954 10512 36358 10568
rect 36414 10512 36419 10568
rect 32305 10510 36419 10512
rect 32305 10507 32371 10510
rect 35893 10507 35959 10510
rect 36353 10507 36419 10510
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 34930 10368 35246 10369
rect 34930 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35246 10368
rect 34930 10303 35246 10304
rect 31845 10162 31911 10165
rect 32305 10162 32371 10165
rect 32489 10162 32555 10165
rect 33593 10162 33659 10165
rect 31845 10160 33659 10162
rect 31845 10104 31850 10160
rect 31906 10104 32310 10160
rect 32366 10104 32494 10160
rect 32550 10104 33598 10160
rect 33654 10104 33659 10160
rect 31845 10102 33659 10104
rect 31845 10099 31911 10102
rect 32305 10099 32371 10102
rect 32489 10099 32555 10102
rect 33593 10099 33659 10102
rect 4870 9824 5186 9825
rect 4870 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5186 9824
rect 4870 9759 5186 9760
rect 35590 9824 35906 9825
rect 35590 9760 35596 9824
rect 35660 9760 35676 9824
rect 35740 9760 35756 9824
rect 35820 9760 35836 9824
rect 35900 9760 35906 9824
rect 35590 9759 35906 9760
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 34930 9280 35246 9281
rect 34930 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35246 9280
rect 34930 9215 35246 9216
rect 4870 8736 5186 8737
rect 4870 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5186 8736
rect 4870 8671 5186 8672
rect 35590 8736 35906 8737
rect 35590 8672 35596 8736
rect 35660 8672 35676 8736
rect 35740 8672 35756 8736
rect 35820 8672 35836 8736
rect 35900 8672 35906 8736
rect 35590 8671 35906 8672
rect 36854 8196 36860 8260
rect 36924 8258 36930 8260
rect 59200 8258 60000 8288
rect 36924 8198 60000 8258
rect 36924 8196 36930 8198
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 34930 8192 35246 8193
rect 34930 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35246 8192
rect 59200 8168 60000 8198
rect 34930 8127 35246 8128
rect 4870 7648 5186 7649
rect 4870 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5186 7648
rect 4870 7583 5186 7584
rect 35590 7648 35906 7649
rect 35590 7584 35596 7648
rect 35660 7584 35676 7648
rect 35740 7584 35756 7648
rect 35820 7584 35836 7648
rect 35900 7584 35906 7648
rect 35590 7583 35906 7584
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 34930 7039 35246 7040
rect 4870 6560 5186 6561
rect 4870 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5186 6560
rect 4870 6495 5186 6496
rect 35590 6560 35906 6561
rect 35590 6496 35596 6560
rect 35660 6496 35676 6560
rect 35740 6496 35756 6560
rect 35820 6496 35836 6560
rect 35900 6496 35906 6560
rect 35590 6495 35906 6496
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 34930 5951 35246 5952
rect 4870 5472 5186 5473
rect 4870 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5186 5472
rect 4870 5407 5186 5408
rect 35590 5472 35906 5473
rect 35590 5408 35596 5472
rect 35660 5408 35676 5472
rect 35740 5408 35756 5472
rect 35820 5408 35836 5472
rect 35900 5408 35906 5472
rect 35590 5407 35906 5408
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 34930 4863 35246 4864
rect 4870 4384 5186 4385
rect 4870 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5186 4384
rect 4870 4319 5186 4320
rect 35590 4384 35906 4385
rect 35590 4320 35596 4384
rect 35660 4320 35676 4384
rect 35740 4320 35756 4384
rect 35820 4320 35836 4384
rect 35900 4320 35906 4384
rect 35590 4319 35906 4320
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 4870 3296 5186 3297
rect 4870 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5186 3296
rect 4870 3231 5186 3232
rect 35590 3296 35906 3297
rect 35590 3232 35596 3296
rect 35660 3232 35676 3296
rect 35740 3232 35756 3296
rect 35820 3232 35836 3296
rect 35900 3232 35906 3296
rect 35590 3231 35906 3232
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 34930 2687 35246 2688
rect 4870 2208 5186 2209
rect 4870 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5186 2208
rect 4870 2143 5186 2144
rect 35590 2208 35906 2209
rect 35590 2144 35596 2208
rect 35660 2144 35676 2208
rect 35740 2144 35756 2208
rect 35820 2144 35836 2208
rect 35900 2144 35906 2208
rect 35590 2143 35906 2144
<< via3 >>
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 4876 37020 4940 37024
rect 4876 36964 4880 37020
rect 4880 36964 4936 37020
rect 4936 36964 4940 37020
rect 4876 36960 4940 36964
rect 4956 37020 5020 37024
rect 4956 36964 4960 37020
rect 4960 36964 5016 37020
rect 5016 36964 5020 37020
rect 4956 36960 5020 36964
rect 5036 37020 5100 37024
rect 5036 36964 5040 37020
rect 5040 36964 5096 37020
rect 5096 36964 5100 37020
rect 5036 36960 5100 36964
rect 5116 37020 5180 37024
rect 5116 36964 5120 37020
rect 5120 36964 5176 37020
rect 5176 36964 5180 37020
rect 5116 36960 5180 36964
rect 35596 37020 35660 37024
rect 35596 36964 35600 37020
rect 35600 36964 35656 37020
rect 35656 36964 35660 37020
rect 35596 36960 35660 36964
rect 35676 37020 35740 37024
rect 35676 36964 35680 37020
rect 35680 36964 35736 37020
rect 35736 36964 35740 37020
rect 35676 36960 35740 36964
rect 35756 37020 35820 37024
rect 35756 36964 35760 37020
rect 35760 36964 35816 37020
rect 35816 36964 35820 37020
rect 35756 36960 35820 36964
rect 35836 37020 35900 37024
rect 35836 36964 35840 37020
rect 35840 36964 35896 37020
rect 35896 36964 35900 37020
rect 35836 36960 35900 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 4876 35932 4940 35936
rect 4876 35876 4880 35932
rect 4880 35876 4936 35932
rect 4936 35876 4940 35932
rect 4876 35872 4940 35876
rect 4956 35932 5020 35936
rect 4956 35876 4960 35932
rect 4960 35876 5016 35932
rect 5016 35876 5020 35932
rect 4956 35872 5020 35876
rect 5036 35932 5100 35936
rect 5036 35876 5040 35932
rect 5040 35876 5096 35932
rect 5096 35876 5100 35932
rect 5036 35872 5100 35876
rect 5116 35932 5180 35936
rect 5116 35876 5120 35932
rect 5120 35876 5176 35932
rect 5176 35876 5180 35932
rect 5116 35872 5180 35876
rect 35596 35932 35660 35936
rect 35596 35876 35600 35932
rect 35600 35876 35656 35932
rect 35656 35876 35660 35932
rect 35596 35872 35660 35876
rect 35676 35932 35740 35936
rect 35676 35876 35680 35932
rect 35680 35876 35736 35932
rect 35736 35876 35740 35932
rect 35676 35872 35740 35876
rect 35756 35932 35820 35936
rect 35756 35876 35760 35932
rect 35760 35876 35816 35932
rect 35816 35876 35820 35932
rect 35756 35872 35820 35876
rect 35836 35932 35900 35936
rect 35836 35876 35840 35932
rect 35840 35876 35896 35932
rect 35896 35876 35900 35932
rect 35836 35872 35900 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 4876 34844 4940 34848
rect 4876 34788 4880 34844
rect 4880 34788 4936 34844
rect 4936 34788 4940 34844
rect 4876 34784 4940 34788
rect 4956 34844 5020 34848
rect 4956 34788 4960 34844
rect 4960 34788 5016 34844
rect 5016 34788 5020 34844
rect 4956 34784 5020 34788
rect 5036 34844 5100 34848
rect 5036 34788 5040 34844
rect 5040 34788 5096 34844
rect 5096 34788 5100 34844
rect 5036 34784 5100 34788
rect 5116 34844 5180 34848
rect 5116 34788 5120 34844
rect 5120 34788 5176 34844
rect 5176 34788 5180 34844
rect 5116 34784 5180 34788
rect 35596 34844 35660 34848
rect 35596 34788 35600 34844
rect 35600 34788 35656 34844
rect 35656 34788 35660 34844
rect 35596 34784 35660 34788
rect 35676 34844 35740 34848
rect 35676 34788 35680 34844
rect 35680 34788 35736 34844
rect 35736 34788 35740 34844
rect 35676 34784 35740 34788
rect 35756 34844 35820 34848
rect 35756 34788 35760 34844
rect 35760 34788 35816 34844
rect 35816 34788 35820 34844
rect 35756 34784 35820 34788
rect 35836 34844 35900 34848
rect 35836 34788 35840 34844
rect 35840 34788 35896 34844
rect 35896 34788 35900 34844
rect 35836 34784 35900 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 4876 33756 4940 33760
rect 4876 33700 4880 33756
rect 4880 33700 4936 33756
rect 4936 33700 4940 33756
rect 4876 33696 4940 33700
rect 4956 33756 5020 33760
rect 4956 33700 4960 33756
rect 4960 33700 5016 33756
rect 5016 33700 5020 33756
rect 4956 33696 5020 33700
rect 5036 33756 5100 33760
rect 5036 33700 5040 33756
rect 5040 33700 5096 33756
rect 5096 33700 5100 33756
rect 5036 33696 5100 33700
rect 5116 33756 5180 33760
rect 5116 33700 5120 33756
rect 5120 33700 5176 33756
rect 5176 33700 5180 33756
rect 5116 33696 5180 33700
rect 35596 33756 35660 33760
rect 35596 33700 35600 33756
rect 35600 33700 35656 33756
rect 35656 33700 35660 33756
rect 35596 33696 35660 33700
rect 35676 33756 35740 33760
rect 35676 33700 35680 33756
rect 35680 33700 35736 33756
rect 35736 33700 35740 33756
rect 35676 33696 35740 33700
rect 35756 33756 35820 33760
rect 35756 33700 35760 33756
rect 35760 33700 35816 33756
rect 35816 33700 35820 33756
rect 35756 33696 35820 33700
rect 35836 33756 35900 33760
rect 35836 33700 35840 33756
rect 35840 33700 35896 33756
rect 35896 33700 35900 33756
rect 35836 33696 35900 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 4876 32668 4940 32672
rect 4876 32612 4880 32668
rect 4880 32612 4936 32668
rect 4936 32612 4940 32668
rect 4876 32608 4940 32612
rect 4956 32668 5020 32672
rect 4956 32612 4960 32668
rect 4960 32612 5016 32668
rect 5016 32612 5020 32668
rect 4956 32608 5020 32612
rect 5036 32668 5100 32672
rect 5036 32612 5040 32668
rect 5040 32612 5096 32668
rect 5096 32612 5100 32668
rect 5036 32608 5100 32612
rect 5116 32668 5180 32672
rect 5116 32612 5120 32668
rect 5120 32612 5176 32668
rect 5176 32612 5180 32668
rect 5116 32608 5180 32612
rect 35596 32668 35660 32672
rect 35596 32612 35600 32668
rect 35600 32612 35656 32668
rect 35656 32612 35660 32668
rect 35596 32608 35660 32612
rect 35676 32668 35740 32672
rect 35676 32612 35680 32668
rect 35680 32612 35736 32668
rect 35736 32612 35740 32668
rect 35676 32608 35740 32612
rect 35756 32668 35820 32672
rect 35756 32612 35760 32668
rect 35760 32612 35816 32668
rect 35816 32612 35820 32668
rect 35756 32608 35820 32612
rect 35836 32668 35900 32672
rect 35836 32612 35840 32668
rect 35840 32612 35896 32668
rect 35896 32612 35900 32668
rect 35836 32608 35900 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 4876 31580 4940 31584
rect 4876 31524 4880 31580
rect 4880 31524 4936 31580
rect 4936 31524 4940 31580
rect 4876 31520 4940 31524
rect 4956 31580 5020 31584
rect 4956 31524 4960 31580
rect 4960 31524 5016 31580
rect 5016 31524 5020 31580
rect 4956 31520 5020 31524
rect 5036 31580 5100 31584
rect 5036 31524 5040 31580
rect 5040 31524 5096 31580
rect 5096 31524 5100 31580
rect 5036 31520 5100 31524
rect 5116 31580 5180 31584
rect 5116 31524 5120 31580
rect 5120 31524 5176 31580
rect 5176 31524 5180 31580
rect 5116 31520 5180 31524
rect 35596 31580 35660 31584
rect 35596 31524 35600 31580
rect 35600 31524 35656 31580
rect 35656 31524 35660 31580
rect 35596 31520 35660 31524
rect 35676 31580 35740 31584
rect 35676 31524 35680 31580
rect 35680 31524 35736 31580
rect 35736 31524 35740 31580
rect 35676 31520 35740 31524
rect 35756 31580 35820 31584
rect 35756 31524 35760 31580
rect 35760 31524 35816 31580
rect 35816 31524 35820 31580
rect 35756 31520 35820 31524
rect 35836 31580 35900 31584
rect 35836 31524 35840 31580
rect 35840 31524 35896 31580
rect 35896 31524 35900 31580
rect 35836 31520 35900 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 4876 30492 4940 30496
rect 4876 30436 4880 30492
rect 4880 30436 4936 30492
rect 4936 30436 4940 30492
rect 4876 30432 4940 30436
rect 4956 30492 5020 30496
rect 4956 30436 4960 30492
rect 4960 30436 5016 30492
rect 5016 30436 5020 30492
rect 4956 30432 5020 30436
rect 5036 30492 5100 30496
rect 5036 30436 5040 30492
rect 5040 30436 5096 30492
rect 5096 30436 5100 30492
rect 5036 30432 5100 30436
rect 5116 30492 5180 30496
rect 5116 30436 5120 30492
rect 5120 30436 5176 30492
rect 5176 30436 5180 30492
rect 5116 30432 5180 30436
rect 35596 30492 35660 30496
rect 35596 30436 35600 30492
rect 35600 30436 35656 30492
rect 35656 30436 35660 30492
rect 35596 30432 35660 30436
rect 35676 30492 35740 30496
rect 35676 30436 35680 30492
rect 35680 30436 35736 30492
rect 35736 30436 35740 30492
rect 35676 30432 35740 30436
rect 35756 30492 35820 30496
rect 35756 30436 35760 30492
rect 35760 30436 35816 30492
rect 35816 30436 35820 30492
rect 35756 30432 35820 30436
rect 35836 30492 35900 30496
rect 35836 30436 35840 30492
rect 35840 30436 35896 30492
rect 35896 30436 35900 30492
rect 35836 30432 35900 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 4876 29404 4940 29408
rect 4876 29348 4880 29404
rect 4880 29348 4936 29404
rect 4936 29348 4940 29404
rect 4876 29344 4940 29348
rect 4956 29404 5020 29408
rect 4956 29348 4960 29404
rect 4960 29348 5016 29404
rect 5016 29348 5020 29404
rect 4956 29344 5020 29348
rect 5036 29404 5100 29408
rect 5036 29348 5040 29404
rect 5040 29348 5096 29404
rect 5096 29348 5100 29404
rect 5036 29344 5100 29348
rect 5116 29404 5180 29408
rect 5116 29348 5120 29404
rect 5120 29348 5176 29404
rect 5176 29348 5180 29404
rect 5116 29344 5180 29348
rect 35596 29404 35660 29408
rect 35596 29348 35600 29404
rect 35600 29348 35656 29404
rect 35656 29348 35660 29404
rect 35596 29344 35660 29348
rect 35676 29404 35740 29408
rect 35676 29348 35680 29404
rect 35680 29348 35736 29404
rect 35736 29348 35740 29404
rect 35676 29344 35740 29348
rect 35756 29404 35820 29408
rect 35756 29348 35760 29404
rect 35760 29348 35816 29404
rect 35816 29348 35820 29404
rect 35756 29344 35820 29348
rect 35836 29404 35900 29408
rect 35836 29348 35840 29404
rect 35840 29348 35896 29404
rect 35896 29348 35900 29404
rect 35836 29344 35900 29348
rect 28028 29064 28092 29068
rect 28028 29008 28078 29064
rect 28078 29008 28092 29064
rect 28028 29004 28092 29008
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 4876 28316 4940 28320
rect 4876 28260 4880 28316
rect 4880 28260 4936 28316
rect 4936 28260 4940 28316
rect 4876 28256 4940 28260
rect 4956 28316 5020 28320
rect 4956 28260 4960 28316
rect 4960 28260 5016 28316
rect 5016 28260 5020 28316
rect 4956 28256 5020 28260
rect 5036 28316 5100 28320
rect 5036 28260 5040 28316
rect 5040 28260 5096 28316
rect 5096 28260 5100 28316
rect 5036 28256 5100 28260
rect 5116 28316 5180 28320
rect 5116 28260 5120 28316
rect 5120 28260 5176 28316
rect 5176 28260 5180 28316
rect 5116 28256 5180 28260
rect 35596 28316 35660 28320
rect 35596 28260 35600 28316
rect 35600 28260 35656 28316
rect 35656 28260 35660 28316
rect 35596 28256 35660 28260
rect 35676 28316 35740 28320
rect 35676 28260 35680 28316
rect 35680 28260 35736 28316
rect 35736 28260 35740 28316
rect 35676 28256 35740 28260
rect 35756 28316 35820 28320
rect 35756 28260 35760 28316
rect 35760 28260 35816 28316
rect 35816 28260 35820 28316
rect 35756 28256 35820 28260
rect 35836 28316 35900 28320
rect 35836 28260 35840 28316
rect 35840 28260 35896 28316
rect 35896 28260 35900 28316
rect 35836 28256 35900 28260
rect 39988 28188 40052 28252
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 4876 27228 4940 27232
rect 4876 27172 4880 27228
rect 4880 27172 4936 27228
rect 4936 27172 4940 27228
rect 4876 27168 4940 27172
rect 4956 27228 5020 27232
rect 4956 27172 4960 27228
rect 4960 27172 5016 27228
rect 5016 27172 5020 27228
rect 4956 27168 5020 27172
rect 5036 27228 5100 27232
rect 5036 27172 5040 27228
rect 5040 27172 5096 27228
rect 5096 27172 5100 27228
rect 5036 27168 5100 27172
rect 5116 27228 5180 27232
rect 5116 27172 5120 27228
rect 5120 27172 5176 27228
rect 5176 27172 5180 27228
rect 5116 27168 5180 27172
rect 35596 27228 35660 27232
rect 35596 27172 35600 27228
rect 35600 27172 35656 27228
rect 35656 27172 35660 27228
rect 35596 27168 35660 27172
rect 35676 27228 35740 27232
rect 35676 27172 35680 27228
rect 35680 27172 35736 27228
rect 35736 27172 35740 27228
rect 35676 27168 35740 27172
rect 35756 27228 35820 27232
rect 35756 27172 35760 27228
rect 35760 27172 35816 27228
rect 35816 27172 35820 27228
rect 35756 27168 35820 27172
rect 35836 27228 35900 27232
rect 35836 27172 35840 27228
rect 35840 27172 35896 27228
rect 35896 27172 35900 27228
rect 35836 27168 35900 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 4876 26140 4940 26144
rect 4876 26084 4880 26140
rect 4880 26084 4936 26140
rect 4936 26084 4940 26140
rect 4876 26080 4940 26084
rect 4956 26140 5020 26144
rect 4956 26084 4960 26140
rect 4960 26084 5016 26140
rect 5016 26084 5020 26140
rect 4956 26080 5020 26084
rect 5036 26140 5100 26144
rect 5036 26084 5040 26140
rect 5040 26084 5096 26140
rect 5096 26084 5100 26140
rect 5036 26080 5100 26084
rect 5116 26140 5180 26144
rect 5116 26084 5120 26140
rect 5120 26084 5176 26140
rect 5176 26084 5180 26140
rect 5116 26080 5180 26084
rect 35596 26140 35660 26144
rect 35596 26084 35600 26140
rect 35600 26084 35656 26140
rect 35656 26084 35660 26140
rect 35596 26080 35660 26084
rect 35676 26140 35740 26144
rect 35676 26084 35680 26140
rect 35680 26084 35736 26140
rect 35736 26084 35740 26140
rect 35676 26080 35740 26084
rect 35756 26140 35820 26144
rect 35756 26084 35760 26140
rect 35760 26084 35816 26140
rect 35816 26084 35820 26140
rect 35756 26080 35820 26084
rect 35836 26140 35900 26144
rect 35836 26084 35840 26140
rect 35840 26084 35896 26140
rect 35896 26084 35900 26140
rect 35836 26080 35900 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 36124 25120 36188 25124
rect 36124 25064 36138 25120
rect 36138 25064 36188 25120
rect 36124 25060 36188 25064
rect 49740 25196 49804 25260
rect 4876 25052 4940 25056
rect 4876 24996 4880 25052
rect 4880 24996 4936 25052
rect 4936 24996 4940 25052
rect 4876 24992 4940 24996
rect 4956 25052 5020 25056
rect 4956 24996 4960 25052
rect 4960 24996 5016 25052
rect 5016 24996 5020 25052
rect 4956 24992 5020 24996
rect 5036 25052 5100 25056
rect 5036 24996 5040 25052
rect 5040 24996 5096 25052
rect 5096 24996 5100 25052
rect 5036 24992 5100 24996
rect 5116 25052 5180 25056
rect 5116 24996 5120 25052
rect 5120 24996 5176 25052
rect 5176 24996 5180 25052
rect 5116 24992 5180 24996
rect 35596 25052 35660 25056
rect 35596 24996 35600 25052
rect 35600 24996 35656 25052
rect 35656 24996 35660 25052
rect 35596 24992 35660 24996
rect 35676 25052 35740 25056
rect 35676 24996 35680 25052
rect 35680 24996 35736 25052
rect 35736 24996 35740 25052
rect 35676 24992 35740 24996
rect 35756 25052 35820 25056
rect 35756 24996 35760 25052
rect 35760 24996 35816 25052
rect 35816 24996 35820 25052
rect 35756 24992 35820 24996
rect 35836 25052 35900 25056
rect 35836 24996 35840 25052
rect 35840 24996 35896 25052
rect 35896 24996 35900 25052
rect 35836 24992 35900 24996
rect 25268 24848 25332 24852
rect 25268 24792 25318 24848
rect 25318 24792 25332 24848
rect 25268 24788 25332 24792
rect 48452 24788 48516 24852
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 4876 23964 4940 23968
rect 4876 23908 4880 23964
rect 4880 23908 4936 23964
rect 4936 23908 4940 23964
rect 4876 23904 4940 23908
rect 4956 23964 5020 23968
rect 4956 23908 4960 23964
rect 4960 23908 5016 23964
rect 5016 23908 5020 23964
rect 4956 23904 5020 23908
rect 5036 23964 5100 23968
rect 5036 23908 5040 23964
rect 5040 23908 5096 23964
rect 5096 23908 5100 23964
rect 5036 23904 5100 23908
rect 5116 23964 5180 23968
rect 5116 23908 5120 23964
rect 5120 23908 5176 23964
rect 5176 23908 5180 23964
rect 5116 23904 5180 23908
rect 35596 23964 35660 23968
rect 35596 23908 35600 23964
rect 35600 23908 35656 23964
rect 35656 23908 35660 23964
rect 35596 23904 35660 23908
rect 35676 23964 35740 23968
rect 35676 23908 35680 23964
rect 35680 23908 35736 23964
rect 35736 23908 35740 23964
rect 35676 23904 35740 23908
rect 35756 23964 35820 23968
rect 35756 23908 35760 23964
rect 35760 23908 35816 23964
rect 35816 23908 35820 23964
rect 35756 23904 35820 23908
rect 35836 23964 35900 23968
rect 35836 23908 35840 23964
rect 35840 23908 35896 23964
rect 35896 23908 35900 23964
rect 35836 23904 35900 23908
rect 40724 23836 40788 23900
rect 27660 23564 27724 23628
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 36124 23080 36188 23084
rect 36124 23024 36174 23080
rect 36174 23024 36188 23080
rect 36124 23020 36188 23024
rect 49004 22944 49068 22948
rect 49004 22888 49018 22944
rect 49018 22888 49068 22944
rect 49004 22884 49068 22888
rect 4876 22876 4940 22880
rect 4876 22820 4880 22876
rect 4880 22820 4936 22876
rect 4936 22820 4940 22876
rect 4876 22816 4940 22820
rect 4956 22876 5020 22880
rect 4956 22820 4960 22876
rect 4960 22820 5016 22876
rect 5016 22820 5020 22876
rect 4956 22816 5020 22820
rect 5036 22876 5100 22880
rect 5036 22820 5040 22876
rect 5040 22820 5096 22876
rect 5096 22820 5100 22876
rect 5036 22816 5100 22820
rect 5116 22876 5180 22880
rect 5116 22820 5120 22876
rect 5120 22820 5176 22876
rect 5176 22820 5180 22876
rect 5116 22816 5180 22820
rect 35596 22876 35660 22880
rect 35596 22820 35600 22876
rect 35600 22820 35656 22876
rect 35656 22820 35660 22876
rect 35596 22816 35660 22820
rect 35676 22876 35740 22880
rect 35676 22820 35680 22876
rect 35680 22820 35736 22876
rect 35736 22820 35740 22876
rect 35676 22816 35740 22820
rect 35756 22876 35820 22880
rect 35756 22820 35760 22876
rect 35760 22820 35816 22876
rect 35816 22820 35820 22876
rect 35756 22816 35820 22820
rect 35836 22876 35900 22880
rect 35836 22820 35840 22876
rect 35840 22820 35896 22876
rect 35896 22820 35900 22876
rect 35836 22816 35900 22820
rect 39620 22340 39684 22404
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 28028 21932 28092 21996
rect 4876 21788 4940 21792
rect 4876 21732 4880 21788
rect 4880 21732 4936 21788
rect 4936 21732 4940 21788
rect 4876 21728 4940 21732
rect 4956 21788 5020 21792
rect 4956 21732 4960 21788
rect 4960 21732 5016 21788
rect 5016 21732 5020 21788
rect 4956 21728 5020 21732
rect 5036 21788 5100 21792
rect 5036 21732 5040 21788
rect 5040 21732 5096 21788
rect 5096 21732 5100 21788
rect 5036 21728 5100 21732
rect 5116 21788 5180 21792
rect 5116 21732 5120 21788
rect 5120 21732 5176 21788
rect 5176 21732 5180 21788
rect 5116 21728 5180 21732
rect 35596 21788 35660 21792
rect 35596 21732 35600 21788
rect 35600 21732 35656 21788
rect 35656 21732 35660 21788
rect 35596 21728 35660 21732
rect 35676 21788 35740 21792
rect 35676 21732 35680 21788
rect 35680 21732 35736 21788
rect 35736 21732 35740 21788
rect 35676 21728 35740 21732
rect 35756 21788 35820 21792
rect 35756 21732 35760 21788
rect 35760 21732 35816 21788
rect 35816 21732 35820 21788
rect 35756 21728 35820 21732
rect 35836 21788 35900 21792
rect 35836 21732 35840 21788
rect 35840 21732 35896 21788
rect 35896 21732 35900 21788
rect 35836 21728 35900 21732
rect 49188 21660 49252 21724
rect 39988 21388 40052 21452
rect 41276 21252 41340 21316
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 49004 20980 49068 21044
rect 41276 20844 41340 20908
rect 48820 20768 48884 20772
rect 48820 20712 48834 20768
rect 48834 20712 48884 20768
rect 48820 20708 48884 20712
rect 4876 20700 4940 20704
rect 4876 20644 4880 20700
rect 4880 20644 4936 20700
rect 4936 20644 4940 20700
rect 4876 20640 4940 20644
rect 4956 20700 5020 20704
rect 4956 20644 4960 20700
rect 4960 20644 5016 20700
rect 5016 20644 5020 20700
rect 4956 20640 5020 20644
rect 5036 20700 5100 20704
rect 5036 20644 5040 20700
rect 5040 20644 5096 20700
rect 5096 20644 5100 20700
rect 5036 20640 5100 20644
rect 5116 20700 5180 20704
rect 5116 20644 5120 20700
rect 5120 20644 5176 20700
rect 5176 20644 5180 20700
rect 5116 20640 5180 20644
rect 35596 20700 35660 20704
rect 35596 20644 35600 20700
rect 35600 20644 35656 20700
rect 35656 20644 35660 20700
rect 35596 20640 35660 20644
rect 35676 20700 35740 20704
rect 35676 20644 35680 20700
rect 35680 20644 35736 20700
rect 35736 20644 35740 20700
rect 35676 20640 35740 20644
rect 35756 20700 35820 20704
rect 35756 20644 35760 20700
rect 35760 20644 35816 20700
rect 35816 20644 35820 20700
rect 35756 20640 35820 20644
rect 35836 20700 35900 20704
rect 35836 20644 35840 20700
rect 35840 20644 35896 20700
rect 35896 20644 35900 20700
rect 35836 20640 35900 20644
rect 48452 20572 48516 20636
rect 25268 20436 25332 20500
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 48820 20028 48884 20092
rect 49740 19680 49804 19684
rect 49740 19624 49790 19680
rect 49790 19624 49804 19680
rect 49740 19620 49804 19624
rect 4876 19612 4940 19616
rect 4876 19556 4880 19612
rect 4880 19556 4936 19612
rect 4936 19556 4940 19612
rect 4876 19552 4940 19556
rect 4956 19612 5020 19616
rect 4956 19556 4960 19612
rect 4960 19556 5016 19612
rect 5016 19556 5020 19612
rect 4956 19552 5020 19556
rect 5036 19612 5100 19616
rect 5036 19556 5040 19612
rect 5040 19556 5096 19612
rect 5096 19556 5100 19612
rect 5036 19552 5100 19556
rect 5116 19612 5180 19616
rect 5116 19556 5120 19612
rect 5120 19556 5176 19612
rect 5176 19556 5180 19612
rect 5116 19552 5180 19556
rect 35596 19612 35660 19616
rect 35596 19556 35600 19612
rect 35600 19556 35656 19612
rect 35656 19556 35660 19612
rect 35596 19552 35660 19556
rect 35676 19612 35740 19616
rect 35676 19556 35680 19612
rect 35680 19556 35736 19612
rect 35736 19556 35740 19612
rect 35676 19552 35740 19556
rect 35756 19612 35820 19616
rect 35756 19556 35760 19612
rect 35760 19556 35816 19612
rect 35816 19556 35820 19612
rect 35756 19552 35820 19556
rect 35836 19612 35900 19616
rect 35836 19556 35840 19612
rect 35840 19556 35896 19612
rect 35896 19556 35900 19612
rect 35836 19552 35900 19556
rect 49188 19484 49252 19548
rect 25452 19212 25516 19276
rect 48636 19212 48700 19276
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 36860 18592 36924 18596
rect 36860 18536 36874 18592
rect 36874 18536 36924 18592
rect 36860 18532 36924 18536
rect 4876 18524 4940 18528
rect 4876 18468 4880 18524
rect 4880 18468 4936 18524
rect 4936 18468 4940 18524
rect 4876 18464 4940 18468
rect 4956 18524 5020 18528
rect 4956 18468 4960 18524
rect 4960 18468 5016 18524
rect 5016 18468 5020 18524
rect 4956 18464 5020 18468
rect 5036 18524 5100 18528
rect 5036 18468 5040 18524
rect 5040 18468 5096 18524
rect 5096 18468 5100 18524
rect 5036 18464 5100 18468
rect 5116 18524 5180 18528
rect 5116 18468 5120 18524
rect 5120 18468 5176 18524
rect 5176 18468 5180 18524
rect 5116 18464 5180 18468
rect 35596 18524 35660 18528
rect 35596 18468 35600 18524
rect 35600 18468 35656 18524
rect 35656 18468 35660 18524
rect 35596 18464 35660 18468
rect 35676 18524 35740 18528
rect 35676 18468 35680 18524
rect 35680 18468 35736 18524
rect 35736 18468 35740 18524
rect 35676 18464 35740 18468
rect 35756 18524 35820 18528
rect 35756 18468 35760 18524
rect 35760 18468 35816 18524
rect 35816 18468 35820 18524
rect 35756 18464 35820 18468
rect 35836 18524 35900 18528
rect 35836 18468 35840 18524
rect 35840 18468 35896 18524
rect 35896 18468 35900 18524
rect 35836 18464 35900 18468
rect 41092 18048 41156 18052
rect 41092 17992 41142 18048
rect 41142 17992 41156 18048
rect 41092 17988 41156 17992
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 4876 17436 4940 17440
rect 4876 17380 4880 17436
rect 4880 17380 4936 17436
rect 4936 17380 4940 17436
rect 4876 17376 4940 17380
rect 4956 17436 5020 17440
rect 4956 17380 4960 17436
rect 4960 17380 5016 17436
rect 5016 17380 5020 17436
rect 4956 17376 5020 17380
rect 5036 17436 5100 17440
rect 5036 17380 5040 17436
rect 5040 17380 5096 17436
rect 5096 17380 5100 17436
rect 5036 17376 5100 17380
rect 5116 17436 5180 17440
rect 5116 17380 5120 17436
rect 5120 17380 5176 17436
rect 5176 17380 5180 17436
rect 5116 17376 5180 17380
rect 35596 17436 35660 17440
rect 35596 17380 35600 17436
rect 35600 17380 35656 17436
rect 35656 17380 35660 17436
rect 35596 17376 35660 17380
rect 35676 17436 35740 17440
rect 35676 17380 35680 17436
rect 35680 17380 35736 17436
rect 35736 17380 35740 17436
rect 35676 17376 35740 17380
rect 35756 17436 35820 17440
rect 35756 17380 35760 17436
rect 35760 17380 35816 17436
rect 35816 17380 35820 17436
rect 35756 17376 35820 17380
rect 35836 17436 35900 17440
rect 35836 17380 35840 17436
rect 35840 17380 35896 17436
rect 35896 17380 35900 17436
rect 35836 17376 35900 17380
rect 40724 17308 40788 17372
rect 39620 17036 39684 17100
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 25452 16764 25516 16828
rect 25268 16492 25332 16556
rect 4876 16348 4940 16352
rect 4876 16292 4880 16348
rect 4880 16292 4936 16348
rect 4936 16292 4940 16348
rect 4876 16288 4940 16292
rect 4956 16348 5020 16352
rect 4956 16292 4960 16348
rect 4960 16292 5016 16348
rect 5016 16292 5020 16348
rect 4956 16288 5020 16292
rect 5036 16348 5100 16352
rect 5036 16292 5040 16348
rect 5040 16292 5096 16348
rect 5096 16292 5100 16348
rect 5036 16288 5100 16292
rect 5116 16348 5180 16352
rect 5116 16292 5120 16348
rect 5120 16292 5176 16348
rect 5176 16292 5180 16348
rect 5116 16288 5180 16292
rect 35596 16348 35660 16352
rect 35596 16292 35600 16348
rect 35600 16292 35656 16348
rect 35656 16292 35660 16348
rect 35596 16288 35660 16292
rect 35676 16348 35740 16352
rect 35676 16292 35680 16348
rect 35680 16292 35736 16348
rect 35736 16292 35740 16348
rect 35676 16288 35740 16292
rect 35756 16348 35820 16352
rect 35756 16292 35760 16348
rect 35760 16292 35816 16348
rect 35816 16292 35820 16348
rect 35756 16288 35820 16292
rect 35836 16348 35900 16352
rect 35836 16292 35840 16348
rect 35840 16292 35896 16348
rect 35896 16292 35900 16348
rect 35836 16288 35900 16292
rect 48636 16280 48700 16284
rect 48636 16224 48650 16280
rect 48650 16224 48700 16280
rect 48636 16220 48700 16224
rect 49740 16280 49804 16284
rect 49740 16224 49754 16280
rect 49754 16224 49804 16280
rect 49740 16220 49804 16224
rect 41276 15948 41340 16012
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 4876 15260 4940 15264
rect 4876 15204 4880 15260
rect 4880 15204 4936 15260
rect 4936 15204 4940 15260
rect 4876 15200 4940 15204
rect 4956 15260 5020 15264
rect 4956 15204 4960 15260
rect 4960 15204 5016 15260
rect 5016 15204 5020 15260
rect 4956 15200 5020 15204
rect 5036 15260 5100 15264
rect 5036 15204 5040 15260
rect 5040 15204 5096 15260
rect 5096 15204 5100 15260
rect 5036 15200 5100 15204
rect 5116 15260 5180 15264
rect 5116 15204 5120 15260
rect 5120 15204 5176 15260
rect 5176 15204 5180 15260
rect 5116 15200 5180 15204
rect 35596 15260 35660 15264
rect 35596 15204 35600 15260
rect 35600 15204 35656 15260
rect 35656 15204 35660 15260
rect 35596 15200 35660 15204
rect 35676 15260 35740 15264
rect 35676 15204 35680 15260
rect 35680 15204 35736 15260
rect 35736 15204 35740 15260
rect 35676 15200 35740 15204
rect 35756 15260 35820 15264
rect 35756 15204 35760 15260
rect 35760 15204 35816 15260
rect 35816 15204 35820 15260
rect 35756 15200 35820 15204
rect 35836 15260 35900 15264
rect 35836 15204 35840 15260
rect 35840 15204 35896 15260
rect 35896 15204 35900 15260
rect 35836 15200 35900 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 4876 14172 4940 14176
rect 4876 14116 4880 14172
rect 4880 14116 4936 14172
rect 4936 14116 4940 14172
rect 4876 14112 4940 14116
rect 4956 14172 5020 14176
rect 4956 14116 4960 14172
rect 4960 14116 5016 14172
rect 5016 14116 5020 14172
rect 4956 14112 5020 14116
rect 5036 14172 5100 14176
rect 5036 14116 5040 14172
rect 5040 14116 5096 14172
rect 5096 14116 5100 14172
rect 5036 14112 5100 14116
rect 5116 14172 5180 14176
rect 5116 14116 5120 14172
rect 5120 14116 5176 14172
rect 5176 14116 5180 14172
rect 5116 14112 5180 14116
rect 35596 14172 35660 14176
rect 35596 14116 35600 14172
rect 35600 14116 35656 14172
rect 35656 14116 35660 14172
rect 35596 14112 35660 14116
rect 35676 14172 35740 14176
rect 35676 14116 35680 14172
rect 35680 14116 35736 14172
rect 35736 14116 35740 14172
rect 35676 14112 35740 14116
rect 35756 14172 35820 14176
rect 35756 14116 35760 14172
rect 35760 14116 35816 14172
rect 35816 14116 35820 14172
rect 35756 14112 35820 14116
rect 35836 14172 35900 14176
rect 35836 14116 35840 14172
rect 35840 14116 35896 14172
rect 35896 14116 35900 14172
rect 35836 14112 35900 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 41092 13560 41156 13564
rect 41092 13504 41106 13560
rect 41106 13504 41156 13560
rect 41092 13500 41156 13504
rect 4876 13084 4940 13088
rect 4876 13028 4880 13084
rect 4880 13028 4936 13084
rect 4936 13028 4940 13084
rect 4876 13024 4940 13028
rect 4956 13084 5020 13088
rect 4956 13028 4960 13084
rect 4960 13028 5016 13084
rect 5016 13028 5020 13084
rect 4956 13024 5020 13028
rect 5036 13084 5100 13088
rect 5036 13028 5040 13084
rect 5040 13028 5096 13084
rect 5096 13028 5100 13084
rect 5036 13024 5100 13028
rect 5116 13084 5180 13088
rect 5116 13028 5120 13084
rect 5120 13028 5176 13084
rect 5176 13028 5180 13084
rect 5116 13024 5180 13028
rect 35596 13084 35660 13088
rect 35596 13028 35600 13084
rect 35600 13028 35656 13084
rect 35656 13028 35660 13084
rect 35596 13024 35660 13028
rect 35676 13084 35740 13088
rect 35676 13028 35680 13084
rect 35680 13028 35736 13084
rect 35736 13028 35740 13084
rect 35676 13024 35740 13028
rect 35756 13084 35820 13088
rect 35756 13028 35760 13084
rect 35760 13028 35816 13084
rect 35816 13028 35820 13084
rect 35756 13024 35820 13028
rect 35836 13084 35900 13088
rect 35836 13028 35840 13084
rect 35840 13028 35896 13084
rect 35896 13028 35900 13084
rect 35836 13024 35900 13028
rect 27660 13016 27724 13020
rect 27660 12960 27674 13016
rect 27674 12960 27724 13016
rect 27660 12956 27724 12960
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 4876 11996 4940 12000
rect 4876 11940 4880 11996
rect 4880 11940 4936 11996
rect 4936 11940 4940 11996
rect 4876 11936 4940 11940
rect 4956 11996 5020 12000
rect 4956 11940 4960 11996
rect 4960 11940 5016 11996
rect 5016 11940 5020 11996
rect 4956 11936 5020 11940
rect 5036 11996 5100 12000
rect 5036 11940 5040 11996
rect 5040 11940 5096 11996
rect 5096 11940 5100 11996
rect 5036 11936 5100 11940
rect 5116 11996 5180 12000
rect 5116 11940 5120 11996
rect 5120 11940 5176 11996
rect 5176 11940 5180 11996
rect 5116 11936 5180 11940
rect 35596 11996 35660 12000
rect 35596 11940 35600 11996
rect 35600 11940 35656 11996
rect 35656 11940 35660 11996
rect 35596 11936 35660 11940
rect 35676 11996 35740 12000
rect 35676 11940 35680 11996
rect 35680 11940 35736 11996
rect 35736 11940 35740 11996
rect 35676 11936 35740 11940
rect 35756 11996 35820 12000
rect 35756 11940 35760 11996
rect 35760 11940 35816 11996
rect 35816 11940 35820 11996
rect 35756 11936 35820 11940
rect 35836 11996 35900 12000
rect 35836 11940 35840 11996
rect 35840 11940 35896 11996
rect 35896 11940 35900 11996
rect 35836 11936 35900 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 4876 10908 4940 10912
rect 4876 10852 4880 10908
rect 4880 10852 4936 10908
rect 4936 10852 4940 10908
rect 4876 10848 4940 10852
rect 4956 10908 5020 10912
rect 4956 10852 4960 10908
rect 4960 10852 5016 10908
rect 5016 10852 5020 10908
rect 4956 10848 5020 10852
rect 5036 10908 5100 10912
rect 5036 10852 5040 10908
rect 5040 10852 5096 10908
rect 5096 10852 5100 10908
rect 5036 10848 5100 10852
rect 5116 10908 5180 10912
rect 5116 10852 5120 10908
rect 5120 10852 5176 10908
rect 5176 10852 5180 10908
rect 5116 10848 5180 10852
rect 35596 10908 35660 10912
rect 35596 10852 35600 10908
rect 35600 10852 35656 10908
rect 35656 10852 35660 10908
rect 35596 10848 35660 10852
rect 35676 10908 35740 10912
rect 35676 10852 35680 10908
rect 35680 10852 35736 10908
rect 35736 10852 35740 10908
rect 35676 10848 35740 10852
rect 35756 10908 35820 10912
rect 35756 10852 35760 10908
rect 35760 10852 35816 10908
rect 35816 10852 35820 10908
rect 35756 10848 35820 10852
rect 35836 10908 35900 10912
rect 35836 10852 35840 10908
rect 35840 10852 35896 10908
rect 35896 10852 35900 10908
rect 35836 10848 35900 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 4876 9820 4940 9824
rect 4876 9764 4880 9820
rect 4880 9764 4936 9820
rect 4936 9764 4940 9820
rect 4876 9760 4940 9764
rect 4956 9820 5020 9824
rect 4956 9764 4960 9820
rect 4960 9764 5016 9820
rect 5016 9764 5020 9820
rect 4956 9760 5020 9764
rect 5036 9820 5100 9824
rect 5036 9764 5040 9820
rect 5040 9764 5096 9820
rect 5096 9764 5100 9820
rect 5036 9760 5100 9764
rect 5116 9820 5180 9824
rect 5116 9764 5120 9820
rect 5120 9764 5176 9820
rect 5176 9764 5180 9820
rect 5116 9760 5180 9764
rect 35596 9820 35660 9824
rect 35596 9764 35600 9820
rect 35600 9764 35656 9820
rect 35656 9764 35660 9820
rect 35596 9760 35660 9764
rect 35676 9820 35740 9824
rect 35676 9764 35680 9820
rect 35680 9764 35736 9820
rect 35736 9764 35740 9820
rect 35676 9760 35740 9764
rect 35756 9820 35820 9824
rect 35756 9764 35760 9820
rect 35760 9764 35816 9820
rect 35816 9764 35820 9820
rect 35756 9760 35820 9764
rect 35836 9820 35900 9824
rect 35836 9764 35840 9820
rect 35840 9764 35896 9820
rect 35896 9764 35900 9820
rect 35836 9760 35900 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 4876 8732 4940 8736
rect 4876 8676 4880 8732
rect 4880 8676 4936 8732
rect 4936 8676 4940 8732
rect 4876 8672 4940 8676
rect 4956 8732 5020 8736
rect 4956 8676 4960 8732
rect 4960 8676 5016 8732
rect 5016 8676 5020 8732
rect 4956 8672 5020 8676
rect 5036 8732 5100 8736
rect 5036 8676 5040 8732
rect 5040 8676 5096 8732
rect 5096 8676 5100 8732
rect 5036 8672 5100 8676
rect 5116 8732 5180 8736
rect 5116 8676 5120 8732
rect 5120 8676 5176 8732
rect 5176 8676 5180 8732
rect 5116 8672 5180 8676
rect 35596 8732 35660 8736
rect 35596 8676 35600 8732
rect 35600 8676 35656 8732
rect 35656 8676 35660 8732
rect 35596 8672 35660 8676
rect 35676 8732 35740 8736
rect 35676 8676 35680 8732
rect 35680 8676 35736 8732
rect 35736 8676 35740 8732
rect 35676 8672 35740 8676
rect 35756 8732 35820 8736
rect 35756 8676 35760 8732
rect 35760 8676 35816 8732
rect 35816 8676 35820 8732
rect 35756 8672 35820 8676
rect 35836 8732 35900 8736
rect 35836 8676 35840 8732
rect 35840 8676 35896 8732
rect 35896 8676 35900 8732
rect 35836 8672 35900 8676
rect 36860 8196 36924 8260
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 4876 7644 4940 7648
rect 4876 7588 4880 7644
rect 4880 7588 4936 7644
rect 4936 7588 4940 7644
rect 4876 7584 4940 7588
rect 4956 7644 5020 7648
rect 4956 7588 4960 7644
rect 4960 7588 5016 7644
rect 5016 7588 5020 7644
rect 4956 7584 5020 7588
rect 5036 7644 5100 7648
rect 5036 7588 5040 7644
rect 5040 7588 5096 7644
rect 5096 7588 5100 7644
rect 5036 7584 5100 7588
rect 5116 7644 5180 7648
rect 5116 7588 5120 7644
rect 5120 7588 5176 7644
rect 5176 7588 5180 7644
rect 5116 7584 5180 7588
rect 35596 7644 35660 7648
rect 35596 7588 35600 7644
rect 35600 7588 35656 7644
rect 35656 7588 35660 7644
rect 35596 7584 35660 7588
rect 35676 7644 35740 7648
rect 35676 7588 35680 7644
rect 35680 7588 35736 7644
rect 35736 7588 35740 7644
rect 35676 7584 35740 7588
rect 35756 7644 35820 7648
rect 35756 7588 35760 7644
rect 35760 7588 35816 7644
rect 35816 7588 35820 7644
rect 35756 7584 35820 7588
rect 35836 7644 35900 7648
rect 35836 7588 35840 7644
rect 35840 7588 35896 7644
rect 35896 7588 35900 7644
rect 35836 7584 35900 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 4876 6556 4940 6560
rect 4876 6500 4880 6556
rect 4880 6500 4936 6556
rect 4936 6500 4940 6556
rect 4876 6496 4940 6500
rect 4956 6556 5020 6560
rect 4956 6500 4960 6556
rect 4960 6500 5016 6556
rect 5016 6500 5020 6556
rect 4956 6496 5020 6500
rect 5036 6556 5100 6560
rect 5036 6500 5040 6556
rect 5040 6500 5096 6556
rect 5096 6500 5100 6556
rect 5036 6496 5100 6500
rect 5116 6556 5180 6560
rect 5116 6500 5120 6556
rect 5120 6500 5176 6556
rect 5176 6500 5180 6556
rect 5116 6496 5180 6500
rect 35596 6556 35660 6560
rect 35596 6500 35600 6556
rect 35600 6500 35656 6556
rect 35656 6500 35660 6556
rect 35596 6496 35660 6500
rect 35676 6556 35740 6560
rect 35676 6500 35680 6556
rect 35680 6500 35736 6556
rect 35736 6500 35740 6556
rect 35676 6496 35740 6500
rect 35756 6556 35820 6560
rect 35756 6500 35760 6556
rect 35760 6500 35816 6556
rect 35816 6500 35820 6556
rect 35756 6496 35820 6500
rect 35836 6556 35900 6560
rect 35836 6500 35840 6556
rect 35840 6500 35896 6556
rect 35896 6500 35900 6556
rect 35836 6496 35900 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 4876 5468 4940 5472
rect 4876 5412 4880 5468
rect 4880 5412 4936 5468
rect 4936 5412 4940 5468
rect 4876 5408 4940 5412
rect 4956 5468 5020 5472
rect 4956 5412 4960 5468
rect 4960 5412 5016 5468
rect 5016 5412 5020 5468
rect 4956 5408 5020 5412
rect 5036 5468 5100 5472
rect 5036 5412 5040 5468
rect 5040 5412 5096 5468
rect 5096 5412 5100 5468
rect 5036 5408 5100 5412
rect 5116 5468 5180 5472
rect 5116 5412 5120 5468
rect 5120 5412 5176 5468
rect 5176 5412 5180 5468
rect 5116 5408 5180 5412
rect 35596 5468 35660 5472
rect 35596 5412 35600 5468
rect 35600 5412 35656 5468
rect 35656 5412 35660 5468
rect 35596 5408 35660 5412
rect 35676 5468 35740 5472
rect 35676 5412 35680 5468
rect 35680 5412 35736 5468
rect 35736 5412 35740 5468
rect 35676 5408 35740 5412
rect 35756 5468 35820 5472
rect 35756 5412 35760 5468
rect 35760 5412 35816 5468
rect 35816 5412 35820 5468
rect 35756 5408 35820 5412
rect 35836 5468 35900 5472
rect 35836 5412 35840 5468
rect 35840 5412 35896 5468
rect 35896 5412 35900 5468
rect 35836 5408 35900 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 4876 4380 4940 4384
rect 4876 4324 4880 4380
rect 4880 4324 4936 4380
rect 4936 4324 4940 4380
rect 4876 4320 4940 4324
rect 4956 4380 5020 4384
rect 4956 4324 4960 4380
rect 4960 4324 5016 4380
rect 5016 4324 5020 4380
rect 4956 4320 5020 4324
rect 5036 4380 5100 4384
rect 5036 4324 5040 4380
rect 5040 4324 5096 4380
rect 5096 4324 5100 4380
rect 5036 4320 5100 4324
rect 5116 4380 5180 4384
rect 5116 4324 5120 4380
rect 5120 4324 5176 4380
rect 5176 4324 5180 4380
rect 5116 4320 5180 4324
rect 35596 4380 35660 4384
rect 35596 4324 35600 4380
rect 35600 4324 35656 4380
rect 35656 4324 35660 4380
rect 35596 4320 35660 4324
rect 35676 4380 35740 4384
rect 35676 4324 35680 4380
rect 35680 4324 35736 4380
rect 35736 4324 35740 4380
rect 35676 4320 35740 4324
rect 35756 4380 35820 4384
rect 35756 4324 35760 4380
rect 35760 4324 35816 4380
rect 35816 4324 35820 4380
rect 35756 4320 35820 4324
rect 35836 4380 35900 4384
rect 35836 4324 35840 4380
rect 35840 4324 35896 4380
rect 35896 4324 35900 4380
rect 35836 4320 35900 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 4876 3292 4940 3296
rect 4876 3236 4880 3292
rect 4880 3236 4936 3292
rect 4936 3236 4940 3292
rect 4876 3232 4940 3236
rect 4956 3292 5020 3296
rect 4956 3236 4960 3292
rect 4960 3236 5016 3292
rect 5016 3236 5020 3292
rect 4956 3232 5020 3236
rect 5036 3292 5100 3296
rect 5036 3236 5040 3292
rect 5040 3236 5096 3292
rect 5096 3236 5100 3292
rect 5036 3232 5100 3236
rect 5116 3292 5180 3296
rect 5116 3236 5120 3292
rect 5120 3236 5176 3292
rect 5176 3236 5180 3292
rect 5116 3232 5180 3236
rect 35596 3292 35660 3296
rect 35596 3236 35600 3292
rect 35600 3236 35656 3292
rect 35656 3236 35660 3292
rect 35596 3232 35660 3236
rect 35676 3292 35740 3296
rect 35676 3236 35680 3292
rect 35680 3236 35736 3292
rect 35736 3236 35740 3292
rect 35676 3232 35740 3236
rect 35756 3292 35820 3296
rect 35756 3236 35760 3292
rect 35760 3236 35816 3292
rect 35816 3236 35820 3292
rect 35756 3232 35820 3236
rect 35836 3292 35900 3296
rect 35836 3236 35840 3292
rect 35840 3236 35896 3292
rect 35896 3236 35900 3292
rect 35836 3232 35900 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 4876 2204 4940 2208
rect 4876 2148 4880 2204
rect 4880 2148 4936 2204
rect 4936 2148 4940 2204
rect 4876 2144 4940 2148
rect 4956 2204 5020 2208
rect 4956 2148 4960 2204
rect 4960 2148 5016 2204
rect 5016 2148 5020 2204
rect 4956 2144 5020 2148
rect 5036 2204 5100 2208
rect 5036 2148 5040 2204
rect 5040 2148 5096 2204
rect 5096 2148 5100 2204
rect 5036 2144 5100 2148
rect 5116 2204 5180 2208
rect 5116 2148 5120 2204
rect 5120 2148 5176 2204
rect 5176 2148 5180 2204
rect 5116 2144 5180 2148
rect 35596 2204 35660 2208
rect 35596 2148 35600 2204
rect 35600 2148 35656 2204
rect 35656 2148 35660 2204
rect 35596 2144 35660 2148
rect 35676 2204 35740 2208
rect 35676 2148 35680 2204
rect 35680 2148 35736 2204
rect 35736 2148 35740 2204
rect 35676 2144 35740 2148
rect 35756 2204 35820 2208
rect 35756 2148 35760 2204
rect 35760 2148 35816 2204
rect 35816 2148 35820 2204
rect 35756 2144 35820 2148
rect 35836 2204 35900 2208
rect 35836 2148 35840 2204
rect 35840 2148 35896 2204
rect 35896 2148 35900 2204
rect 35836 2144 35900 2148
<< metal4 >>
rect 4208 37568 4528 37584
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 4868 37024 5188 37584
rect 4868 36960 4876 37024
rect 4940 36960 4956 37024
rect 5020 36960 5036 37024
rect 5100 36960 5116 37024
rect 5180 36960 5188 37024
rect 4868 35936 5188 36960
rect 4868 35872 4876 35936
rect 4940 35872 4956 35936
rect 5020 35872 5036 35936
rect 5100 35872 5116 35936
rect 5180 35872 5188 35936
rect 4868 34848 5188 35872
rect 4868 34784 4876 34848
rect 4940 34784 4956 34848
rect 5020 34784 5036 34848
rect 5100 34784 5116 34848
rect 5180 34784 5188 34848
rect 4868 33760 5188 34784
rect 4868 33696 4876 33760
rect 4940 33696 4956 33760
rect 5020 33696 5036 33760
rect 5100 33696 5116 33760
rect 5180 33696 5188 33760
rect 4868 32672 5188 33696
rect 4868 32608 4876 32672
rect 4940 32608 4956 32672
rect 5020 32608 5036 32672
rect 5100 32608 5116 32672
rect 5180 32608 5188 32672
rect 4868 31584 5188 32608
rect 4868 31520 4876 31584
rect 4940 31520 4956 31584
rect 5020 31520 5036 31584
rect 5100 31520 5116 31584
rect 5180 31520 5188 31584
rect 4868 30496 5188 31520
rect 4868 30432 4876 30496
rect 4940 30432 4956 30496
rect 5020 30432 5036 30496
rect 5100 30432 5116 30496
rect 5180 30432 5188 30496
rect 4868 29408 5188 30432
rect 4868 29344 4876 29408
rect 4940 29344 4956 29408
rect 5020 29344 5036 29408
rect 5100 29344 5116 29408
rect 5180 29344 5188 29408
rect 4868 28320 5188 29344
rect 34928 37568 35248 37584
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 28027 29068 28093 29069
rect 28027 29004 28028 29068
rect 28092 29004 28093 29068
rect 28027 29003 28093 29004
rect 4868 28256 4876 28320
rect 4940 28256 4956 28320
rect 5020 28256 5036 28320
rect 5100 28256 5116 28320
rect 5180 28256 5188 28320
rect 4868 27232 5188 28256
rect 4868 27168 4876 27232
rect 4940 27168 4956 27232
rect 5020 27168 5036 27232
rect 5100 27168 5116 27232
rect 5180 27168 5188 27232
rect 4868 26144 5188 27168
rect 4868 26080 4876 26144
rect 4940 26080 4956 26144
rect 5020 26080 5036 26144
rect 5100 26080 5116 26144
rect 5180 26080 5188 26144
rect 4868 25056 5188 26080
rect 4868 24992 4876 25056
rect 4940 24992 4956 25056
rect 5020 24992 5036 25056
rect 5100 24992 5116 25056
rect 5180 24992 5188 25056
rect 4868 23968 5188 24992
rect 25267 24852 25333 24853
rect 25267 24788 25268 24852
rect 25332 24788 25333 24852
rect 25267 24787 25333 24788
rect 4868 23904 4876 23968
rect 4940 23904 4956 23968
rect 5020 23904 5036 23968
rect 5100 23904 5116 23968
rect 5180 23904 5188 23968
rect 4868 22880 5188 23904
rect 4868 22816 4876 22880
rect 4940 22816 4956 22880
rect 5020 22816 5036 22880
rect 5100 22816 5116 22880
rect 5180 22816 5188 22880
rect 4868 21792 5188 22816
rect 4868 21728 4876 21792
rect 4940 21728 4956 21792
rect 5020 21728 5036 21792
rect 5100 21728 5116 21792
rect 5180 21728 5188 21792
rect 4868 20704 5188 21728
rect 4868 20640 4876 20704
rect 4940 20640 4956 20704
rect 5020 20640 5036 20704
rect 5100 20640 5116 20704
rect 5180 20640 5188 20704
rect 4868 19616 5188 20640
rect 25270 20501 25330 24787
rect 27659 23628 27725 23629
rect 27659 23564 27660 23628
rect 27724 23564 27725 23628
rect 27659 23563 27725 23564
rect 25267 20500 25333 20501
rect 25267 20436 25268 20500
rect 25332 20436 25333 20500
rect 25267 20435 25333 20436
rect 4868 19552 4876 19616
rect 4940 19552 4956 19616
rect 5020 19552 5036 19616
rect 5100 19552 5116 19616
rect 5180 19552 5188 19616
rect 4868 18528 5188 19552
rect 4868 18464 4876 18528
rect 4940 18464 4956 18528
rect 5020 18464 5036 18528
rect 5100 18464 5116 18528
rect 5180 18464 5188 18528
rect 4868 17440 5188 18464
rect 4868 17376 4876 17440
rect 4940 17376 4956 17440
rect 5020 17376 5036 17440
rect 5100 17376 5116 17440
rect 5180 17376 5188 17440
rect 4868 16352 5188 17376
rect 25270 16557 25330 20435
rect 25451 19276 25517 19277
rect 25451 19212 25452 19276
rect 25516 19212 25517 19276
rect 25451 19211 25517 19212
rect 25454 16829 25514 19211
rect 25451 16828 25517 16829
rect 25451 16764 25452 16828
rect 25516 16764 25517 16828
rect 25451 16763 25517 16764
rect 25267 16556 25333 16557
rect 25267 16492 25268 16556
rect 25332 16492 25333 16556
rect 25267 16491 25333 16492
rect 4868 16288 4876 16352
rect 4940 16288 4956 16352
rect 5020 16288 5036 16352
rect 5100 16288 5116 16352
rect 5180 16288 5188 16352
rect 4868 15264 5188 16288
rect 4868 15200 4876 15264
rect 4940 15200 4956 15264
rect 5020 15200 5036 15264
rect 5100 15200 5116 15264
rect 5180 15200 5188 15264
rect 4868 14176 5188 15200
rect 4868 14112 4876 14176
rect 4940 14112 4956 14176
rect 5020 14112 5036 14176
rect 5100 14112 5116 14176
rect 5180 14112 5188 14176
rect 4868 13088 5188 14112
rect 4868 13024 4876 13088
rect 4940 13024 4956 13088
rect 5020 13024 5036 13088
rect 5100 13024 5116 13088
rect 5180 13024 5188 13088
rect 4868 12000 5188 13024
rect 27662 13021 27722 23563
rect 28030 21997 28090 29003
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 28027 21996 28093 21997
rect 28027 21932 28028 21996
rect 28092 21932 28093 21996
rect 28027 21931 28093 21932
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 27659 13020 27725 13021
rect 27659 12956 27660 13020
rect 27724 12956 27725 13020
rect 27659 12955 27725 12956
rect 4868 11936 4876 12000
rect 4940 11936 4956 12000
rect 5020 11936 5036 12000
rect 5100 11936 5116 12000
rect 5180 11936 5188 12000
rect 4868 10912 5188 11936
rect 4868 10848 4876 10912
rect 4940 10848 4956 10912
rect 5020 10848 5036 10912
rect 5100 10848 5116 10912
rect 5180 10848 5188 10912
rect 4868 9824 5188 10848
rect 4868 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5188 9824
rect 4868 8736 5188 9760
rect 4868 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5188 8736
rect 4868 7648 5188 8672
rect 4868 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5188 7648
rect 4868 6560 5188 7584
rect 4868 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5188 6560
rect 4868 5472 5188 6496
rect 4868 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5188 5472
rect 4868 4384 5188 5408
rect 4868 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5188 4384
rect 4868 3296 5188 4320
rect 4868 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5188 3296
rect 4868 2208 5188 3232
rect 4868 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5188 2208
rect 4868 2128 5188 2144
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
rect 35588 37024 35908 37584
rect 35588 36960 35596 37024
rect 35660 36960 35676 37024
rect 35740 36960 35756 37024
rect 35820 36960 35836 37024
rect 35900 36960 35908 37024
rect 35588 35936 35908 36960
rect 35588 35872 35596 35936
rect 35660 35872 35676 35936
rect 35740 35872 35756 35936
rect 35820 35872 35836 35936
rect 35900 35872 35908 35936
rect 35588 34848 35908 35872
rect 35588 34784 35596 34848
rect 35660 34784 35676 34848
rect 35740 34784 35756 34848
rect 35820 34784 35836 34848
rect 35900 34784 35908 34848
rect 35588 33760 35908 34784
rect 35588 33696 35596 33760
rect 35660 33696 35676 33760
rect 35740 33696 35756 33760
rect 35820 33696 35836 33760
rect 35900 33696 35908 33760
rect 35588 32672 35908 33696
rect 35588 32608 35596 32672
rect 35660 32608 35676 32672
rect 35740 32608 35756 32672
rect 35820 32608 35836 32672
rect 35900 32608 35908 32672
rect 35588 31584 35908 32608
rect 35588 31520 35596 31584
rect 35660 31520 35676 31584
rect 35740 31520 35756 31584
rect 35820 31520 35836 31584
rect 35900 31520 35908 31584
rect 35588 30496 35908 31520
rect 35588 30432 35596 30496
rect 35660 30432 35676 30496
rect 35740 30432 35756 30496
rect 35820 30432 35836 30496
rect 35900 30432 35908 30496
rect 35588 29408 35908 30432
rect 35588 29344 35596 29408
rect 35660 29344 35676 29408
rect 35740 29344 35756 29408
rect 35820 29344 35836 29408
rect 35900 29344 35908 29408
rect 35588 28320 35908 29344
rect 35588 28256 35596 28320
rect 35660 28256 35676 28320
rect 35740 28256 35756 28320
rect 35820 28256 35836 28320
rect 35900 28256 35908 28320
rect 35588 27232 35908 28256
rect 39987 28252 40053 28253
rect 39987 28188 39988 28252
rect 40052 28188 40053 28252
rect 39987 28187 40053 28188
rect 35588 27168 35596 27232
rect 35660 27168 35676 27232
rect 35740 27168 35756 27232
rect 35820 27168 35836 27232
rect 35900 27168 35908 27232
rect 35588 26144 35908 27168
rect 35588 26080 35596 26144
rect 35660 26080 35676 26144
rect 35740 26080 35756 26144
rect 35820 26080 35836 26144
rect 35900 26080 35908 26144
rect 35588 25056 35908 26080
rect 36123 25124 36189 25125
rect 36123 25060 36124 25124
rect 36188 25060 36189 25124
rect 36123 25059 36189 25060
rect 35588 24992 35596 25056
rect 35660 24992 35676 25056
rect 35740 24992 35756 25056
rect 35820 24992 35836 25056
rect 35900 24992 35908 25056
rect 35588 23968 35908 24992
rect 35588 23904 35596 23968
rect 35660 23904 35676 23968
rect 35740 23904 35756 23968
rect 35820 23904 35836 23968
rect 35900 23904 35908 23968
rect 35588 22880 35908 23904
rect 36126 23085 36186 25059
rect 36123 23084 36189 23085
rect 36123 23020 36124 23084
rect 36188 23020 36189 23084
rect 36123 23019 36189 23020
rect 35588 22816 35596 22880
rect 35660 22816 35676 22880
rect 35740 22816 35756 22880
rect 35820 22816 35836 22880
rect 35900 22816 35908 22880
rect 35588 21792 35908 22816
rect 39619 22404 39685 22405
rect 39619 22340 39620 22404
rect 39684 22340 39685 22404
rect 39619 22339 39685 22340
rect 35588 21728 35596 21792
rect 35660 21728 35676 21792
rect 35740 21728 35756 21792
rect 35820 21728 35836 21792
rect 35900 21728 35908 21792
rect 35588 20704 35908 21728
rect 35588 20640 35596 20704
rect 35660 20640 35676 20704
rect 35740 20640 35756 20704
rect 35820 20640 35836 20704
rect 35900 20640 35908 20704
rect 35588 19616 35908 20640
rect 35588 19552 35596 19616
rect 35660 19552 35676 19616
rect 35740 19552 35756 19616
rect 35820 19552 35836 19616
rect 35900 19552 35908 19616
rect 35588 18528 35908 19552
rect 36859 18596 36925 18597
rect 36859 18532 36860 18596
rect 36924 18532 36925 18596
rect 36859 18531 36925 18532
rect 35588 18464 35596 18528
rect 35660 18464 35676 18528
rect 35740 18464 35756 18528
rect 35820 18464 35836 18528
rect 35900 18464 35908 18528
rect 35588 17440 35908 18464
rect 35588 17376 35596 17440
rect 35660 17376 35676 17440
rect 35740 17376 35756 17440
rect 35820 17376 35836 17440
rect 35900 17376 35908 17440
rect 35588 16352 35908 17376
rect 35588 16288 35596 16352
rect 35660 16288 35676 16352
rect 35740 16288 35756 16352
rect 35820 16288 35836 16352
rect 35900 16288 35908 16352
rect 35588 15264 35908 16288
rect 35588 15200 35596 15264
rect 35660 15200 35676 15264
rect 35740 15200 35756 15264
rect 35820 15200 35836 15264
rect 35900 15200 35908 15264
rect 35588 14176 35908 15200
rect 35588 14112 35596 14176
rect 35660 14112 35676 14176
rect 35740 14112 35756 14176
rect 35820 14112 35836 14176
rect 35900 14112 35908 14176
rect 35588 13088 35908 14112
rect 35588 13024 35596 13088
rect 35660 13024 35676 13088
rect 35740 13024 35756 13088
rect 35820 13024 35836 13088
rect 35900 13024 35908 13088
rect 35588 12000 35908 13024
rect 35588 11936 35596 12000
rect 35660 11936 35676 12000
rect 35740 11936 35756 12000
rect 35820 11936 35836 12000
rect 35900 11936 35908 12000
rect 35588 10912 35908 11936
rect 35588 10848 35596 10912
rect 35660 10848 35676 10912
rect 35740 10848 35756 10912
rect 35820 10848 35836 10912
rect 35900 10848 35908 10912
rect 35588 9824 35908 10848
rect 35588 9760 35596 9824
rect 35660 9760 35676 9824
rect 35740 9760 35756 9824
rect 35820 9760 35836 9824
rect 35900 9760 35908 9824
rect 35588 8736 35908 9760
rect 35588 8672 35596 8736
rect 35660 8672 35676 8736
rect 35740 8672 35756 8736
rect 35820 8672 35836 8736
rect 35900 8672 35908 8736
rect 35588 7648 35908 8672
rect 36862 8261 36922 18531
rect 39622 17101 39682 22339
rect 39990 21453 40050 28187
rect 49739 25260 49805 25261
rect 49739 25196 49740 25260
rect 49804 25196 49805 25260
rect 49739 25195 49805 25196
rect 48451 24852 48517 24853
rect 48451 24788 48452 24852
rect 48516 24788 48517 24852
rect 48451 24787 48517 24788
rect 40723 23900 40789 23901
rect 40723 23836 40724 23900
rect 40788 23836 40789 23900
rect 40723 23835 40789 23836
rect 39987 21452 40053 21453
rect 39987 21388 39988 21452
rect 40052 21388 40053 21452
rect 39987 21387 40053 21388
rect 40726 17373 40786 23835
rect 41275 21316 41341 21317
rect 41275 21252 41276 21316
rect 41340 21252 41341 21316
rect 41275 21251 41341 21252
rect 41278 20909 41338 21251
rect 41275 20908 41341 20909
rect 41275 20844 41276 20908
rect 41340 20844 41341 20908
rect 41275 20843 41341 20844
rect 41091 18052 41157 18053
rect 41091 17988 41092 18052
rect 41156 17988 41157 18052
rect 41091 17987 41157 17988
rect 40723 17372 40789 17373
rect 40723 17308 40724 17372
rect 40788 17308 40789 17372
rect 40723 17307 40789 17308
rect 39619 17100 39685 17101
rect 39619 17036 39620 17100
rect 39684 17036 39685 17100
rect 39619 17035 39685 17036
rect 41094 13565 41154 17987
rect 41278 16013 41338 20843
rect 48454 20637 48514 24787
rect 49003 22948 49069 22949
rect 49003 22884 49004 22948
rect 49068 22884 49069 22948
rect 49003 22883 49069 22884
rect 49006 21045 49066 22883
rect 49187 21724 49253 21725
rect 49187 21660 49188 21724
rect 49252 21660 49253 21724
rect 49187 21659 49253 21660
rect 49003 21044 49069 21045
rect 49003 20980 49004 21044
rect 49068 20980 49069 21044
rect 49003 20979 49069 20980
rect 48819 20772 48885 20773
rect 48819 20708 48820 20772
rect 48884 20708 48885 20772
rect 48819 20707 48885 20708
rect 48451 20636 48517 20637
rect 48451 20572 48452 20636
rect 48516 20572 48517 20636
rect 48451 20571 48517 20572
rect 48822 20093 48882 20707
rect 48819 20092 48885 20093
rect 48819 20028 48820 20092
rect 48884 20028 48885 20092
rect 48819 20027 48885 20028
rect 49190 19549 49250 21659
rect 49742 19685 49802 25195
rect 49739 19684 49805 19685
rect 49739 19620 49740 19684
rect 49804 19620 49805 19684
rect 49739 19619 49805 19620
rect 49187 19548 49253 19549
rect 49187 19484 49188 19548
rect 49252 19484 49253 19548
rect 49187 19483 49253 19484
rect 48635 19276 48701 19277
rect 48635 19212 48636 19276
rect 48700 19212 48701 19276
rect 48635 19211 48701 19212
rect 48638 16285 48698 19211
rect 49742 16285 49802 19619
rect 48635 16284 48701 16285
rect 48635 16220 48636 16284
rect 48700 16220 48701 16284
rect 48635 16219 48701 16220
rect 49739 16284 49805 16285
rect 49739 16220 49740 16284
rect 49804 16220 49805 16284
rect 49739 16219 49805 16220
rect 41275 16012 41341 16013
rect 41275 15948 41276 16012
rect 41340 15948 41341 16012
rect 41275 15947 41341 15948
rect 41091 13564 41157 13565
rect 41091 13500 41092 13564
rect 41156 13500 41157 13564
rect 41091 13499 41157 13500
rect 36859 8260 36925 8261
rect 36859 8196 36860 8260
rect 36924 8196 36925 8260
rect 36859 8195 36925 8196
rect 35588 7584 35596 7648
rect 35660 7584 35676 7648
rect 35740 7584 35756 7648
rect 35820 7584 35836 7648
rect 35900 7584 35908 7648
rect 35588 6560 35908 7584
rect 35588 6496 35596 6560
rect 35660 6496 35676 6560
rect 35740 6496 35756 6560
rect 35820 6496 35836 6560
rect 35900 6496 35908 6560
rect 35588 5472 35908 6496
rect 35588 5408 35596 5472
rect 35660 5408 35676 5472
rect 35740 5408 35756 5472
rect 35820 5408 35836 5472
rect 35900 5408 35908 5472
rect 35588 4384 35908 5408
rect 35588 4320 35596 4384
rect 35660 4320 35676 4384
rect 35740 4320 35756 4384
rect 35820 4320 35836 4384
rect 35900 4320 35908 4384
rect 35588 3296 35908 4320
rect 35588 3232 35596 3296
rect 35660 3232 35676 3296
rect 35740 3232 35756 3296
rect 35820 3232 35836 3296
rect 35900 3232 35908 3296
rect 35588 2208 35908 3232
rect 35588 2144 35596 2208
rect 35660 2144 35676 2208
rect 35740 2144 35756 2208
rect 35820 2144 35836 2208
rect 35900 2144 35908 2208
rect 35588 2128 35908 2144
use sky130_fd_sc_hd__inv_2  _0722_
timestamp 18001
transform 1 0 27324 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0723_
timestamp 18001
transform -1 0 33212 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0724_
timestamp 18001
transform -1 0 21344 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0725_
timestamp 18001
transform -1 0 42320 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0726_
timestamp 18001
transform -1 0 39836 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0727_
timestamp 18001
transform 1 0 44528 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0728_
timestamp 18001
transform -1 0 42872 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0729_
timestamp 18001
transform -1 0 42688 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0730_
timestamp 18001
transform 1 0 37812 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0731_
timestamp 18001
transform -1 0 38364 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or4b_2  _0732_
timestamp 18001
transform -1 0 32752 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__or4b_2  _0733_
timestamp 18001
transform 1 0 27232 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _0734_
timestamp 18001
transform 1 0 32844 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _0735_
timestamp 18001
transform -1 0 37996 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_1  _0736_
timestamp 18001
transform -1 0 36340 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _0737_
timestamp 18001
transform 1 0 27048 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0738_
timestamp 18001
transform -1 0 31004 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0739_
timestamp 18001
transform 1 0 28520 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0740_
timestamp 18001
transform -1 0 31464 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0741_
timestamp 18001
transform 1 0 30176 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0742_
timestamp 18001
transform 1 0 33396 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0743_
timestamp 18001
transform 1 0 32844 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0744_
timestamp 18001
transform -1 0 34500 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0745_
timestamp 18001
transform -1 0 27692 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0746_
timestamp 18001
transform -1 0 28704 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _0747_
timestamp 18001
transform 1 0 26864 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0748_
timestamp 18001
transform -1 0 27416 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0749_
timestamp 18001
transform 1 0 35144 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nand3_1  _0750_
timestamp 18001
transform 1 0 35420 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0751_
timestamp 18001
transform 1 0 36708 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a41o_1  _0752_
timestamp 18001
transform -1 0 36340 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _0753_
timestamp 18001
transform -1 0 36616 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0754_
timestamp 18001
transform 1 0 36524 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__nor4_2  _0755_
timestamp 18001
transform 1 0 29808 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__inv_2  _0756_
timestamp 18001
transform 1 0 30820 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0757_
timestamp 18001
transform -1 0 23828 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0758_
timestamp 18001
transform -1 0 23460 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0759_
timestamp 18001
transform -1 0 26588 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0760_
timestamp 18001
transform 1 0 25760 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0761_
timestamp 18001
transform 1 0 14720 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or4bb_1  _0762_
timestamp 18001
transform -1 0 20976 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__or4_1  _0763_
timestamp 18001
transform -1 0 18400 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0764_
timestamp 18001
transform 1 0 15088 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0765_
timestamp 18001
transform -1 0 16744 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0766_
timestamp 18001
transform -1 0 20976 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__or4b_2  _0767_
timestamp 18001
transform 1 0 20976 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0768_
timestamp 18001
transform -1 0 19964 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0769_
timestamp 18001
transform -1 0 20516 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or4_2  _0770_
timestamp 18001
transform 1 0 16100 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0771_
timestamp 18001
transform -1 0 16100 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__or4b_2  _0772_
timestamp 18001
transform 1 0 16652 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__nor4_4  _0773_
timestamp 18001
transform -1 0 17940 0 1 7616
box -38 -48 1602 592
use sky130_fd_sc_hd__nor2_1  _0774_
timestamp 18001
transform -1 0 15548 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0775_
timestamp 18001
transform -1 0 16928 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0776_
timestamp 18001
transform 1 0 15824 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0777_
timestamp 18001
transform -1 0 14812 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0778_
timestamp 18001
transform -1 0 14904 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0779_
timestamp 18001
transform -1 0 14352 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0780_
timestamp 18001
transform -1 0 15548 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0781_
timestamp 18001
transform 1 0 13892 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0782_
timestamp 18001
transform -1 0 13064 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0783_
timestamp 18001
transform -1 0 13064 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0784_
timestamp 18001
transform 1 0 15916 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0785_
timestamp 18001
transform -1 0 16100 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_1  _0786_
timestamp 18001
transform 1 0 16100 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__and4_1  _0787_
timestamp 18001
transform 1 0 15916 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0788_
timestamp 18001
transform 1 0 17940 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0789_
timestamp 18001
transform -1 0 17664 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0790_
timestamp 18001
transform -1 0 18584 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0791_
timestamp 18001
transform 1 0 17388 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _0792_
timestamp 18001
transform 1 0 17756 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0793_
timestamp 18001
transform 1 0 18400 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _0794_
timestamp 18001
transform 1 0 20976 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0795_
timestamp 18001
transform 1 0 20332 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0796_
timestamp 18001
transform -1 0 21436 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0797_
timestamp 18001
transform 1 0 21068 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _0798_
timestamp 18001
transform -1 0 20792 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0799_
timestamp 18001
transform 1 0 20976 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0800_
timestamp 18001
transform 1 0 23000 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0801_
timestamp 18001
transform 1 0 21528 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _0802_
timestamp 18001
transform -1 0 20424 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0803_
timestamp 18001
transform 1 0 22264 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0804_
timestamp 18001
transform -1 0 22172 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__and4_1  _0805_
timestamp 18001
transform -1 0 21620 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0806_
timestamp 18001
transform 1 0 21712 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0807_
timestamp 18001
transform -1 0 23276 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0808_
timestamp 18001
transform 1 0 21804 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0809_
timestamp 18001
transform -1 0 21712 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0810_
timestamp 18001
transform 1 0 22172 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _0811_
timestamp 18001
transform 1 0 22632 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0812_
timestamp 18001
transform 1 0 15916 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0813_
timestamp 18001
transform 1 0 16744 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0814_
timestamp 18001
transform -1 0 18860 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__and4_1  _0815_
timestamp 18001
transform -1 0 20516 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0816_
timestamp 18001
transform 1 0 18032 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0817_
timestamp 18001
transform 1 0 12880 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0818_
timestamp 18001
transform -1 0 14444 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0819_
timestamp 18001
transform -1 0 13984 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _0820_
timestamp 18001
transform -1 0 17296 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0821_
timestamp 18001
transform 1 0 14444 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0822_
timestamp 18001
transform -1 0 12880 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0823_
timestamp 18001
transform 1 0 14076 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0824_
timestamp 18001
transform 1 0 14720 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _0825_
timestamp 18001
transform -1 0 15916 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0826_
timestamp 18001
transform -1 0 15088 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0827_
timestamp 18001
transform 1 0 19596 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0828_
timestamp 18001
transform -1 0 19596 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0829_
timestamp 18001
transform -1 0 18860 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _0830_
timestamp 18001
transform -1 0 17388 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0831_
timestamp 18001
transform 1 0 19596 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0832_
timestamp 18001
transform -1 0 17020 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0833_
timestamp 18001
transform -1 0 18676 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__and4_1  _0834_
timestamp 18001
transform -1 0 17848 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0835_
timestamp 18001
transform 1 0 17020 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0836_
timestamp 18001
transform 1 0 12328 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0837_
timestamp 18001
transform -1 0 12972 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0838_
timestamp 18001
transform -1 0 13524 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0839_
timestamp 18001
transform 1 0 12144 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0840_
timestamp 18001
transform 1 0 14720 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0841_
timestamp 18001
transform 1 0 12420 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0842_
timestamp 18001
transform 1 0 14812 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0843_
timestamp 18001
transform -1 0 26772 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0844_
timestamp 18001
transform 1 0 17756 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__or4b_1  _0845_
timestamp 18001
transform -1 0 19964 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _0846_
timestamp 18001
transform 1 0 19228 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0847_
timestamp 18001
transform 1 0 23368 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0848_
timestamp 18001
transform -1 0 25208 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0849_
timestamp 18001
transform 1 0 26956 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0850_
timestamp 18001
transform -1 0 27416 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0851_
timestamp 18001
transform 1 0 23184 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _0852_
timestamp 18001
transform 1 0 23644 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0853_
timestamp 18001
transform -1 0 26588 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0854_
timestamp 18001
transform -1 0 29256 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0855_
timestamp 18001
transform -1 0 29348 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0856_
timestamp 18001
transform -1 0 29072 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0857_
timestamp 18001
transform -1 0 30728 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _0858_
timestamp 18001
transform -1 0 29900 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0859_
timestamp 18001
transform 1 0 28244 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0860_
timestamp 18001
transform 1 0 31740 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0861_
timestamp 18001
transform 1 0 32660 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0862_
timestamp 18001
transform 1 0 32384 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0863_
timestamp 18001
transform 1 0 32108 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0864_
timestamp 18001
transform 1 0 34684 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0865_
timestamp 18001
transform 1 0 33764 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0866_
timestamp 18001
transform 1 0 34040 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0867_
timestamp 18001
transform -1 0 34592 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__or4b_1  _0868_
timestamp 18001
transform 1 0 32752 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__or4b_1  _0869_
timestamp 18001
transform -1 0 35420 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0870_
timestamp 18001
transform -1 0 33856 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__and3_2  _0871_
timestamp 18001
transform -1 0 34132 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_2  _0872_
timestamp 18001
transform 1 0 24380 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0873_
timestamp 18001
transform 1 0 33764 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0874_
timestamp 18001
transform 1 0 33304 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_1  _0875_
timestamp 18001
transform -1 0 33028 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0876_
timestamp 18001
transform 1 0 38640 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0877_
timestamp 18001
transform 1 0 36432 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _0878_
timestamp 18001
transform -1 0 37904 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0879_
timestamp 18001
transform -1 0 38180 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0880_
timestamp 18001
transform -1 0 37168 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _0881_
timestamp 18001
transform 1 0 37076 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0882_
timestamp 18001
transform 1 0 37628 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0883_
timestamp 18001
transform -1 0 37076 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _0884_
timestamp 18001
transform 1 0 36524 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0885_
timestamp 18001
transform -1 0 35052 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0886_
timestamp 18001
transform -1 0 34592 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0887_
timestamp 18001
transform 1 0 36064 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0888_
timestamp 18001
transform -1 0 30728 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0889_
timestamp 18001
transform 1 0 30452 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  _0890_
timestamp 18001
transform -1 0 29440 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0891_
timestamp 18001
transform 1 0 33120 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0892_
timestamp 18001
transform 1 0 33856 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0893_
timestamp 18001
transform -1 0 31004 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0894_
timestamp 18001
transform 1 0 29900 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__a21boi_1  _0895_
timestamp 18001
transform 1 0 33396 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _0896_
timestamp 18001
transform 1 0 33948 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0897_
timestamp 18001
transform 1 0 32292 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0898_
timestamp 18001
transform -1 0 33304 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _0899_
timestamp 18001
transform -1 0 31188 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0900_
timestamp 18001
transform 1 0 30360 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0901_
timestamp 18001
transform 1 0 30912 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0902_
timestamp 18001
transform 1 0 18584 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _0903_
timestamp 18001
transform -1 0 34500 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _0904_
timestamp 18001
transform 1 0 33212 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0905_
timestamp 18001
transform 1 0 31924 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0906_
timestamp 18001
transform 1 0 37168 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__o41a_2  _0907_
timestamp 18001
transform -1 0 37168 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__inv_2  _0908_
timestamp 18001
transform 1 0 37536 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  _0909_
timestamp 18001
transform 1 0 35604 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0910_
timestamp 18001
transform -1 0 37168 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__o32a_1  _0911_
timestamp 18001
transform -1 0 37076 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0912_
timestamp 18001
transform 1 0 38732 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or4b_4  _0913_
timestamp 18001
transform 1 0 32108 0 -1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__nor2_1  _0914_
timestamp 18001
transform -1 0 28060 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0915_
timestamp 18001
transform -1 0 54924 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0916_
timestamp 18001
transform -1 0 37076 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or4b_2  _0917_
timestamp 18001
transform 1 0 31280 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0918_
timestamp 18001
transform -1 0 31096 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0919_
timestamp 18001
transform -1 0 37536 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _0920_
timestamp 18001
transform -1 0 36248 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__and3_2  _0921_
timestamp 18001
transform -1 0 37812 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0922_
timestamp 18001
transform 1 0 32568 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0923_
timestamp 18001
transform -1 0 48484 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _0924_
timestamp 18001
transform 1 0 45356 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0925_
timestamp 18001
transform 1 0 29992 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _0926_
timestamp 18001
transform 1 0 30912 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0927_
timestamp 18001
transform 1 0 27508 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _0928_
timestamp 18001
transform 1 0 28060 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0929_
timestamp 18001
transform -1 0 43056 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _0930_
timestamp 18001
transform 1 0 41124 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0931_
timestamp 18001
transform -1 0 43056 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _0932_
timestamp 18001
transform 1 0 41308 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0933_
timestamp 18001
transform -1 0 36892 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0934_
timestamp 18001
transform -1 0 37260 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0935_
timestamp 18001
transform -1 0 36616 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _0936_
timestamp 18001
transform -1 0 34592 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0937_
timestamp 18001
transform 1 0 40756 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _0938_
timestamp 18001
transform 1 0 42044 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0939_
timestamp 18001
transform 1 0 29900 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0940_
timestamp 18001
transform 1 0 30636 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _0941_
timestamp 18001
transform -1 0 47012 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0942_
timestamp 18001
transform 1 0 46368 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _0943_
timestamp 18001
transform 1 0 30268 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0944_
timestamp 18001
transform 1 0 32108 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0945_
timestamp 18001
transform 1 0 25760 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _0946_
timestamp 18001
transform -1 0 26404 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0947_
timestamp 18001
transform -1 0 45724 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0948_
timestamp 18001
transform 1 0 44344 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0949_
timestamp 18001
transform -1 0 43700 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _0950_
timestamp 18001
transform 1 0 41676 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0951_
timestamp 18001
transform -1 0 35972 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _0952_
timestamp 18001
transform 1 0 34684 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0953_
timestamp 18001
transform -1 0 44344 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _0954_
timestamp 18001
transform 1 0 42504 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0955_
timestamp 18001
transform 1 0 31096 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0956_
timestamp 18001
transform -1 0 31740 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _0957_
timestamp 18001
transform -1 0 47196 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0958_
timestamp 18001
transform 1 0 46368 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0959_
timestamp 18001
transform 1 0 26956 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _0960_
timestamp 18001
transform 1 0 27968 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0961_
timestamp 18001
transform -1 0 24104 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _0962_
timestamp 18001
transform 1 0 22816 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0963_
timestamp 18001
transform 1 0 47564 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _0964_
timestamp 18001
transform -1 0 48944 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0965_
timestamp 18001
transform -1 0 45356 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0966_
timestamp 18001
transform 1 0 44988 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0967_
timestamp 18001
transform 1 0 35052 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _0968_
timestamp 18001
transform 1 0 35144 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0969_
timestamp 18001
transform 1 0 43516 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _0970_
timestamp 18001
transform 1 0 44252 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0971_
timestamp 18001
transform 1 0 29532 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0972_
timestamp 18001
transform -1 0 29900 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0973_
timestamp 18001
transform -1 0 49036 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _0974_
timestamp 18001
transform 1 0 48484 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0975_
timestamp 18001
transform 1 0 25944 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0976_
timestamp 18001
transform 1 0 25944 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0977_
timestamp 18001
transform -1 0 22816 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _0978_
timestamp 18001
transform -1 0 22080 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0979_
timestamp 18001
transform -1 0 47104 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0980_
timestamp 18001
transform 1 0 45908 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _0981_
timestamp 18001
transform -1 0 47104 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0982_
timestamp 18001
transform 1 0 44988 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0983_
timestamp 18001
transform 1 0 35604 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _0984_
timestamp 18001
transform -1 0 36892 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0985_
timestamp 18001
transform -1 0 45080 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _0986_
timestamp 18001
transform 1 0 43792 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0987_
timestamp 18001
transform 1 0 27048 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0988_
timestamp 18001
transform 1 0 27324 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0989_
timestamp 18001
transform -1 0 49680 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _0990_
timestamp 18001
transform 1 0 48852 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0991_
timestamp 18001
transform -1 0 23828 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _0992_
timestamp 18001
transform 1 0 22816 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _0993_
timestamp 18001
transform -1 0 20332 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0994_
timestamp 18001
transform 1 0 18584 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _0995_
timestamp 18001
transform -1 0 48944 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _0996_
timestamp 18001
transform 1 0 46000 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _0997_
timestamp 18001
transform 1 0 48024 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _0998_
timestamp 18001
transform -1 0 49312 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0999_
timestamp 18001
transform -1 0 37168 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1000_
timestamp 18001
transform 1 0 35880 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1001_
timestamp 18001
transform 1 0 42412 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1002_
timestamp 18001
transform 1 0 42780 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1003_
timestamp 18001
transform -1 0 23828 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1004_
timestamp 18001
transform 1 0 22908 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1005_
timestamp 18001
transform 1 0 50232 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1006_
timestamp 18001
transform 1 0 51428 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1007_
timestamp 18001
transform -1 0 22540 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1008_
timestamp 18001
transform 1 0 21804 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1009_
timestamp 18001
transform -1 0 20700 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1010_
timestamp 18001
transform 1 0 19228 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1011_
timestamp 18001
transform -1 0 48944 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1012_
timestamp 18001
transform 1 0 46828 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1013_
timestamp 18001
transform 1 0 48944 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1014_
timestamp 18001
transform 1 0 50140 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1015_
timestamp 18001
transform -1 0 36156 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1016_
timestamp 18001
transform 1 0 35328 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1017_
timestamp 18001
transform 1 0 39928 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1018_
timestamp 18001
transform 1 0 40480 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1019_
timestamp 18001
transform -1 0 22540 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1020_
timestamp 18001
transform 1 0 21160 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1021_
timestamp 18001
transform 1 0 51336 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1022_
timestamp 18001
transform 1 0 51980 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1023_
timestamp 18001
transform 1 0 19596 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1024_
timestamp 18001
transform 1 0 20056 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1025_
timestamp 18001
transform -1 0 20424 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1026_
timestamp 18001
transform 1 0 18860 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1027_
timestamp 18001
transform -1 0 50048 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1028_
timestamp 18001
transform 1 0 49404 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1029_
timestamp 18001
transform 1 0 50692 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1030_
timestamp 18001
transform 1 0 51612 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1031_
timestamp 18001
transform 1 0 35512 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1032_
timestamp 18001
transform 1 0 36156 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1033_
timestamp 18001
transform -1 0 38732 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1034_
timestamp 18001
transform 1 0 37720 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1035_
timestamp 18001
transform -1 0 20148 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1036_
timestamp 18001
transform 1 0 18860 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1037_
timestamp 18001
transform 1 0 52808 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1038_
timestamp 18001
transform 1 0 53452 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1039_
timestamp 18001
transform -1 0 20056 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1040_
timestamp 18001
transform 1 0 18768 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1041_
timestamp 18001
transform -1 0 19964 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1042_
timestamp 18001
transform 1 0 19964 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1043_
timestamp 18001
transform 1 0 50140 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1044_
timestamp 18001
transform 1 0 50692 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1045_
timestamp 18001
transform 1 0 53268 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1046_
timestamp 18001
transform 1 0 53452 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1047_
timestamp 18001
transform 1 0 34500 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1048_
timestamp 18001
transform 1 0 34868 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1049_
timestamp 18001
transform -1 0 37076 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1050_
timestamp 18001
transform 1 0 35696 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1051_
timestamp 18001
transform -1 0 19964 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1052_
timestamp 18001
transform 1 0 18492 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1053_
timestamp 18001
transform 1 0 55292 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1054_
timestamp 18001
transform -1 0 56580 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1055_
timestamp 18001
transform -1 0 20148 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1056_
timestamp 18001
transform 1 0 18860 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1057_
timestamp 18001
transform -1 0 22632 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1058_
timestamp 18001
transform -1 0 21436 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1059_
timestamp 18001
transform 1 0 51520 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1060_
timestamp 18001
transform 1 0 52440 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1061_
timestamp 18001
transform 1 0 54464 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1062_
timestamp 18001
transform -1 0 55660 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1063_
timestamp 18001
transform -1 0 34040 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1064_
timestamp 18001
transform 1 0 32752 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1065_
timestamp 18001
transform -1 0 36156 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1066_
timestamp 18001
transform 1 0 34868 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1067_
timestamp 18001
transform 1 0 19228 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1068_
timestamp 18001
transform 1 0 19228 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1069_
timestamp 18001
transform -1 0 57592 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1070_
timestamp 18001
transform 1 0 56580 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1071_
timestamp 18001
transform -1 0 20792 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1072_
timestamp 18001
transform 1 0 18492 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1073_
timestamp 18001
transform -1 0 24012 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1074_
timestamp 18001
transform 1 0 22632 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1075_
timestamp 18001
transform -1 0 53452 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1076_
timestamp 18001
transform 1 0 51612 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1077_
timestamp 18001
transform 1 0 55660 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1078_
timestamp 18001
transform -1 0 56856 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1079_
timestamp 18001
transform -1 0 32936 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1080_
timestamp 18001
transform 1 0 32108 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1081_
timestamp 18001
transform -1 0 36340 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1082_
timestamp 18001
transform 1 0 34684 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1083_
timestamp 18001
transform -1 0 20424 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1084_
timestamp 18001
transform -1 0 20332 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1085_
timestamp 18001
transform 1 0 56304 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1086_
timestamp 18001
transform 1 0 56212 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1087_
timestamp 18001
transform -1 0 25760 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1088_
timestamp 18001
transform 1 0 21804 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1089_
timestamp 18001
transform -1 0 25576 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1090_
timestamp 18001
transform 1 0 24380 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1091_
timestamp 18001
transform 1 0 54004 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1092_
timestamp 18001
transform 1 0 56028 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1093_
timestamp 18001
transform 1 0 54556 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1094_
timestamp 18001
transform -1 0 55844 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1095_
timestamp 18001
transform 1 0 32108 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1096_
timestamp 18001
transform 1 0 33028 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1097_
timestamp 18001
transform -1 0 37260 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1098_
timestamp 18001
transform 1 0 35972 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1099_
timestamp 18001
transform -1 0 22908 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1100_
timestamp 18001
transform 1 0 21988 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1101_
timestamp 18001
transform 1 0 53452 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1102_
timestamp 18001
transform 1 0 54280 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1103_
timestamp 18001
transform -1 0 24104 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1104_
timestamp 18001
transform 1 0 23644 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1105_
timestamp 18001
transform -1 0 26404 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1106_
timestamp 18001
transform 1 0 25116 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1107_
timestamp 18001
transform 1 0 55200 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1108_
timestamp 18001
transform 1 0 56120 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1109_
timestamp 18001
transform 1 0 51796 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1110_
timestamp 18001
transform -1 0 52624 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1111_
timestamp 18001
transform -1 0 32752 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1112_
timestamp 18001
transform 1 0 31372 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1113_
timestamp 18001
transform 1 0 40572 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1114_
timestamp 18001
transform -1 0 41860 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1115_
timestamp 18001
transform -1 0 24012 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1116_
timestamp 18001
transform 1 0 22724 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1117_
timestamp 18001
transform 1 0 52716 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1118_
timestamp 18001
transform 1 0 52716 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1119_
timestamp 18001
transform -1 0 26772 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1120_
timestamp 18001
transform -1 0 26864 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1121_
timestamp 18001
transform -1 0 28152 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1122_
timestamp 18001
transform 1 0 27692 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1123_
timestamp 18001
transform 1 0 53176 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1124_
timestamp 18001
transform -1 0 54648 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1125_
timestamp 18001
transform 1 0 49128 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1126_
timestamp 18001
transform 1 0 50876 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1127_
timestamp 18001
transform 1 0 32108 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1128_
timestamp 18001
transform 1 0 32384 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1129_
timestamp 18001
transform 1 0 38364 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1130_
timestamp 18001
transform 1 0 39008 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1131_
timestamp 18001
transform -1 0 26312 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1132_
timestamp 18001
transform -1 0 25944 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1133_
timestamp 18001
transform 1 0 49956 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1134_
timestamp 18001
transform 1 0 50600 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1135_
timestamp 18001
transform 1 0 28244 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1136_
timestamp 18001
transform 1 0 29532 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1137_
timestamp 18001
transform 1 0 28336 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1138_
timestamp 18001
transform 1 0 28520 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1139_
timestamp 18001
transform 1 0 50324 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1140_
timestamp 18001
transform 1 0 50508 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1141_
timestamp 18001
transform -1 0 48576 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1142_
timestamp 18001
transform 1 0 47472 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1143_
timestamp 18001
transform 1 0 32108 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1144_
timestamp 18001
transform 1 0 32108 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1145_
timestamp 18001
transform -1 0 39560 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1146_
timestamp 18001
transform 1 0 37904 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1147_
timestamp 18001
transform 1 0 24288 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1148_
timestamp 18001
transform 1 0 25576 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1149_
timestamp 18001
transform 1 0 46828 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o22a_1  _1150_
timestamp 18001
transform 1 0 47564 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1151_
timestamp 18001
transform 1 0 28888 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o22a_1  _1152_
timestamp 18001
transform -1 0 30176 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1153_
timestamp 18001
transform -1 0 29072 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o22a_1  _1154_
timestamp 18001
transform 1 0 27968 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1155_
timestamp 18001
transform 1 0 52716 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o22a_1  _1156_
timestamp 18001
transform -1 0 54096 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1157_
timestamp 18001
transform 1 0 44988 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__o22a_1  _1158_
timestamp 18001
transform 1 0 44988 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1159_
timestamp 18001
transform 1 0 33120 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _1160_
timestamp 18001
transform 1 0 31372 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1161_
timestamp 18001
transform -1 0 39560 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o22a_1  _1162_
timestamp 18001
transform 1 0 38456 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1163_
timestamp 18001
transform -1 0 26864 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1164_
timestamp 18001
transform 1 0 26128 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__or4b_4  _1165_
timestamp 18001
transform -1 0 32844 0 1 7616
box -38 -48 1050 592
use sky130_fd_sc_hd__nor2_1  _1166_
timestamp 18001
transform 1 0 27140 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1167_
timestamp 18001
transform -1 0 26404 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1168_
timestamp 18001
transform -1 0 36708 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__nand4b_1  _1169_
timestamp 18001
transform 1 0 32936 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _1170_
timestamp 18001
transform 1 0 33488 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__or4_2  _1171_
timestamp 18001
transform -1 0 33672 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1172_
timestamp 18001
transform -1 0 39008 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _1173_
timestamp 18001
transform 1 0 40020 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _1174_
timestamp 18001
transform -1 0 44804 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__nand3b_1  _1175_
timestamp 18001
transform -1 0 44344 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_1  _1176_
timestamp 18001
transform 1 0 40204 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1177_
timestamp 18001
transform 1 0 40204 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_2  _1178_
timestamp 18001
transform -1 0 44896 0 1 29376
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_1  _1179_
timestamp 18001
transform -1 0 44528 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1180_
timestamp 18001
transform -1 0 40940 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1181_
timestamp 18001
transform 1 0 41216 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_2  _1182_
timestamp 18001
transform 1 0 40480 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__or4bb_1  _1183_
timestamp 18001
transform 1 0 33304 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__or4bb_1  _1184_
timestamp 18001
transform 1 0 34132 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__or4_4  _1185_
timestamp 18001
transform -1 0 34500 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _1186_
timestamp 18001
transform 1 0 37904 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1187_
timestamp 18001
transform -1 0 43148 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1188_
timestamp 18001
transform 1 0 44988 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1189_
timestamp 18001
transform 1 0 43608 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1190_
timestamp 18001
transform 1 0 43056 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_2  _1191_
timestamp 18001
transform 1 0 42412 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1192_
timestamp 18001
transform -1 0 41400 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1193_
timestamp 18001
transform 1 0 41860 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1194_
timestamp 18001
transform -1 0 39100 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1195_
timestamp 18001
transform 1 0 37260 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _1196_
timestamp 18001
transform 1 0 40112 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__o211ai_2  _1197_
timestamp 18001
transform 1 0 40940 0 1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__o22a_1  _1198_
timestamp 18001
transform 1 0 40940 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1199_
timestamp 18001
transform -1 0 40388 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1200_
timestamp 18001
transform 1 0 39836 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1201_
timestamp 18001
transform 1 0 43424 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _1202_
timestamp 18001
transform 1 0 43608 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__and4bb_1  _1203_
timestamp 18001
transform 1 0 42872 0 -1 29376
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _1204_
timestamp 18001
transform -1 0 45448 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_2  _1205_
timestamp 18001
transform 1 0 42872 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1206_
timestamp 18001
transform -1 0 42780 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1207_
timestamp 18001
transform 1 0 44344 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_4  _1208_
timestamp 18001
transform 1 0 43148 0 -1 28288
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _1209_
timestamp 18001
transform 1 0 45632 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1210_
timestamp 18001
transform -1 0 46552 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1211_
timestamp 18001
transform 1 0 43148 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1212_
timestamp 18001
transform 1 0 43424 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1213_
timestamp 18001
transform 1 0 46460 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1214_
timestamp 18001
transform 1 0 25944 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1215_
timestamp 18001
transform 1 0 26036 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1216_
timestamp 18001
transform 1 0 28336 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1217_
timestamp 18001
transform 1 0 27508 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1218_
timestamp 18001
transform 1 0 29532 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1219_
timestamp 18001
transform 1 0 32292 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1220_
timestamp 18001
transform 1 0 30912 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1221_
timestamp 18001
transform 1 0 33304 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__or4b_4  _1222_
timestamp 18001
transform 1 0 27968 0 1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__or2_1  _1223_
timestamp 18001
transform 1 0 33764 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _1224_
timestamp 18001
transform 1 0 39100 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_1  _1225_
timestamp 18001
transform -1 0 24840 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1226_
timestamp 18001
transform -1 0 26496 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1227_
timestamp 18001
transform 1 0 25208 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1228_
timestamp 18001
transform 1 0 26496 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__o21bai_1  _1229_
timestamp 18001
transform 1 0 25760 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _1230_
timestamp 18001
transform 1 0 26220 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1231_
timestamp 18001
transform 1 0 26956 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1232_
timestamp 18001
transform -1 0 26680 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__o21bai_1  _1233_
timestamp 18001
transform 1 0 25484 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1234_
timestamp 18001
transform -1 0 23460 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1235_
timestamp 18001
transform 1 0 21804 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1236_
timestamp 18001
transform -1 0 21988 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1237_
timestamp 18001
transform 1 0 20240 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1238_
timestamp 18001
transform 1 0 16928 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1239_
timestamp 18001
transform 1 0 16652 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1240_
timestamp 18001
transform -1 0 16560 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1241_
timestamp 18001
transform -1 0 18216 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1242_
timestamp 18001
transform -1 0 18216 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _1243_
timestamp 18001
transform -1 0 18768 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _1244_
timestamp 18001
transform -1 0 16376 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1245_
timestamp 18001
transform 1 0 17940 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1246_
timestamp 18001
transform -1 0 15640 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1247_
timestamp 18001
transform 1 0 18124 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1248_
timestamp 18001
transform 1 0 18768 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1249_
timestamp 18001
transform 1 0 18492 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1250_
timestamp 18001
transform 1 0 19228 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1251_
timestamp 18001
transform 1 0 19964 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1252_
timestamp 18001
transform -1 0 22540 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1253_
timestamp 18001
transform -1 0 23184 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1254_
timestamp 18001
transform -1 0 22080 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1255_
timestamp 18001
transform -1 0 23184 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1256_
timestamp 18001
transform 1 0 24840 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1257_
timestamp 18001
transform -1 0 25024 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1258_
timestamp 18001
transform -1 0 26404 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1259_
timestamp 18001
transform 1 0 25300 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_4  _1260_
timestamp 18001
transform 1 0 28152 0 -1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__nor2_1  _1261_
timestamp 18001
transform 1 0 32844 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1262_
timestamp 18001
transform 1 0 28888 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1263_
timestamp 18001
transform -1 0 28060 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or4b_4  _1264_
timestamp 18001
transform 1 0 28060 0 1 7616
box -38 -48 1050 592
use sky130_fd_sc_hd__o22a_1  _1265_
timestamp 18001
transform -1 0 32844 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1266_
timestamp 18001
transform -1 0 29256 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1267_
timestamp 18001
transform 1 0 31096 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__o22ai_1  _1268_
timestamp 18001
transform -1 0 33764 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1269_
timestamp 18001
transform 1 0 34684 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _1270_
timestamp 18001
transform -1 0 29440 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1271_
timestamp 18001
transform 1 0 34408 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1272_
timestamp 18001
transform 1 0 37904 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1273_
timestamp 18001
transform -1 0 36524 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_2  _1274_
timestamp 18001
transform 1 0 36064 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1275_
timestamp 18001
transform -1 0 39284 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _1276_
timestamp 18001
transform 1 0 35972 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _1277_
timestamp 18001
transform -1 0 32844 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1278_
timestamp 18001
transform 1 0 32016 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1279_
timestamp 18001
transform -1 0 37720 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1280_
timestamp 18001
transform -1 0 33856 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1281_
timestamp 18001
transform -1 0 30452 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1282_
timestamp 18001
transform 1 0 35788 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1283_
timestamp 18001
transform -1 0 32936 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1284_
timestamp 18001
transform -1 0 38548 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nor4_1  _1285_
timestamp 18001
transform -1 0 37996 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1286_
timestamp 18001
transform -1 0 33488 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_4  _1287_
timestamp 18001
transform -1 0 35972 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1288_
timestamp 18001
transform 1 0 32108 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1289_
timestamp 18001
transform 1 0 39836 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1290_
timestamp 18001
transform -1 0 38272 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1291_
timestamp 18001
transform -1 0 36800 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _1292_
timestamp 18001
transform 1 0 34960 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1293_
timestamp 18001
transform -1 0 36248 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _1294_
timestamp 18001
transform 1 0 35328 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a311o_1  _1295_
timestamp 18001
transform -1 0 35512 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _1296_
timestamp 18001
transform -1 0 35512 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1297_
timestamp 18001
transform 1 0 42412 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1298_
timestamp 18001
transform 1 0 38364 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1299_
timestamp 18001
transform -1 0 33580 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1300_
timestamp 18001
transform -1 0 29716 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1301_
timestamp 18001
transform 1 0 32200 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1302_
timestamp 18001
transform 1 0 31924 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_2  _1303_
timestamp 18001
transform -1 0 32752 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1304_
timestamp 18001
transform 1 0 36708 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a2111oi_1  _1305_
timestamp 18001
transform 1 0 28612 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _1306_
timestamp 18001
transform -1 0 31464 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_1  _1307_
timestamp 18001
transform 1 0 30636 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1308_
timestamp 18001
transform 1 0 30268 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _1309_
timestamp 18001
transform -1 0 31832 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1310_
timestamp 18001
transform -1 0 30820 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1311_
timestamp 18001
transform 1 0 32108 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1312_
timestamp 18001
transform 1 0 30636 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _1313_
timestamp 18001
transform 1 0 29532 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1314_
timestamp 18001
transform 1 0 33488 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1315_
timestamp 18001
transform 1 0 29900 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _1316_
timestamp 18001
transform 1 0 28244 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1317_
timestamp 18001
transform 1 0 29256 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o32ai_1  _1318_
timestamp 18001
transform -1 0 29440 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1319_
timestamp 18001
transform -1 0 30268 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _1320_
timestamp 18001
transform -1 0 30268 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__o31a_1  _1321_
timestamp 18001
transform 1 0 28520 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1322_
timestamp 18001
transform 1 0 27232 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1323_
timestamp 18001
transform -1 0 27968 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o22a_1  _1324_
timestamp 18001
transform 1 0 27968 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a2111o_1  _1325_
timestamp 18001
transform 1 0 32660 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _1326_
timestamp 18001
transform 1 0 32568 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__o2bb2a_1  _1327_
timestamp 18001
transform -1 0 33580 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1328_
timestamp 18001
transform 1 0 33028 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__a21bo_1  _1329_
timestamp 18001
transform 1 0 39836 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1330_
timestamp 18001
transform -1 0 39192 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1331_
timestamp 18001
transform -1 0 39652 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1332_
timestamp 18001
transform 1 0 38640 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1333_
timestamp 18001
transform -1 0 39836 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1334_
timestamp 18001
transform -1 0 40204 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1335_
timestamp 18001
transform 1 0 40572 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a31oi_1  _1336_
timestamp 18001
transform -1 0 38916 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1337_
timestamp 18001
transform -1 0 39560 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__o311a_1  _1338_
timestamp 18001
transform 1 0 37628 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _1339_
timestamp 18001
transform 1 0 36432 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_1  _1340_
timestamp 18001
transform -1 0 36984 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1341_
timestamp 18001
transform -1 0 36340 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a221oi_1  _1342_
timestamp 18001
transform -1 0 39560 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_1  _1343_
timestamp 18001
transform 1 0 39008 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1344_
timestamp 18001
transform -1 0 31188 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1345_
timestamp 18001
transform 1 0 29532 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1346_
timestamp 18001
transform 1 0 41400 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _1347_
timestamp 18001
transform 1 0 39100 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1348_
timestamp 18001
transform -1 0 39744 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _1349_
timestamp 18001
transform 1 0 38824 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1350_
timestamp 18001
transform -1 0 40480 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__and4b_1  _1351_
timestamp 18001
transform -1 0 40572 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1352_
timestamp 18001
transform -1 0 39836 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__a21boi_2  _1353_
timestamp 18001
transform -1 0 41308 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__o211a_1  _1354_
timestamp 18001
transform -1 0 42320 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _1355_
timestamp 18001
transform 1 0 43240 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1356_
timestamp 18001
transform 1 0 40572 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_2  _1357_
timestamp 18001
transform 1 0 39468 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1358_
timestamp 18001
transform 1 0 39008 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1359_
timestamp 18001
transform -1 0 43700 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__a2111o_1  _1360_
timestamp 18001
transform -1 0 42228 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__a21bo_1  _1361_
timestamp 18001
transform -1 0 56764 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1362_
timestamp 18001
transform -1 0 23368 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nand4_1  _1363_
timestamp 18001
transform -1 0 22264 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1364_
timestamp 18001
transform 1 0 20516 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1365_
timestamp 18001
transform -1 0 22356 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1366_
timestamp 18001
transform 1 0 20792 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1367_
timestamp 18001
transform 1 0 23460 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and4b_1  _1368_
timestamp 18001
transform 1 0 22264 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1369_
timestamp 18001
transform -1 0 22908 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__nand4b_1  _1370_
timestamp 18001
transform 1 0 22080 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1371_
timestamp 18001
transform -1 0 23828 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__and2_4  _1372_
timestamp 18001
transform 1 0 43240 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__and3_4  _1373_
timestamp 18001
transform 1 0 39560 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__and3_4  _1374_
timestamp 18001
transform -1 0 40664 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__and3_4  _1375_
timestamp 18001
transform 1 0 38732 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _1376_
timestamp 18001
transform 1 0 42688 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__and3_4  _1377_
timestamp 18001
transform 1 0 43332 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__and3_4  _1378_
timestamp 18001
transform 1 0 42504 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1379_
timestamp 18001
transform -1 0 50416 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__and3_4  _1380_
timestamp 18001
transform 1 0 43056 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__and3_4  _1381_
timestamp 18001
transform 1 0 42228 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__and2_2  _1382_
timestamp 18001
transform 1 0 38272 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__and2_4  _1383_
timestamp 18001
transform 1 0 42504 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__and3_4  _1384_
timestamp 18001
transform 1 0 42412 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__and2_2  _1385_
timestamp 18001
transform 1 0 44344 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__and3_4  _1386_
timestamp 18001
transform 1 0 42412 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__and3_4  _1387_
timestamp 18001
transform 1 0 39560 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__and2_4  _1388_
timestamp 18001
transform 1 0 38088 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _1389_
timestamp 18001
transform 1 0 39836 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1390_
timestamp 18001
transform -1 0 49036 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1391_
timestamp 18001
transform -1 0 49864 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1392_
timestamp 18001
transform -1 0 50416 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1393_
timestamp 18001
transform 1 0 48852 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1394_
timestamp 18001
transform 1 0 48300 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1395_
timestamp 18001
transform 1 0 46000 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1396_
timestamp 18001
transform 1 0 47656 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1397_
timestamp 18001
transform 1 0 49404 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1398_
timestamp 18001
transform -1 0 57500 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1399_
timestamp 18001
transform 1 0 24196 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1400_
timestamp 18001
transform 1 0 24840 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1401_
timestamp 18001
transform 1 0 24472 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1402_
timestamp 18001
transform 1 0 27968 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1403_
timestamp 18001
transform 1 0 25392 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1404_
timestamp 18001
transform 1 0 25852 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1405_
timestamp 18001
transform 1 0 37904 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1406_
timestamp 18001
transform -1 0 31832 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1407_
timestamp 18001
transform 1 0 25208 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1408_
timestamp 18001
transform 1 0 26588 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1409_
timestamp 18001
transform 1 0 21896 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1410_
timestamp 18001
transform 1 0 24472 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1411_
timestamp 18001
transform 1 0 24932 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1412_
timestamp 18001
transform 1 0 25484 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1413_
timestamp 18001
transform -1 0 28796 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1414_
timestamp 18001
transform -1 0 26772 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1415_
timestamp 18001
transform 1 0 25484 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1416_
timestamp 18001
transform -1 0 26312 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1417_
timestamp 18001
transform -1 0 30636 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _1418_
timestamp 18001
transform 1 0 25576 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1419_
timestamp 18001
transform -1 0 25484 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1420_
timestamp 18001
transform 1 0 23276 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1421_
timestamp 18001
transform 1 0 48760 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1422_
timestamp 18001
transform 1 0 49680 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1423_
timestamp 18001
transform 1 0 49036 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1424_
timestamp 18001
transform 1 0 50048 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_1  _1425_
timestamp 18001
transform -1 0 43884 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1426_
timestamp 18001
transform -1 0 42504 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1427_
timestamp 18001
transform -1 0 50876 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1428_
timestamp 18001
transform 1 0 44896 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1429_
timestamp 18001
transform 1 0 47380 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1430_
timestamp 18001
transform 1 0 48208 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1431_
timestamp 18001
transform -1 0 50048 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1432_
timestamp 18001
transform 1 0 49036 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1433_
timestamp 18001
transform 1 0 49956 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1434_
timestamp 18001
transform -1 0 44436 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1435_
timestamp 18001
transform -1 0 57592 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1436_
timestamp 18001
transform 1 0 47380 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1437_
timestamp 18001
transform -1 0 49496 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1438_
timestamp 18001
transform 1 0 46828 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1439_
timestamp 18001
transform -1 0 49128 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1440_
timestamp 18001
transform 1 0 48300 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1441_
timestamp 18001
transform -1 0 50876 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1442_
timestamp 18001
transform 1 0 44068 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1443_
timestamp 18001
transform 1 0 47564 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1444_
timestamp 18001
transform 1 0 49036 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1445_
timestamp 18001
transform -1 0 57592 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1446_
timestamp 18001
transform -1 0 29992 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1447_
timestamp 18001
transform 1 0 34224 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1448_
timestamp 18001
transform -1 0 35696 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _1449_
timestamp 18001
transform -1 0 38456 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1450_
timestamp 18001
transform 1 0 36616 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1451_
timestamp 18001
transform -1 0 38272 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1452_
timestamp 18001
transform -1 0 39192 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1453_
timestamp 18001
transform -1 0 37812 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1454_
timestamp 18001
transform -1 0 33856 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1455_
timestamp 18001
transform 1 0 33120 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1456_
timestamp 18001
transform -1 0 34592 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1457_
timestamp 18001
transform 1 0 34040 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1458_
timestamp 18001
transform -1 0 34592 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1459_
timestamp 18001
transform -1 0 29348 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1460_
timestamp 18001
transform 1 0 42412 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1461_
timestamp 18001
transform 1 0 43056 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1462_
timestamp 18001
transform -1 0 40480 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1463_
timestamp 18001
transform 1 0 39652 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1464_
timestamp 18001
transform 1 0 38548 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1465_
timestamp 18001
transform 1 0 39928 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1466_
timestamp 18001
transform 1 0 37720 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1467_
timestamp 18001
transform 1 0 39284 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1468_
timestamp 18001
transform 1 0 39836 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1469_
timestamp 18001
transform 1 0 40664 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1470_
timestamp 18001
transform -1 0 57500 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1471_
timestamp 18001
transform 1 0 26220 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1472_
timestamp 18001
transform 1 0 24012 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1473_
timestamp 18001
transform 1 0 24380 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1474_
timestamp 18001
transform 1 0 24380 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1475_
timestamp 18001
transform -1 0 29440 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1476_
timestamp 18001
transform 1 0 26312 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1477_
timestamp 18001
transform 1 0 25300 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1478_
timestamp 18001
transform -1 0 31096 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__a2111o_1  _1479_
timestamp 18001
transform 1 0 25392 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__or4_1  _1480_
timestamp 18001
transform -1 0 25392 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1481_
timestamp 18001
transform 1 0 16100 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _1482_
timestamp 18001
transform 1 0 28428 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1483_
timestamp 18001
transform -1 0 28980 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1484_
timestamp 18001
transform -1 0 29808 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1485_
timestamp 18001
transform -1 0 30544 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _1486_
timestamp 18001
transform -1 0 37168 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1487_
timestamp 18001
transform -1 0 40664 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1488_
timestamp 18001
transform 1 0 45172 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1489_
timestamp 18001
transform 1 0 30728 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1490_
timestamp 18001
transform 1 0 27508 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1491_
timestamp 18001
transform 1 0 40388 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1492_
timestamp 18001
transform 1 0 40480 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _1493_
timestamp 18001
transform 1 0 34132 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1494_
timestamp 18001
transform -1 0 42320 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1495_
timestamp 18001
transform 1 0 30176 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1496_
timestamp 18001
transform 1 0 46000 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1497_
timestamp 18001
transform -1 0 32476 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1498_
timestamp 18001
transform -1 0 27416 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1499_
timestamp 18001
transform 1 0 44068 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1500_
timestamp 18001
transform 1 0 40848 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _1501_
timestamp 18001
transform 1 0 33580 0 -1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1502_
timestamp 18001
transform 1 0 42412 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1503_
timestamp 18001
transform -1 0 33120 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1504_
timestamp 18001
transform 1 0 45632 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1505_
timestamp 18001
transform 1 0 27600 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1506_
timestamp 18001
transform 1 0 22080 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1507_
timestamp 18001
transform -1 0 48484 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1508_
timestamp 18001
transform -1 0 44896 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _1509_
timestamp 18001
transform 1 0 34776 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1510_
timestamp 18001
transform -1 0 44988 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1511_
timestamp 18001
transform 1 0 29348 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1512_
timestamp 18001
transform 1 0 48116 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1513_
timestamp 18001
transform -1 0 26864 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1514_
timestamp 18001
transform 1 0 21804 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1515_
timestamp 18001
transform 1 0 45632 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1516_
timestamp 18001
transform 1 0 44988 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _1517_
timestamp 18001
transform -1 0 38088 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1518_
timestamp 18001
transform 1 0 43424 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1519_
timestamp 18001
transform 1 0 26956 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1520_
timestamp 18001
transform 1 0 48760 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1521_
timestamp 18001
transform 1 0 22264 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1522_
timestamp 18001
transform 1 0 19228 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1523_
timestamp 18001
transform 1 0 45540 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1524_
timestamp 18001
transform -1 0 48944 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _1525_
timestamp 18001
transform -1 0 36800 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1526_
timestamp 18001
transform 1 0 42596 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1527_
timestamp 18001
transform 1 0 22356 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1528_
timestamp 18001
transform 1 0 50140 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1529_
timestamp 18001
transform -1 0 22264 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1530_
timestamp 18001
transform 1 0 18216 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1531_
timestamp 18001
transform 1 0 46552 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1532_
timestamp 18001
transform 1 0 49680 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _1533_
timestamp 18001
transform 1 0 34684 0 1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1534_
timestamp 18001
transform 1 0 40020 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1535_
timestamp 18001
transform 1 0 20516 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1536_
timestamp 18001
transform 1 0 51428 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1537_
timestamp 18001
transform 1 0 18216 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1538_
timestamp 18001
transform 1 0 17940 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1539_
timestamp 18001
transform 1 0 48852 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1540_
timestamp 18001
transform 1 0 51428 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _1541_
timestamp 18001
transform -1 0 37076 0 -1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1542_
timestamp 18001
transform 1 0 37260 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1543_
timestamp 18001
transform 1 0 17020 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1544_
timestamp 18001
transform 1 0 52992 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1545_
timestamp 18001
transform 1 0 17296 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1546_
timestamp 18001
transform 1 0 17296 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1547_
timestamp 18001
transform 1 0 50140 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1548_
timestamp 18001
transform 1 0 53360 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _1549_
timestamp 18001
transform 1 0 34684 0 1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1550_
timestamp 18001
transform 1 0 34868 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1551_
timestamp 18001
transform 1 0 16652 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1552_
timestamp 18001
transform -1 0 56764 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1553_
timestamp 18001
transform 1 0 18492 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1554_
timestamp 18001
transform 1 0 21804 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1555_
timestamp 18001
transform 1 0 52716 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1556_
timestamp 18001
transform 1 0 55292 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _1557_
timestamp 18001
transform 1 0 32476 0 1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1558_
timestamp 18001
transform 1 0 33580 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1559_
timestamp 18001
transform 1 0 17848 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1560_
timestamp 18001
transform 1 0 55936 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1561_
timestamp 18001
transform 1 0 19228 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1562_
timestamp 18001
transform 1 0 21436 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1563_
timestamp 18001
transform 1 0 52164 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1564_
timestamp 18001
transform -1 0 58144 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _1565_
timestamp 18001
transform 1 0 30544 0 1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1566_
timestamp 18001
transform 1 0 33488 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1567_
timestamp 18001
transform -1 0 21068 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1568_
timestamp 18001
transform 1 0 55936 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1569_
timestamp 18001
transform 1 0 21804 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1570_
timestamp 18001
transform 1 0 23184 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1571_
timestamp 18001
transform -1 0 56304 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1572_
timestamp 18001
transform -1 0 56212 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _1573_
timestamp 18001
transform 1 0 31096 0 1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1574_
timestamp 18001
transform 1 0 35328 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1575_
timestamp 18001
transform 1 0 21436 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1576_
timestamp 18001
transform 1 0 54096 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1577_
timestamp 18001
transform 1 0 22448 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1578_
timestamp 18001
transform 1 0 25024 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1579_
timestamp 18001
transform 1 0 55936 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1580_
timestamp 18001
transform 1 0 52716 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _1581_
timestamp 18001
transform 1 0 31004 0 1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1582_
timestamp 18001
transform 1 0 41216 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1583_
timestamp 18001
transform 1 0 21804 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1584_
timestamp 18001
transform 1 0 52440 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1585_
timestamp 18001
transform 1 0 26956 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1586_
timestamp 18001
transform 1 0 27324 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1587_
timestamp 18001
transform 1 0 54004 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1588_
timestamp 18001
transform -1 0 52072 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _1589_
timestamp 18001
transform -1 0 32384 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1590_
timestamp 18001
transform 1 0 37904 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1591_
timestamp 18001
transform -1 0 26588 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1592_
timestamp 18001
transform 1 0 50600 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1593_
timestamp 18001
transform 1 0 29624 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1594_
timestamp 18001
transform 1 0 28336 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1595_
timestamp 18001
transform 1 0 50416 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1596_
timestamp 18001
transform 1 0 47564 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _1597_
timestamp 18001
transform 1 0 31188 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1598_
timestamp 18001
transform 1 0 37076 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1599_
timestamp 18001
transform 1 0 25024 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1600_
timestamp 18001
transform 1 0 46460 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1601_
timestamp 18001
transform -1 0 29440 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1602_
timestamp 18001
transform 1 0 27508 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1603_
timestamp 18001
transform -1 0 53728 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1604_
timestamp 18001
transform 1 0 44252 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _1605_
timestamp 18001
transform 1 0 31188 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1606_
timestamp 18001
transform 1 0 37904 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1607_
timestamp 18001
transform -1 0 25576 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _1608_
timestamp 18001
transform -1 0 39192 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1609_
timestamp 18001
transform -1 0 39744 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1610_
timestamp 18001
transform 1 0 34684 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1611_
timestamp 18001
transform 1 0 24932 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfxtp_1  _1612_
timestamp 18001
transform -1 0 36984 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfrtp_4  _1613_
timestamp 18001
transform 1 0 37352 0 -1 29376
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _1614_
timestamp 18001
transform 1 0 35972 0 1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _1615_
timestamp 18001
transform 1 0 37628 0 1 27200
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1616_
timestamp 18001
transform 1 0 42780 0 -1 30464
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1617_
timestamp 18001
transform -1 0 47472 0 1 29376
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _1618_
timestamp 18001
transform 1 0 46368 0 1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1619_
timestamp 18001
transform 1 0 55476 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1620_
timestamp 18001
transform 1 0 25208 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1621_
timestamp 18001
transform 1 0 25024 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1622_
timestamp 18001
transform 1 0 27692 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1623_
timestamp 18001
transform 1 0 25668 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1624_
timestamp 18001
transform 1 0 29532 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1625_
timestamp 18001
transform 1 0 32108 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1626_
timestamp 18001
transform 1 0 30084 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1627_
timestamp 18001
transform 1 0 32752 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1628_
timestamp 18001
transform 1 0 40204 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1629_
timestamp 18001
transform 1 0 23092 0 -1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1630_
timestamp 18001
transform 1 0 25024 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1631_
timestamp 18001
transform -1 0 28888 0 1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1632_
timestamp 18001
transform -1 0 27876 0 1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1633_
timestamp 18001
transform 1 0 25024 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1634_
timestamp 18001
transform 1 0 20792 0 1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1635_
timestamp 18001
transform 1 0 19872 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1636_
timestamp 18001
transform 1 0 17296 0 -1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1637_
timestamp 18001
transform 1 0 14352 0 1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1638_
timestamp 18001
transform 1 0 17204 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1639_
timestamp 18001
transform 1 0 13892 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1640_
timestamp 18001
transform -1 0 17388 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1641_
timestamp 18001
transform 1 0 18032 0 -1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1642_
timestamp 18001
transform 1 0 20240 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1643_
timestamp 18001
transform 1 0 22080 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1644_
timestamp 18001
transform 1 0 22540 0 -1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1645_
timestamp 18001
transform -1 0 26864 0 -1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1646_
timestamp 18001
transform -1 0 27784 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1647_
timestamp 18001
transform 1 0 42504 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1648_
timestamp 18001
transform 1 0 28612 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1649_
timestamp 18001
transform 1 0 24564 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1650_
timestamp 18001
transform 1 0 32568 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1651_
timestamp 18001
transform 1 0 41676 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _1652_
timestamp 18001
transform -1 0 36616 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1653_
timestamp 18001
transform 1 0 38640 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1654_
timestamp 18001
transform -1 0 29440 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1655_
timestamp 18001
transform 1 0 23644 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1656_
timestamp 18001
transform 1 0 24380 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1657_
timestamp 18001
transform 1 0 26956 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1658_
timestamp 18001
transform 1 0 26220 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1659_
timestamp 18001
transform 1 0 28060 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1660_
timestamp 18001
transform 1 0 29992 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1661_
timestamp 18001
transform 1 0 30636 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1662_
timestamp 18001
transform 1 0 32108 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1663_
timestamp 18001
transform 1 0 31464 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1664_
timestamp 18001
transform 1 0 15548 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1665_
timestamp 18001
transform -1 0 16560 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1666_
timestamp 18001
transform 1 0 12788 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1667_
timestamp 18001
transform 1 0 12052 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1668_
timestamp 18001
transform 1 0 12144 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1669_
timestamp 18001
transform 1 0 14076 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1670_
timestamp 18001
transform -1 0 18492 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1671_
timestamp 18001
transform -1 0 19504 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1672_
timestamp 18001
transform 1 0 19228 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1673_
timestamp 18001
transform -1 0 23644 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1674_
timestamp 18001
transform -1 0 24288 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1675_
timestamp 18001
transform 1 0 19136 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1676_
timestamp 18001
transform -1 0 24840 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1677_
timestamp 18001
transform -1 0 24012 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1678_
timestamp 18001
transform -1 0 24288 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1679_
timestamp 18001
transform -1 0 23828 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1680_
timestamp 18001
transform 1 0 16560 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1681_
timestamp 18001
transform 1 0 18308 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1682_
timestamp 18001
transform 1 0 13064 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1683_
timestamp 18001
transform 1 0 12144 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1684_
timestamp 18001
transform 1 0 12144 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1685_
timestamp 18001
transform 1 0 12144 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1686_
timestamp 18001
transform -1 0 22816 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1687_
timestamp 18001
transform 1 0 19412 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1688_
timestamp 18001
transform 1 0 15364 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1689_
timestamp 18001
transform 1 0 17296 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1690_
timestamp 18001
transform 1 0 12972 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1691_
timestamp 18001
transform 1 0 11960 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1692_
timestamp 18001
transform 1 0 12880 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1693_
timestamp 18001
transform -1 0 17296 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1694_
timestamp 18001
transform 1 0 25576 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1695_
timestamp 18001
transform 1 0 28244 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1696_
timestamp 18001
transform 1 0 28704 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1697_
timestamp 18001
transform 1 0 32108 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1698_
timestamp 18001
transform -1 0 35788 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1699_
timestamp 18001
transform 1 0 31004 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1700_
timestamp 18001
transform 1 0 36892 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1701_
timestamp 18001
transform -1 0 39100 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1702_
timestamp 18001
transform 1 0 37260 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1703_
timestamp 18001
transform 1 0 35788 0 1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1704_
timestamp 18001
transform 1 0 28428 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1705_
timestamp 18001
transform 1 0 29532 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1706_
timestamp 18001
transform 1 0 32936 0 -1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1707_
timestamp 18001
transform 1 0 30176 0 -1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1708_
timestamp 18001
transform 1 0 29072 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1709_
timestamp 18001
transform 1 0 55660 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1710_
timestamp 18001
transform 1 0 19688 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1711_
timestamp 18001
transform 1 0 19688 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1712_
timestamp 18001
transform 1 0 23920 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1713_
timestamp 18001
transform 1 0 23460 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_1  _1714_
timestamp 18001
transform 1 0 56856 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1715_
timestamp 18001
transform 1 0 21804 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1716_
timestamp 18001
transform 1 0 22816 0 1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1717_
timestamp 18001
transform 1 0 56856 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1718_
timestamp 18001
transform 1 0 56856 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1719_
timestamp 18001
transform 1 0 28520 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1720_
timestamp 18001
transform 1 0 56856 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1721_
timestamp 18001
transform -1 0 16468 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _1722__161
timestamp 18001
transform 1 0 45080 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1722_
timestamp 18001
transform -1 0 44804 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1723__162
timestamp 18001
transform 1 0 41400 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1723_
timestamp 18001
transform -1 0 41400 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1724_
timestamp 18001
transform 1 0 37260 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1724__163
timestamp 18001
transform 1 0 37260 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1725__164
timestamp 18001
transform 1 0 42044 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1725_
timestamp 18001
transform -1 0 42044 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1726_
timestamp 18001
transform 1 0 42412 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1726__165
timestamp 18001
transform 1 0 42412 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1727__166
timestamp 18001
transform 1 0 44804 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1727_
timestamp 18001
transform -1 0 44436 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1728_
timestamp 18001
transform -1 0 38180 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1728__167
timestamp 18001
transform 1 0 38180 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1729_
timestamp 18001
transform -1 0 36248 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1729__168
timestamp 18001
transform 1 0 36248 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1730__169
timestamp 18001
transform 1 0 35604 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1730_
timestamp 18001
transform -1 0 35144 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1731_
timestamp 18001
transform 1 0 34408 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1731__170
timestamp 18001
transform -1 0 34408 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1732_
timestamp 18001
transform 1 0 43608 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1732__171
timestamp 18001
transform 1 0 43608 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1733__172
timestamp 18001
transform 1 0 43332 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1733_
timestamp 18001
transform -1 0 43332 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1734__173
timestamp 18001
transform 1 0 38824 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1734_
timestamp 18001
transform -1 0 38824 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1735__174
timestamp 18001
transform 1 0 40756 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1735_
timestamp 18001
transform -1 0 40756 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1736__126
timestamp 18001
transform -1 0 48116 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1736_
timestamp 18001
transform -1 0 47380 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1737__127
timestamp 18001
transform 1 0 24472 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1737_
timestamp 18001
transform 1 0 24748 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1738__128
timestamp 18001
transform -1 0 35236 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1738_
timestamp 18001
transform -1 0 34960 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1739__129
timestamp 18001
transform -1 0 47840 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1739_
timestamp 18001
transform -1 0 47012 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1740_
timestamp 18001
transform 1 0 32108 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1740__130
timestamp 18001
transform 1 0 32016 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1741__131
timestamp 18001
transform -1 0 41032 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1741_
timestamp 18001
transform -1 0 40756 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1742__132
timestamp 18001
transform -1 0 37076 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1742_
timestamp 18001
transform -1 0 36800 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1743__133
timestamp 18001
transform -1 0 29348 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1743_
timestamp 18001
transform -1 0 29072 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1744__134
timestamp 18001
transform -1 0 28152 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1744_
timestamp 18001
transform -1 0 27876 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1745_
timestamp 18001
transform -1 0 25484 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1745__135
timestamp 18001
transform 1 0 25116 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1746__136
timestamp 18001
transform -1 0 41676 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1746_
timestamp 18001
transform -1 0 41400 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1747__137
timestamp 18001
transform -1 0 39100 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1747_
timestamp 18001
transform -1 0 38824 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1748_
timestamp 18001
transform 1 0 35236 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1748__138
timestamp 18001
transform -1 0 35512 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1749__139
timestamp 18001
transform -1 0 38456 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1749_
timestamp 18001
transform -1 0 38180 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1750__140
timestamp 18001
transform -1 0 42320 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1750_
timestamp 18001
transform -1 0 42044 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1751__141
timestamp 18001
transform 1 0 26588 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1751_
timestamp 18001
transform 1 0 26956 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1752_
timestamp 18001
transform -1 0 36892 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1752__175
timestamp 18001
transform 1 0 36892 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1753_
timestamp 18001
transform -1 0 39468 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1753__176
timestamp 18001
transform 1 0 39468 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1754__177
timestamp 18001
transform 1 0 40112 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1754_
timestamp 18001
transform -1 0 40112 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1755_
timestamp 18001
transform 1 0 35236 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1755__178
timestamp 18001
transform 1 0 35328 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1756_
timestamp 18001
transform 1 0 42412 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1756__142
timestamp 18001
transform 1 0 42320 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1757__143
timestamp 18001
transform -1 0 44252 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1757_
timestamp 18001
transform -1 0 43976 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1758__144
timestamp 18001
transform -1 0 44896 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1758_
timestamp 18001
transform -1 0 44620 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1759__145
timestamp 18001
transform -1 0 36432 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1759_
timestamp 18001
transform -1 0 36156 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1760__146
timestamp 18001
transform -1 0 40388 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1760_
timestamp 18001
transform -1 0 40112 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1761__147
timestamp 18001
transform -1 0 33304 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1761_
timestamp 18001
transform -1 0 33028 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1762__148
timestamp 18001
transform -1 0 34592 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1762_
timestamp 18001
transform -1 0 34316 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1763__149
timestamp 18001
transform -1 0 32016 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1763_
timestamp 18001
transform -1 0 31740 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1764_
timestamp 18001
transform 1 0 46184 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1764__150
timestamp 18001
transform -1 0 46460 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1765_
timestamp 18001
transform 1 0 37260 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1765__151
timestamp 18001
transform 1 0 37168 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1766__152
timestamp 18001
transform -1 0 43608 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1766_
timestamp 18001
transform -1 0 43332 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1767__153
timestamp 18001
transform -1 0 33948 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1767_
timestamp 18001
transform -1 0 33672 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1768__154
timestamp 18001
transform -1 0 31372 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1768_
timestamp 18001
transform -1 0 31096 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1769__155
timestamp 18001
transform -1 0 30636 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1769_
timestamp 18001
transform -1 0 30360 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1770_
timestamp 18001
transform -1 0 57684 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1771__156
timestamp 18001
transform -1 0 39744 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1771_
timestamp 18001
transform -1 0 39468 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1772_
timestamp 18001
transform 1 0 31648 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1773_
timestamp 18001
transform -1 0 57684 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1774__157
timestamp 18001
transform -1 0 29992 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1774_
timestamp 18001
transform -1 0 29716 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1775__158
timestamp 18001
transform -1 0 45540 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1775_
timestamp 18001
transform -1 0 45264 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1776__159
timestamp 18001
transform -1 0 26220 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1776_
timestamp 18001
transform -1 0 25944 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _1777__160
timestamp 18001
transform -1 0 46184 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1777_
timestamp 18001
transform -1 0 45908 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0734__Y
timestamp 18001
transform -1 0 33488 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0871__X
timestamp 18001
transform 1 0 35052 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0872__B
timestamp 18001
transform 1 0 25024 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0902__X
timestamp 18001
transform -1 0 20332 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0909__A2
timestamp 18001
transform 1 0 35420 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0911__B2
timestamp 18001
transform 1 0 37812 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0915__A
timestamp 18001
transform 1 0 54464 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0915__Y
timestamp 18001
transform 1 0 54924 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0916__A
timestamp 18001
transform 1 0 36432 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0921__A
timestamp 18001
transform 1 0 36984 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0922__A
timestamp 18001
transform 1 0 33028 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0928__B1
timestamp 18001
transform 1 0 28704 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0929__A1
timestamp 18001
transform 1 0 43056 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0930__A1
timestamp 18001
transform 1 0 41768 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0930__A2
timestamp 18001
transform 1 0 40940 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0932__A2
timestamp 18001
transform 1 0 41124 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0933__B1
timestamp 18001
transform 1 0 36340 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0939__C1
timestamp 18001
transform 1 0 31188 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0941__C1
timestamp 18001
transform 1 0 47656 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0943__C1
timestamp 18001
transform 1 0 31740 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0947__A1
timestamp 18001
transform -1 0 45724 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0947__C1
timestamp 18001
transform -1 0 45540 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0948__A2
timestamp 18001
transform 1 0 44160 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0950__A2
timestamp 18001
transform 1 0 41492 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0955__C1
timestamp 18001
transform 1 0 32476 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0957__C1
timestamp 18001
transform 1 0 47196 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0960__B1
timestamp 18001
transform -1 0 29348 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0964__B1
timestamp 18001
transform 1 0 47288 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0965__B1
timestamp 18001
transform 1 0 45356 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0965__C1
timestamp 18001
transform 1 0 44436 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0971__C1
timestamp 18001
transform 1 0 30268 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0975__C1
timestamp 18001
transform 1 0 25760 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0980__A2
timestamp 18001
transform 1 0 45724 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0981__C1
timestamp 18001
transform 1 0 47104 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0992__B1
timestamp 18001
transform 1 0 23460 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0993__C1
timestamp 18001
transform 1 0 20332 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0996__A2
timestamp 18001
transform 1 0 45816 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1008__B1
timestamp 18001
transform 1 0 22448 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1012__B1
timestamp 18001
transform 1 0 47564 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1022__B1
timestamp 18001
transform 1 0 52624 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1029__C1
timestamp 18001
transform 1 0 50508 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1040__B1
timestamp 18001
transform 1 0 20056 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1045__C1
timestamp 18001
transform 1 0 53084 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1055__C1
timestamp 18001
transform 1 0 20792 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1057__C1
timestamp 18001
transform -1 0 22816 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1059__C1
timestamp 18001
transform 1 0 51336 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1073__C1
timestamp 18001
transform -1 0 24196 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1078__B1
timestamp 18001
transform 1 0 56028 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1086__B1
timestamp 18001
transform 1 0 56028 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1089__C1
timestamp 18001
transform 1 0 24656 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1094__B1
timestamp 18001
transform 1 0 55016 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1102__B1
timestamp 18001
transform 1 0 54924 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1103__C1
timestamp 18001
transform 1 0 24840 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1106__B1
timestamp 18001
transform 1 0 25760 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1118__B1
timestamp 18001
transform 1 0 53360 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1119__C1
timestamp 18001
transform 1 0 25852 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1124__B1
timestamp 18001
transform 1 0 53820 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1131__C1
timestamp 18001
transform 1 0 26312 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1135__B1
timestamp 18001
transform 1 0 29348 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1140__B1
timestamp 18001
transform 1 0 51152 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1142__B1
timestamp 18001
transform 1 0 48116 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1147__C1
timestamp 18001
transform 1 0 24104 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1156__B1
timestamp 18001
transform -1 0 54280 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1158__A2
timestamp 18001
transform 1 0 45632 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1162__A2
timestamp 18001
transform 1 0 39560 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1163__B
timestamp 18001
transform 1 0 27232 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1164__A2
timestamp 18001
transform -1 0 26864 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1172__B
timestamp 18001
transform 1 0 38364 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1185__X
timestamp 18001
transform 1 0 34500 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1195__S
timestamp 18001
transform 1 0 36984 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1200__S
timestamp 18001
transform 1 0 39652 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1201__B
timestamp 18001
transform 1 0 43240 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1206__A1
timestamp 18001
transform 1 0 42136 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1210__S
timestamp 18001
transform 1 0 45540 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1213__S
timestamp 18001
transform 1 0 46276 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1214__S
timestamp 18001
transform -1 0 25944 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1215__S
timestamp 18001
transform 1 0 27508 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1216__S
timestamp 18001
transform 1 0 29164 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1217__S
timestamp 18001
transform 1 0 29532 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1218__S
timestamp 18001
transform 1 0 30360 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1219__S
timestamp 18001
transform 1 0 33120 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1220__S
timestamp 18001
transform 1 0 31740 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1325__A1
timestamp 18001
transform 1 0 34132 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1328__A0
timestamp 18001
transform -1 0 34592 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1352__X
timestamp 18001
transform 1 0 39836 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1358__X
timestamp 18001
transform 1 0 40112 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1359__B1
timestamp 18001
transform 1 0 43700 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1360__B1
timestamp 18001
transform -1 0 41216 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1360__D1
timestamp 18001
transform 1 0 41216 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1361__A2
timestamp 18001
transform 1 0 55844 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1372__X
timestamp 18001
transform 1 0 44068 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1373__X
timestamp 18001
transform 1 0 40572 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1374__X
timestamp 18001
transform -1 0 40848 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1375__X
timestamp 18001
transform 1 0 40388 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1377__X
timestamp 18001
transform -1 0 44528 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1378__X
timestamp 18001
transform -1 0 44344 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1379__A2
timestamp 18001
transform 1 0 50416 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1379__B1
timestamp 18001
transform -1 0 49772 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1380__X
timestamp 18001
transform 1 0 44068 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1381__X
timestamp 18001
transform 1 0 43884 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1382__X
timestamp 18001
transform 1 0 38824 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1383__X
timestamp 18001
transform 1 0 43884 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1384__X
timestamp 18001
transform 1 0 43884 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1385__X
timestamp 18001
transform 1 0 45724 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1386__X
timestamp 18001
transform 1 0 43792 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1387__X
timestamp 18001
transform 1 0 40388 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1388__X
timestamp 18001
transform 1 0 38732 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1389__X
timestamp 18001
transform 1 0 40480 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1390__A2
timestamp 18001
transform -1 0 49220 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1390__B1
timestamp 18001
transform 1 0 49036 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1391__A2
timestamp 18001
transform -1 0 49588 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1391__B1
timestamp 18001
transform -1 0 49404 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1392__A2
timestamp 18001
transform -1 0 50600 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1392__B1
timestamp 18001
transform -1 0 50048 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1393__A2
timestamp 18001
transform 1 0 49036 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1393__B1
timestamp 18001
transform 1 0 48576 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1394__A2
timestamp 18001
transform -1 0 48300 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1394__B1
timestamp 18001
transform -1 0 48116 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1395__A2
timestamp 18001
transform -1 0 46000 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1395__B1
timestamp 18001
transform -1 0 45816 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1396__A2
timestamp 18001
transform 1 0 48208 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1396__B1
timestamp 18001
transform -1 0 47472 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1398__A2
timestamp 18001
transform 1 0 56580 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1399__A2
timestamp 18001
transform 1 0 24840 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1399__B1
timestamp 18001
transform 1 0 25024 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1400__A2
timestamp 18001
transform 1 0 25484 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1400__B1
timestamp 18001
transform 1 0 25668 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1401__A2
timestamp 18001
transform 1 0 24656 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1401__B1
timestamp 18001
transform 1 0 24840 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1402__A2
timestamp 18001
transform 1 0 28704 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1402__B1
timestamp 18001
transform 1 0 28888 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1403__A2
timestamp 18001
transform 1 0 26128 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1403__B1
timestamp 18001
transform 1 0 26312 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1404__A2
timestamp 18001
transform 1 0 26588 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1404__B1
timestamp 18001
transform 1 0 27324 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1405__B1
timestamp 18001
transform 1 0 37720 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1406__A2
timestamp 18001
transform 1 0 31832 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1406__B1
timestamp 18001
transform 1 0 32016 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1407__A2
timestamp 18001
transform 1 0 26956 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1407__B1
timestamp 18001
transform 1 0 26680 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1408__X
timestamp 18001
transform -1 0 27324 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1409__A2
timestamp 18001
transform 1 0 23460 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1409__B1
timestamp 18001
transform -1 0 21896 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1409__C1
timestamp 18001
transform 1 0 22632 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1410__A2
timestamp 18001
transform 1 0 25116 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1410__B1
timestamp 18001
transform 1 0 25300 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1411__A2
timestamp 18001
transform -1 0 24932 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1411__B1
timestamp 18001
transform 1 0 26404 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1412__A2
timestamp 18001
transform -1 0 26772 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1412__B1
timestamp 18001
transform 1 0 26404 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1413__A2
timestamp 18001
transform 1 0 28796 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1413__B1
timestamp 18001
transform 1 0 28980 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1414__A2
timestamp 18001
transform 1 0 27140 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1414__B1
timestamp 18001
transform 1 0 26956 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1415__A2
timestamp 18001
transform 1 0 26220 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1416__A2
timestamp 18001
transform -1 0 26680 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1416__B1
timestamp 18001
transform -1 0 26864 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1416__C1
timestamp 18001
transform 1 0 26312 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1417__A2
timestamp 18001
transform -1 0 30820 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1417__B1
timestamp 18001
transform -1 0 31004 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1418__A2
timestamp 18001
transform 1 0 26220 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1420__A2
timestamp 18001
transform 1 0 24012 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1421__A1
timestamp 18001
transform -1 0 48668 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1421__A2
timestamp 18001
transform 1 0 49404 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1421__B1
timestamp 18001
transform 1 0 48852 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1422__A2
timestamp 18001
transform 1 0 49496 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1422__B1
timestamp 18001
transform 1 0 49312 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1423__A2
timestamp 18001
transform -1 0 49864 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1423__B1
timestamp 18001
transform 1 0 48668 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1424__A2
timestamp 18001
transform -1 0 50784 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1425__B1_N
timestamp 18001
transform 1 0 42504 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1427__A2
timestamp 18001
transform -1 0 51060 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1427__B1
timestamp 18001
transform -1 0 50048 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1428__A
timestamp 18001
transform -1 0 44896 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1429__A2
timestamp 18001
transform 1 0 47196 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1429__B1
timestamp 18001
transform -1 0 47196 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1430__A2
timestamp 18001
transform -1 0 48484 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1430__B1
timestamp 18001
transform -1 0 48300 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1431__A2
timestamp 18001
transform 1 0 49220 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1431__B1
timestamp 18001
transform 1 0 49036 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1434__B1
timestamp 18001
transform 1 0 44436 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1435__A2
timestamp 18001
transform 1 0 56672 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1435__B1
timestamp 18001
transform 1 0 56488 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1436__A2
timestamp 18001
transform 1 0 47748 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1436__B1
timestamp 18001
transform 1 0 47564 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1437__A2
timestamp 18001
transform 1 0 49680 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1437__B1
timestamp 18001
transform 1 0 49496 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1438__A2
timestamp 18001
transform 1 0 46644 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1438__B1
timestamp 18001
transform 1 0 46460 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1439__A2
timestamp 18001
transform -1 0 50048 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1439__B1
timestamp 18001
transform 1 0 47288 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1440__A2
timestamp 18001
transform -1 0 49956 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1440__B1
timestamp 18001
transform 1 0 49588 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1441__A2
timestamp 18001
transform 1 0 50140 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1441__B1
timestamp 18001
transform 1 0 49956 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1442__A2
timestamp 18001
transform 1 0 43884 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1442__B1
timestamp 18001
transform 1 0 45816 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1443__A2
timestamp 18001
transform 1 0 47012 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1443__B1
timestamp 18001
transform 1 0 47196 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1445__A2
timestamp 18001
transform 1 0 56672 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1446__B
timestamp 18001
transform -1 0 28888 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1447__A2
timestamp 18001
transform 1 0 34040 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1447__B1
timestamp 18001
transform 1 0 36616 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1448__A2
timestamp 18001
transform 1 0 36800 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1448__B1
timestamp 18001
transform 1 0 36984 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1449__B1
timestamp 18001
transform -1 0 39376 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1450__A2
timestamp 18001
transform -1 0 37444 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1450__B1
timestamp 18001
transform -1 0 37628 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1452__B1
timestamp 18001
transform -1 0 39560 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1455__A2
timestamp 18001
transform 1 0 33856 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1455__B1
timestamp 18001
transform 1 0 34684 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1456__A2
timestamp 18001
transform 1 0 33764 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1456__B1
timestamp 18001
transform 1 0 34776 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1457__A2
timestamp 18001
transform 1 0 34776 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1457__B1
timestamp 18001
transform 1 0 34960 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1460__A2
timestamp 18001
transform 1 0 43240 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1460__B1
timestamp 18001
transform 1 0 43056 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1461__A2
timestamp 18001
transform 1 0 43792 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1461__B1
timestamp 18001
transform 1 0 42872 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1462__A2
timestamp 18001
transform 1 0 41216 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1462__B1
timestamp 18001
transform 1 0 41400 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1463__A2
timestamp 18001
transform 1 0 39468 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1463__B1
timestamp 18001
transform 1 0 40388 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1464__A2
timestamp 18001
transform 1 0 39744 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1464__B1
timestamp 18001
transform 1 0 41124 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1465__A2
timestamp 18001
transform 1 0 40848 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1465__B1
timestamp 18001
transform 1 0 41032 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1466__A2
timestamp 18001
transform 1 0 38364 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1466__B1
timestamp 18001
transform 1 0 38548 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1467__A2
timestamp 18001
transform -1 0 40756 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1467__B1
timestamp 18001
transform -1 0 40940 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1468__A
timestamp 18001
transform 1 0 40388 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1470__A2
timestamp 18001
transform -1 0 56764 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1471__A2
timestamp 18001
transform -1 0 27048 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1471__B1
timestamp 18001
transform -1 0 27232 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1472__A2
timestamp 18001
transform 1 0 24656 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1472__B1
timestamp 18001
transform 1 0 24656 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1473__A2
timestamp 18001
transform 1 0 25484 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1473__B1
timestamp 18001
transform -1 0 25484 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1474__A2
timestamp 18001
transform -1 0 25300 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1474__B1
timestamp 18001
transform 1 0 25116 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1475__A2
timestamp 18001
transform 1 0 29164 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1475__B1
timestamp 18001
transform -1 0 29348 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1476__A2
timestamp 18001
transform 1 0 26956 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1477__A2
timestamp 18001
transform 1 0 25944 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1477__B1
timestamp 18001
transform 1 0 26128 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1478__A2
timestamp 18001
transform 1 0 31832 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1478__B1
timestamp 18001
transform 1 0 32108 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1478__C1
timestamp 18001
transform -1 0 32476 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1479__A2
timestamp 18001
transform 1 0 26404 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1479__D1
timestamp 18001
transform 1 0 26220 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1481__A2
timestamp 18001
transform 1 0 16836 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1491__Q
timestamp 18001
transform 1 0 42320 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1538__RESET_B
timestamp 18001
transform 1 0 20424 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1548__RESET_B
timestamp 18001
transform 1 0 53176 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1554__RESET_B
timestamp 18001
transform 1 0 21528 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1555__RESET_B
timestamp 18001
transform 1 0 52440 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1579__RESET_B
timestamp 18001
transform 1 0 55752 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1587__RESET_B
timestamp 18001
transform 1 0 53820 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1610__RESET_B
timestamp 18001
transform 1 0 34408 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1613__RESET_B
timestamp 18001
transform 1 0 36984 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1614__RESET_B
timestamp 18001
transform 1 0 37904 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1616__RESET_B
timestamp 18001
transform 1 0 42596 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1617__RESET_B
timestamp 18001
transform -1 0 47656 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1618__RESET_B
timestamp 18001
transform 1 0 48300 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1619__D
timestamp 18001
transform 1 0 55292 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1625__RESET_B
timestamp 18001
transform 1 0 31832 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1641__RESET_B
timestamp 18001
transform 1 0 19872 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1644__RESET_B
timestamp 18001
transform 1 0 22356 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1650__Q
timestamp 18001
transform 1 0 34500 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1700__RESET_B
timestamp 18001
transform 1 0 36248 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1701__RESET_B
timestamp 18001
transform 1 0 36524 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1702__RESET_B
timestamp 18001
transform -1 0 37260 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1703__RESET_B
timestamp 18001
transform 1 0 38088 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_clk_A
timestamp 18001
transform -1 0 36984 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_clk_X
timestamp 18001
transform 1 0 36984 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_1_0__f_clk_A
timestamp 18001
transform 1 0 26404 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_1_0__f_clk_X
timestamp 18001
transform 1 0 26956 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_1_1__f_clk_A
timestamp 18001
transform -1 0 45724 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_1_1__f_clk_X
timestamp 18001
transform 1 0 48668 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_0_clk_A
timestamp 18001
transform 1 0 17664 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_1_clk_A
timestamp 18001
transform 1 0 24748 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_2_clk_A
timestamp 18001
transform 1 0 29808 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_3_clk_A
timestamp 18001
transform 1 0 23000 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_4_clk_A
timestamp 18001
transform 1 0 19320 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_5_clk_A
timestamp 18001
transform 1 0 17848 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_6_clk_A
timestamp 18001
transform -1 0 26220 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_7_clk_A
timestamp 18001
transform 1 0 30452 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_8_clk_A
timestamp 18001
transform 1 0 29256 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_9_clk_A
timestamp 18001
transform 1 0 35972 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_10_clk_A
timestamp 18001
transform 1 0 39100 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_11_clk_A
timestamp 18001
transform 1 0 50048 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_12_clk_A
timestamp 18001
transform 1 0 54004 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_13_clk_A
timestamp 18001
transform 1 0 47564 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_14_clk_A
timestamp 18001
transform 1 0 41768 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_15_clk_A
timestamp 18001
transform 1 0 48392 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_16_clk_A
timestamp 18001
transform -1 0 55476 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_17_clk_A
timestamp 18001
transform 1 0 48484 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_18_clk_A
timestamp 18001
transform 1 0 40848 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_19_clk_A
timestamp 18001
transform 1 0 41032 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_20_clk_A
timestamp 18001
transform 1 0 32200 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_21_clk_A
timestamp 18001
transform 1 0 27600 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_22_clk_A
timestamp 18001
transform 1 0 27692 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_23_clk_A
timestamp 18001
transform 1 0 23276 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_24_clk_A
timestamp 18001
transform 1 0 16560 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_25_clk_A
timestamp 18001
transform 1 0 16376 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkload0_A
timestamp 18001
transform 1 0 47288 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout24_A
timestamp 18001
transform -1 0 29716 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout25_X
timestamp 18001
transform -1 0 29164 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout28_A
timestamp 18001
transform 1 0 38364 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout29_A
timestamp 18001
transform 1 0 48668 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout30_A
timestamp 18001
transform -1 0 52164 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout30_X
timestamp 18001
transform 1 0 53452 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout31_X
timestamp 18001
transform 1 0 39560 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout35_A
timestamp 18001
transform -1 0 28336 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout36_A
timestamp 18001
transform 1 0 24472 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout36_X
timestamp 18001
transform 1 0 24656 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout37_A
timestamp 18001
transform -1 0 34408 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout37_X
timestamp 18001
transform -1 0 34776 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout38_A
timestamp 18001
transform 1 0 47196 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout39_A
timestamp 18001
transform -1 0 47472 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout39_X
timestamp 18001
transform 1 0 47472 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout40_X
timestamp 18001
transform 1 0 33488 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout49_A
timestamp 18001
transform -1 0 38548 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout50_A
timestamp 18001
transform 1 0 42596 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout51_A
timestamp 18001
transform 1 0 39560 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout51_X
timestamp 18001
transform -1 0 39560 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout52_A
timestamp 18001
transform -1 0 53452 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout53_A
timestamp 18001
transform 1 0 52716 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout54_A
timestamp 18001
transform -1 0 47564 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout55_A
timestamp 18001
transform -1 0 55844 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout56_X
timestamp 18001
transform 1 0 40664 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout61_A
timestamp 18001
transform 1 0 27324 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout63_A
timestamp 18001
transform -1 0 25944 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout65_A
timestamp 18001
transform 1 0 37260 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout66_A
timestamp 18001
transform 1 0 36800 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout67_A
timestamp 18001
transform -1 0 37628 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout67_X
timestamp 18001
transform -1 0 37812 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout69_A
timestamp 18001
transform -1 0 48484 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout70_A
timestamp 18001
transform 1 0 55660 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout71_A
timestamp 18001
transform 1 0 54556 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout72_A
timestamp 18001
transform -1 0 53176 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout73_A
timestamp 18001
transform -1 0 56488 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout74_A
timestamp 18001
transform 1 0 54740 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout74_X
timestamp 18001
transform 1 0 55476 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout75_A
timestamp 18001
transform -1 0 30360 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout75_X
timestamp 18001
transform -1 0 30176 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout87_A
timestamp 18001
transform 1 0 39376 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout88_A
timestamp 18001
transform 1 0 49956 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout89_A
timestamp 18001
transform 1 0 51612 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout90_A
timestamp 18001
transform -1 0 49680 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout91_A
timestamp 18001
transform -1 0 52992 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout92_X
timestamp 18001
transform 1 0 39560 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout93_X
timestamp 18001
transform -1 0 38548 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout100_A
timestamp 18001
transform 1 0 19964 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout102_A
timestamp 18001
transform 1 0 27508 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout104_A
timestamp 18001
transform 1 0 23552 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout105_A
timestamp 18001
transform -1 0 18216 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout105_X
timestamp 18001
transform 1 0 19780 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout106_A
timestamp 18001
transform -1 0 21068 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout107_A
timestamp 18001
transform 1 0 18032 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout108_A
timestamp 18001
transform 1 0 19688 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout108_X
timestamp 18001
transform 1 0 20240 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout109_A
timestamp 18001
transform 1 0 27968 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout110_A
timestamp 18001
transform 1 0 30636 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout112_A
timestamp 18001
transform 1 0 28060 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout113_A
timestamp 18001
transform -1 0 18584 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout113_X
timestamp 18001
transform 1 0 18584 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout116_A
timestamp 18001
transform 1 0 36708 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout117_A
timestamp 18001
transform 1 0 53268 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout118_A
timestamp 18001
transform 1 0 46184 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout119_A
timestamp 18001
transform -1 0 35052 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout120_A
timestamp 18001
transform 1 0 43056 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout121_A
timestamp 18001
transform 1 0 36708 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout121_X
timestamp 18001
transform 1 0 36524 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout123_A
timestamp 18001
transform 1 0 49680 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout124_A
timestamp 18001
transform 1 0 49312 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout124_X
timestamp 18001
transform 1 0 49496 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout125_A
timestamp 18001
transform -1 0 36708 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout125_X
timestamp 18001
transform 1 0 37260 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 18001
transform -1 0 19412 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 18001
transform -1 0 29164 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 18001
transform -1 0 28428 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 18001
transform -1 0 31648 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 18001
transform -1 0 31464 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 18001
transform -1 0 1840 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk
timestamp 18001
transform -1 0 36800 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_clk
timestamp 18001
transform -1 0 26404 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_clk
timestamp 18001
transform 1 0 45540 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_0_clk
timestamp 18001
transform 1 0 16652 0 -1 18496
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_1_clk
timestamp 18001
transform 1 0 23276 0 1 15232
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_2_clk
timestamp 18001
transform 1 0 29992 0 1 19584
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_3_clk
timestamp 18001
transform 1 0 21988 0 -1 23936
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_4_clk
timestamp 18001
transform 1 0 18308 0 -1 22848
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_5_clk
timestamp 18001
transform 1 0 16376 0 1 31552
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_6_clk
timestamp 18001
transform 1 0 24656 0 1 33728
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_7_clk
timestamp 18001
transform 1 0 30636 0 -1 31552
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_8_clk
timestamp 18001
transform 1 0 29532 0 1 27200
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_9_clk
timestamp 18001
transform -1 0 35880 0 1 23936
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_10_clk
timestamp 18001
transform -1 0 38640 0 -1 30464
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_11_clk
timestamp 18001
transform 1 0 50232 0 -1 28288
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_12_clk
timestamp 18001
transform 1 0 54188 0 1 22848
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_13_clk
timestamp 18001
transform 1 0 46368 0 1 23936
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_14_clk
timestamp 18001
transform 1 0 40756 0 -1 19584
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_15_clk
timestamp 18001
transform 1 0 46552 0 1 16320
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_16_clk
timestamp 18001
transform 1 0 55292 0 1 16320
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_17_clk
timestamp 18001
transform 1 0 49036 0 1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_18_clk
timestamp 18001
transform -1 0 40848 0 1 7616
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_19_clk
timestamp 18001
transform 1 0 40020 0 1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_20_clk
timestamp 18001
transform 1 0 32384 0 -1 16320
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_21_clk
timestamp 18001
transform 1 0 27784 0 1 9792
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_22_clk
timestamp 18001
transform -1 0 28888 0 1 4352
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_23_clk
timestamp 18001
transform 1 0 21988 0 -1 7616
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_24_clk
timestamp 18001
transform -1 0 16100 0 -1 7616
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_leaf_25_clk
timestamp 18001
transform 1 0 15364 0 1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__inv_8  clkload0
timestamp 18001
transform 1 0 45540 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkinv_8  clkload1
timestamp 18001
transform 1 0 16468 0 1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__bufinv_16  clkload2
timestamp 18001
transform 1 0 23368 0 -1 15232
box -38 -48 2246 592
use sky130_fd_sc_hd__inv_4  clkload3
timestamp 18001
transform 1 0 30176 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__inv_6  clkload4
timestamp 18001
transform 1 0 21068 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__inv_12  clkload5
timestamp 18001
transform 1 0 17940 0 1 22848
box -38 -48 1234 592
use sky130_fd_sc_hd__clkinv_8  clkload6
timestamp 18001
transform 1 0 16652 0 -1 32640
box -38 -48 1234 592
use sky130_fd_sc_hd__clkinv_2  clkload7
timestamp 18001
transform 1 0 23920 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_8  clkload8
timestamp 18001
transform 1 0 31372 0 1 31552
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_6  clkload9
timestamp 18001
transform 1 0 29532 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__inv_8  clkload10
timestamp 18001
transform 1 0 32384 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__inv_12  clkload11
timestamp 18001
transform 1 0 27784 0 -1 9792
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_8  clkload12
timestamp 18001
transform 1 0 21620 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkinv_4  clkload13
timestamp 18001
transform 1 0 15088 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__inv_8  clkload14
timestamp 18001
transform 1 0 15364 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__inv_4  clkload15
timestamp 18001
transform 1 0 34868 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__clkinvlp_4  clkload16
timestamp 18001
transform 1 0 38732 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__inv_6  clkload17
timestamp 18001
transform 1 0 49404 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_2  clkload18
timestamp 18001
transform 1 0 46000 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  clkload19
timestamp 18001
transform 1 0 40388 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_2  clkload20
timestamp 18001
transform 1 0 46184 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_8  clkload21
timestamp 18001
transform 1 0 54188 0 1 16320
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_8  clkload22
timestamp 18001
transform -1 0 50692 0 -1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_6  clkload23
timestamp 18001
transform 1 0 39008 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_4  clkload24
timestamp 18001
transform 1 0 41400 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  fanout22
timestamp 18001
transform -1 0 36984 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout23
timestamp 18001
transform -1 0 36616 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  fanout24
timestamp 18001
transform -1 0 29348 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout25
timestamp 18001
transform -1 0 28980 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout26
timestamp 18001
transform -1 0 35696 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout27
timestamp 18001
transform -1 0 38364 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout28
timestamp 18001
transform 1 0 37812 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout29
timestamp 18001
transform -1 0 49036 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout30
timestamp 18001
transform 1 0 52072 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout31
timestamp 18001
transform 1 0 38180 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout32
timestamp 18001
transform 1 0 38640 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout33
timestamp 18001
transform 1 0 38548 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout34
timestamp 18001
transform -1 0 39468 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout35
timestamp 18001
transform -1 0 28152 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout36
timestamp 18001
transform -1 0 24288 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout37
timestamp 18001
transform 1 0 33856 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout38
timestamp 18001
transform 1 0 46460 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout39
timestamp 18001
transform 1 0 46920 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout40
timestamp 18001
transform 1 0 33120 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout41
timestamp 18001
transform -1 0 24748 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout42
timestamp 18001
transform -1 0 27324 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout43
timestamp 18001
transform 1 0 23552 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout44
timestamp 18001
transform -1 0 27140 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout45
timestamp 18001
transform 1 0 36616 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout46
timestamp 18001
transform 1 0 32752 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout47
timestamp 18001
transform 1 0 36432 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout48
timestamp 18001
transform -1 0 36800 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout49
timestamp 18001
transform -1 0 38088 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout50
timestamp 18001
transform 1 0 43424 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout51
timestamp 18001
transform -1 0 39284 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout52
timestamp 18001
transform 1 0 52716 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout53
timestamp 18001
transform -1 0 52532 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout54
timestamp 18001
transform 1 0 47564 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout55
timestamp 18001
transform 1 0 55292 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout56
timestamp 18001
transform 1 0 39192 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout57
timestamp 18001
transform 1 0 25668 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout58
timestamp 18001
transform 1 0 31004 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  fanout59
timestamp 18001
transform 1 0 47564 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout60
timestamp 18001
transform -1 0 24748 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout61
timestamp 18001
transform -1 0 26956 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout62
timestamp 18001
transform 1 0 24472 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout63
timestamp 18001
transform -1 0 26312 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout64
timestamp 18001
transform 1 0 35788 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout65
timestamp 18001
transform -1 0 37812 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout66
timestamp 18001
transform 1 0 35512 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  fanout67
timestamp 18001
transform -1 0 37444 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout68
timestamp 18001
transform 1 0 45908 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout69
timestamp 18001
transform -1 0 47380 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout70
timestamp 18001
transform 1 0 55844 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout71
timestamp 18001
transform 1 0 54188 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout72
timestamp 18001
transform -1 0 52440 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout73
timestamp 18001
transform -1 0 56304 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout74
timestamp 18001
transform 1 0 54924 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  fanout75
timestamp 18001
transform -1 0 29440 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout76
timestamp 18001
transform -1 0 29164 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout77
timestamp 18001
transform 1 0 23000 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout78
timestamp 18001
transform -1 0 27232 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout79
timestamp 18001
transform 1 0 24104 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout80
timestamp 18001
transform 1 0 29532 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout81
timestamp 18001
transform -1 0 26956 0 1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  fanout82
timestamp 18001
transform 1 0 30268 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout83
timestamp 18001
transform 1 0 32752 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout84
timestamp 18001
transform 1 0 29900 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout85
timestamp 18001
transform -1 0 39652 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout86
timestamp 18001
transform -1 0 43700 0 1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  fanout87
timestamp 18001
transform 1 0 39008 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout88
timestamp 18001
transform -1 0 50048 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout89
timestamp 18001
transform -1 0 52164 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout90
timestamp 18001
transform 1 0 49128 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout91
timestamp 18001
transform 1 0 52440 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout92
timestamp 18001
transform 1 0 38640 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout93
timestamp 18001
transform 1 0 37260 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout94
timestamp 18001
transform 1 0 26956 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout95
timestamp 18001
transform 1 0 20332 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout96
timestamp 18001
transform -1 0 18952 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout97
timestamp 18001
transform -1 0 20516 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout98
timestamp 18001
transform 1 0 20424 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout99
timestamp 18001
transform -1 0 18584 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout100
timestamp 18001
transform -1 0 19780 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout101
timestamp 18001
transform -1 0 28244 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout102
timestamp 18001
transform 1 0 26956 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout103
timestamp 18001
transform 1 0 30176 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout104
timestamp 18001
transform 1 0 23736 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout105
timestamp 18001
transform 1 0 19044 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout106
timestamp 18001
transform -1 0 20884 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout107
timestamp 18001
transform -1 0 17940 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout108
timestamp 18001
transform 1 0 19872 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout109
timestamp 18001
transform 1 0 27416 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout110
timestamp 18001
transform 1 0 30820 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout111
timestamp 18001
transform -1 0 27508 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout112
timestamp 18001
transform -1 0 28060 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout113
timestamp 18001
transform 1 0 18768 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout114
timestamp 18001
transform 1 0 36708 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout115
timestamp 18001
transform 1 0 41952 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout116
timestamp 18001
transform -1 0 36708 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout117
timestamp 18001
transform 1 0 52716 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout118
timestamp 18001
transform -1 0 46920 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout119
timestamp 18001
transform 1 0 35052 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout120
timestamp 18001
transform -1 0 43056 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout121
timestamp 18001
transform -1 0 36524 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout122
timestamp 18001
transform 1 0 52716 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout123
timestamp 18001
transform -1 0 49128 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout124
timestamp 18001
transform -1 0 49312 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout125
timestamp 18001
transform 1 0 36708 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_3
timestamp 1636986456
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_15
timestamp 1636986456
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27
timestamp 18001
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29
timestamp 1636986456
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_41
timestamp 1636986456
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_53
timestamp 18001
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_57
timestamp 1636986456
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_69
timestamp 1636986456
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_81
timestamp 18001
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_85
timestamp 1636986456
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_97
timestamp 1636986456
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_109
timestamp 18001
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_113
timestamp 1636986456
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_125
timestamp 1636986456
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_137
timestamp 18001
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_141
timestamp 1636986456
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_153
timestamp 1636986456
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_165
timestamp 18001
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_169
timestamp 1636986456
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_181
timestamp 1636986456
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_193
timestamp 18001
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_202
timestamp 18001
transform 1 0 19688 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_210
timestamp 18001
transform 1 0 20424 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_217
timestamp 18001
transform 1 0 21068 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_225
timestamp 18001
transform 1 0 21804 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_239
timestamp 18001
transform 1 0 23092 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_245
timestamp 18001
transform 1 0 23644 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_251
timestamp 18001
transform 1 0 24196 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_253
timestamp 1636986456
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_265
timestamp 1636986456
transform 1 0 25484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_277
timestamp 18001
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_281
timestamp 1636986456
transform 1 0 26956 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_293
timestamp 18001
transform 1 0 28060 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_332
timestamp 18001
transform 1 0 31648 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_337
timestamp 1636986456
transform 1 0 32108 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_349
timestamp 1636986456
transform 1 0 33212 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_361
timestamp 18001
transform 1 0 34316 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_365
timestamp 18001
transform 1 0 34684 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_371
timestamp 18001
transform 1 0 35236 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_375
timestamp 1636986456
transform 1 0 35604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_387
timestamp 18001
transform 1 0 36708 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_391
timestamp 18001
transform 1 0 37076 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_396
timestamp 1636986456
transform 1 0 37536 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_408
timestamp 1636986456
transform 1 0 38640 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_421
timestamp 1636986456
transform 1 0 39836 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_433
timestamp 1636986456
transform 1 0 40940 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_445
timestamp 18001
transform 1 0 42044 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_452
timestamp 18001
transform 1 0 42688 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_460
timestamp 18001
transform 1 0 43424 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_465
timestamp 18001
transform 1 0 43884 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_473
timestamp 18001
transform 1 0 44620 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_477
timestamp 1636986456
transform 1 0 44988 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_489
timestamp 1636986456
transform 1 0 46092 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_501
timestamp 18001
transform 1 0 47196 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_505
timestamp 1636986456
transform 1 0 47564 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_517
timestamp 1636986456
transform 1 0 48668 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_529
timestamp 18001
transform 1 0 49772 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_533
timestamp 1636986456
transform 1 0 50140 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_545
timestamp 1636986456
transform 1 0 51244 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_557
timestamp 18001
transform 1 0 52348 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_561
timestamp 1636986456
transform 1 0 52716 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_573
timestamp 1636986456
transform 1 0 53820 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_585
timestamp 18001
transform 1 0 54924 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_589
timestamp 1636986456
transform 1 0 55292 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_601
timestamp 1636986456
transform 1 0 56396 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_613
timestamp 18001
transform 1 0 57500 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_617
timestamp 18001
transform 1 0 57868 0 1 2176
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1636986456
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 1636986456
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 1636986456
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_39
timestamp 1636986456
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_51
timestamp 18001
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 18001
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_57
timestamp 1636986456
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_69
timestamp 1636986456
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_81
timestamp 1636986456
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_93
timestamp 1636986456
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_105
timestamp 18001
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_111
timestamp 18001
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_113
timestamp 1636986456
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_125
timestamp 1636986456
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_137
timestamp 1636986456
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_149
timestamp 1636986456
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_161
timestamp 18001
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_167
timestamp 18001
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_169
timestamp 1636986456
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_181
timestamp 1636986456
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_193
timestamp 1636986456
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_205
timestamp 18001
transform 1 0 19964 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_213
timestamp 18001
transform 1 0 20700 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_220
timestamp 18001
transform 1 0 21344 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_247
timestamp 18001
transform 1 0 23828 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_268
timestamp 1636986456
transform 1 0 25760 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_281
timestamp 1636986456
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_335
timestamp 18001
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_358
timestamp 18001
transform 1 0 34040 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_370
timestamp 18001
transform 1 0 35144 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_397
timestamp 18001
transform 1 0 37628 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_453
timestamp 18001
transform 1 0 42780 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_466
timestamp 18001
transform 1 0 43976 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_481
timestamp 1636986456
transform 1 0 45356 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_493
timestamp 18001
transform 1 0 46460 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_501
timestamp 18001
transform 1 0 47196 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_505
timestamp 1636986456
transform 1 0 47564 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_517
timestamp 1636986456
transform 1 0 48668 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_529
timestamp 1636986456
transform 1 0 49772 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_541
timestamp 1636986456
transform 1 0 50876 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_553
timestamp 18001
transform 1 0 51980 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_559
timestamp 18001
transform 1 0 52532 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_561
timestamp 1636986456
transform 1 0 52716 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_573
timestamp 1636986456
transform 1 0 53820 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_585
timestamp 1636986456
transform 1 0 54924 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_597
timestamp 1636986456
transform 1 0 56028 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_609
timestamp 18001
transform 1 0 57132 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_615
timestamp 18001
transform 1 0 57684 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_617
timestamp 18001
transform 1 0 57868 0 -1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1636986456
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1636986456
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 18001
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1636986456
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 1636986456
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_53
timestamp 1636986456
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_65
timestamp 1636986456
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_77
timestamp 18001
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 18001
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_85
timestamp 1636986456
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_97
timestamp 1636986456
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_109
timestamp 1636986456
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_121
timestamp 1636986456
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_133
timestamp 18001
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 18001
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_141
timestamp 1636986456
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_153
timestamp 1636986456
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_165
timestamp 1636986456
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_177
timestamp 1636986456
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_189
timestamp 18001
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_195
timestamp 18001
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_197
timestamp 18001
transform 1 0 19228 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_201
timestamp 18001
transform 1 0 19596 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_222
timestamp 18001
transform 1 0 21528 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_239
timestamp 18001
transform 1 0 23092 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_246
timestamp 18001
transform 1 0 23736 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_253
timestamp 18001
transform 1 0 24380 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_264
timestamp 18001
transform 1 0 25392 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_271
timestamp 18001
transform 1 0 26036 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_294
timestamp 18001
transform 1 0 28152 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_300
timestamp 18001
transform 1 0 28704 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_309
timestamp 18001
transform 1 0 29532 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_320
timestamp 18001
transform 1 0 30544 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_342
timestamp 1636986456
transform 1 0 32568 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_354
timestamp 18001
transform 1 0 33672 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_362
timestamp 18001
transform 1 0 34408 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_365
timestamp 1636986456
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_377
timestamp 1636986456
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_389
timestamp 1636986456
transform 1 0 36892 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_401
timestamp 1636986456
transform 1 0 37996 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_413
timestamp 18001
transform 1 0 39100 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_419
timestamp 18001
transform 1 0 39652 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_421
timestamp 1636986456
transform 1 0 39836 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_433
timestamp 1636986456
transform 1 0 40940 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_445
timestamp 1636986456
transform 1 0 42044 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_457
timestamp 1636986456
transform 1 0 43148 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_469
timestamp 18001
transform 1 0 44252 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_475
timestamp 18001
transform 1 0 44804 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_477
timestamp 1636986456
transform 1 0 44988 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_489
timestamp 1636986456
transform 1 0 46092 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_501
timestamp 1636986456
transform 1 0 47196 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_513
timestamp 1636986456
transform 1 0 48300 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_525
timestamp 18001
transform 1 0 49404 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_531
timestamp 18001
transform 1 0 49956 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_533
timestamp 1636986456
transform 1 0 50140 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_545
timestamp 1636986456
transform 1 0 51244 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_557
timestamp 1636986456
transform 1 0 52348 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_569
timestamp 1636986456
transform 1 0 53452 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_581
timestamp 18001
transform 1 0 54556 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_587
timestamp 18001
transform 1 0 55108 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_589
timestamp 1636986456
transform 1 0 55292 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_601
timestamp 1636986456
transform 1 0 56396 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_613
timestamp 1636986456
transform 1 0 57500 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1636986456
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1636986456
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 1636986456
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 1636986456
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 18001
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 18001
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1636986456
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_69
timestamp 1636986456
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_81
timestamp 1636986456
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_93
timestamp 1636986456
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_105
timestamp 18001
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 18001
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_113
timestamp 1636986456
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_125
timestamp 1636986456
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_137
timestamp 1636986456
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_149
timestamp 1636986456
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_161
timestamp 18001
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_167
timestamp 18001
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_177
timestamp 1636986456
transform 1 0 17388 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_189
timestamp 1636986456
transform 1 0 18492 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_201
timestamp 18001
transform 1 0 19596 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_223
timestamp 18001
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_242
timestamp 18001
transform 1 0 23368 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_263
timestamp 18001
transform 1 0 25300 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_277
timestamp 18001
transform 1 0 26588 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_302
timestamp 1636986456
transform 1 0 28888 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_314
timestamp 1636986456
transform 1 0 29992 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_326
timestamp 18001
transform 1 0 31096 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_334
timestamp 18001
transform 1 0 31832 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_337
timestamp 1636986456
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_349
timestamp 1636986456
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_361
timestamp 1636986456
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_373
timestamp 1636986456
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_385
timestamp 18001
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_391
timestamp 18001
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_393
timestamp 1636986456
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_405
timestamp 1636986456
transform 1 0 38364 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_417
timestamp 1636986456
transform 1 0 39468 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_429
timestamp 1636986456
transform 1 0 40572 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_441
timestamp 18001
transform 1 0 41676 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_447
timestamp 18001
transform 1 0 42228 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_449
timestamp 1636986456
transform 1 0 42412 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_461
timestamp 1636986456
transform 1 0 43516 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_473
timestamp 1636986456
transform 1 0 44620 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_485
timestamp 1636986456
transform 1 0 45724 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_497
timestamp 18001
transform 1 0 46828 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_503
timestamp 18001
transform 1 0 47380 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_505
timestamp 1636986456
transform 1 0 47564 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_517
timestamp 1636986456
transform 1 0 48668 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_529
timestamp 1636986456
transform 1 0 49772 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_541
timestamp 1636986456
transform 1 0 50876 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_553
timestamp 18001
transform 1 0 51980 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_559
timestamp 18001
transform 1 0 52532 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_561
timestamp 1636986456
transform 1 0 52716 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_573
timestamp 1636986456
transform 1 0 53820 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_585
timestamp 1636986456
transform 1 0 54924 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_597
timestamp 1636986456
transform 1 0 56028 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_609
timestamp 18001
transform 1 0 57132 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_615
timestamp 18001
transform 1 0 57684 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_617
timestamp 18001
transform 1 0 57868 0 -1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1636986456
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1636986456
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 18001
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1636986456
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 1636986456
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_53
timestamp 1636986456
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_65
timestamp 1636986456
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_77
timestamp 18001
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 18001
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_85
timestamp 1636986456
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_97
timestamp 1636986456
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_109
timestamp 1636986456
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_121
timestamp 1636986456
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_133
timestamp 18001
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_139
timestamp 18001
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_141
timestamp 1636986456
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_153
timestamp 18001
transform 1 0 15180 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_177
timestamp 1636986456
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_189
timestamp 18001
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_195
timestamp 18001
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_197
timestamp 1636986456
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_209
timestamp 18001
transform 1 0 20332 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_220
timestamp 1636986456
transform 1 0 21344 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_232
timestamp 18001
transform 1 0 22448 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_241
timestamp 18001
transform 1 0 23276 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_247
timestamp 18001
transform 1 0 23828 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_251
timestamp 18001
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_274
timestamp 1636986456
transform 1 0 26312 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_286
timestamp 18001
transform 1 0 27416 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_302
timestamp 18001
transform 1 0 28888 0 1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_309
timestamp 1636986456
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_321
timestamp 18001
transform 1 0 30636 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_326
timestamp 18001
transform 1 0 31096 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_350
timestamp 1636986456
transform 1 0 33304 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_385
timestamp 1636986456
transform 1 0 36524 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_397
timestamp 1636986456
transform 1 0 37628 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_409
timestamp 18001
transform 1 0 38732 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_417
timestamp 18001
transform 1 0 39468 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_421
timestamp 1636986456
transform 1 0 39836 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_433
timestamp 1636986456
transform 1 0 40940 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_445
timestamp 1636986456
transform 1 0 42044 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_457
timestamp 1636986456
transform 1 0 43148 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_469
timestamp 18001
transform 1 0 44252 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_475
timestamp 18001
transform 1 0 44804 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_477
timestamp 1636986456
transform 1 0 44988 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_489
timestamp 1636986456
transform 1 0 46092 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_501
timestamp 1636986456
transform 1 0 47196 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_513
timestamp 1636986456
transform 1 0 48300 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_525
timestamp 18001
transform 1 0 49404 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_531
timestamp 18001
transform 1 0 49956 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_533
timestamp 1636986456
transform 1 0 50140 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_545
timestamp 1636986456
transform 1 0 51244 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_557
timestamp 1636986456
transform 1 0 52348 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_569
timestamp 1636986456
transform 1 0 53452 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_581
timestamp 18001
transform 1 0 54556 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_587
timestamp 18001
transform 1 0 55108 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_589
timestamp 1636986456
transform 1 0 55292 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_601
timestamp 1636986456
transform 1 0 56396 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_613
timestamp 1636986456
transform 1 0 57500 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1636986456
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 1636986456
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_27
timestamp 1636986456
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_39
timestamp 1636986456
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_51
timestamp 18001
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 18001
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 1636986456
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_69
timestamp 1636986456
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_81
timestamp 1636986456
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_93
timestamp 1636986456
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_105
timestamp 18001
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_111
timestamp 18001
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_113
timestamp 1636986456
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_125
timestamp 18001
transform 1 0 12604 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_147
timestamp 18001
transform 1 0 14628 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_172
timestamp 1636986456
transform 1 0 16928 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_184
timestamp 1636986456
transform 1 0 18032 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_196
timestamp 18001
transform 1 0 19136 0 -1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_212
timestamp 1636986456
transform 1 0 20608 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_225
timestamp 1636986456
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_237
timestamp 18001
transform 1 0 22908 0 -1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_266
timestamp 1636986456
transform 1 0 25576 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_278
timestamp 18001
transform 1 0 26680 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_281
timestamp 18001
transform 1 0 26956 0 -1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_309
timestamp 1636986456
transform 1 0 29532 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_321
timestamp 18001
transform 1 0 30636 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_335
timestamp 18001
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_337
timestamp 1636986456
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_349
timestamp 18001
transform 1 0 33212 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_367
timestamp 18001
transform 1 0 34868 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_373
timestamp 18001
transform 1 0 35420 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_390
timestamp 18001
transform 1 0 36984 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_393
timestamp 1636986456
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_405
timestamp 1636986456
transform 1 0 38364 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_417
timestamp 1636986456
transform 1 0 39468 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_429
timestamp 1636986456
transform 1 0 40572 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_441
timestamp 18001
transform 1 0 41676 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_447
timestamp 18001
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_449
timestamp 1636986456
transform 1 0 42412 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_461
timestamp 1636986456
transform 1 0 43516 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_473
timestamp 1636986456
transform 1 0 44620 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_485
timestamp 1636986456
transform 1 0 45724 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_497
timestamp 18001
transform 1 0 46828 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_503
timestamp 18001
transform 1 0 47380 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_505
timestamp 1636986456
transform 1 0 47564 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_517
timestamp 1636986456
transform 1 0 48668 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_529
timestamp 1636986456
transform 1 0 49772 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_541
timestamp 1636986456
transform 1 0 50876 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_553
timestamp 18001
transform 1 0 51980 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_559
timestamp 18001
transform 1 0 52532 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_561
timestamp 1636986456
transform 1 0 52716 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_573
timestamp 1636986456
transform 1 0 53820 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_585
timestamp 1636986456
transform 1 0 54924 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_597
timestamp 1636986456
transform 1 0 56028 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_609
timestamp 18001
transform 1 0 57132 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_615
timestamp 18001
transform 1 0 57684 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_617
timestamp 18001
transform 1 0 57868 0 -1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 1636986456
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 1636986456
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 18001
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 1636986456
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_41
timestamp 1636986456
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_53
timestamp 1636986456
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_65
timestamp 1636986456
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_77
timestamp 18001
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 18001
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_85
timestamp 1636986456
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_97
timestamp 1636986456
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_109
timestamp 1636986456
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_121
timestamp 18001
transform 1 0 12236 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_130
timestamp 18001
transform 1 0 13064 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_138
timestamp 18001
transform 1 0 13800 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_157
timestamp 18001
transform 1 0 15548 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_170
timestamp 18001
transform 1 0 16744 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_178
timestamp 18001
transform 1 0 17480 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_195
timestamp 18001
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_222
timestamp 1636986456
transform 1 0 21528 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_234
timestamp 1636986456
transform 1 0 22632 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_246
timestamp 18001
transform 1 0 23736 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_253
timestamp 1636986456
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_265
timestamp 18001
transform 1 0 25484 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_307
timestamp 18001
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_311
timestamp 18001
transform 1 0 29716 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_343
timestamp 18001
transform 1 0 32660 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_373
timestamp 18001
transform 1 0 35420 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_377
timestamp 18001
transform 1 0 35788 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_401
timestamp 1636986456
transform 1 0 37996 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_413
timestamp 18001
transform 1 0 39100 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_419
timestamp 18001
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_421
timestamp 1636986456
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_433
timestamp 1636986456
transform 1 0 40940 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_445
timestamp 1636986456
transform 1 0 42044 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_457
timestamp 1636986456
transform 1 0 43148 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_469
timestamp 18001
transform 1 0 44252 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_475
timestamp 18001
transform 1 0 44804 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_477
timestamp 1636986456
transform 1 0 44988 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_489
timestamp 1636986456
transform 1 0 46092 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_501
timestamp 1636986456
transform 1 0 47196 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_513
timestamp 1636986456
transform 1 0 48300 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_525
timestamp 18001
transform 1 0 49404 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_531
timestamp 18001
transform 1 0 49956 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_533
timestamp 1636986456
transform 1 0 50140 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_545
timestamp 1636986456
transform 1 0 51244 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_557
timestamp 1636986456
transform 1 0 52348 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_569
timestamp 1636986456
transform 1 0 53452 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_581
timestamp 18001
transform 1 0 54556 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_587
timestamp 18001
transform 1 0 55108 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_589
timestamp 1636986456
transform 1 0 55292 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_601
timestamp 1636986456
transform 1 0 56396 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_613
timestamp 1636986456
transform 1 0 57500 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1636986456
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 1636986456
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_27
timestamp 1636986456
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_39
timestamp 1636986456
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_51
timestamp 18001
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 18001
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_57
timestamp 1636986456
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_69
timestamp 1636986456
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_81
timestamp 1636986456
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_93
timestamp 1636986456
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_105
timestamp 18001
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_111
timestamp 18001
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_113
timestamp 18001
transform 1 0 11500 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_142
timestamp 18001
transform 1 0 14168 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_163
timestamp 18001
transform 1 0 16100 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_167
timestamp 18001
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_169
timestamp 18001
transform 1 0 16652 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_200
timestamp 18001
transform 1 0 19504 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_205
timestamp 18001
transform 1 0 19964 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_223
timestamp 18001
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_245
timestamp 1636986456
transform 1 0 23644 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_257
timestamp 1636986456
transform 1 0 24748 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_269
timestamp 18001
transform 1 0 25852 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_277
timestamp 18001
transform 1 0 26588 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_281
timestamp 18001
transform 1 0 26956 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_297
timestamp 18001
transform 1 0 28428 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_313
timestamp 18001
transform 1 0 29900 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_330
timestamp 18001
transform 1 0 31464 0 -1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_337
timestamp 1636986456
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_349
timestamp 18001
transform 1 0 33212 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_358
timestamp 1636986456
transform 1 0 34040 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_370
timestamp 18001
transform 1 0 35144 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_391
timestamp 18001
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_393
timestamp 1636986456
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_405
timestamp 1636986456
transform 1 0 38364 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_417
timestamp 1636986456
transform 1 0 39468 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_429
timestamp 1636986456
transform 1 0 40572 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_441
timestamp 18001
transform 1 0 41676 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_447
timestamp 18001
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_449
timestamp 1636986456
transform 1 0 42412 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_461
timestamp 1636986456
transform 1 0 43516 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_473
timestamp 1636986456
transform 1 0 44620 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_485
timestamp 1636986456
transform 1 0 45724 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_497
timestamp 18001
transform 1 0 46828 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_503
timestamp 18001
transform 1 0 47380 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_505
timestamp 1636986456
transform 1 0 47564 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_517
timestamp 1636986456
transform 1 0 48668 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_529
timestamp 1636986456
transform 1 0 49772 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_541
timestamp 1636986456
transform 1 0 50876 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_553
timestamp 18001
transform 1 0 51980 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_559
timestamp 18001
transform 1 0 52532 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_561
timestamp 1636986456
transform 1 0 52716 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_573
timestamp 1636986456
transform 1 0 53820 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_585
timestamp 1636986456
transform 1 0 54924 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_597
timestamp 1636986456
transform 1 0 56028 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_609
timestamp 18001
transform 1 0 57132 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_615
timestamp 18001
transform 1 0 57684 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_617
timestamp 18001
transform 1 0 57868 0 -1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1636986456
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 1636986456
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 18001
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 1636986456
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_41
timestamp 1636986456
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_53
timestamp 1636986456
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_65
timestamp 1636986456
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_77
timestamp 18001
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_83
timestamp 18001
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_85
timestamp 1636986456
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_97
timestamp 1636986456
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_109
timestamp 1636986456
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_121
timestamp 1636986456
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_133
timestamp 18001
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_139
timestamp 18001
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_149
timestamp 1636986456
transform 1 0 14812 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_170
timestamp 1636986456
transform 1 0 16744 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_182
timestamp 18001
transform 1 0 17848 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_190
timestamp 18001
transform 1 0 18584 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_197
timestamp 1636986456
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_253
timestamp 18001
transform 1 0 24380 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_261
timestamp 18001
transform 1 0 25116 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_289
timestamp 1636986456
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_301
timestamp 18001
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_307
timestamp 18001
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_309
timestamp 18001
transform 1 0 29532 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_317
timestamp 18001
transform 1 0 30268 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_325
timestamp 1636986456
transform 1 0 31004 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_337
timestamp 18001
transform 1 0 32108 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_350
timestamp 18001
transform 1 0 33304 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_358
timestamp 18001
transform 1 0 34040 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_363
timestamp 18001
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_365
timestamp 18001
transform 1 0 34684 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_377
timestamp 18001
transform 1 0 35788 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_381
timestamp 18001
transform 1 0 36156 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_386
timestamp 18001
transform 1 0 36616 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_390
timestamp 1636986456
transform 1 0 36984 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_402
timestamp 1636986456
transform 1 0 38088 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_414
timestamp 18001
transform 1 0 39192 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_421
timestamp 1636986456
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_433
timestamp 1636986456
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_445
timestamp 1636986456
transform 1 0 42044 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_457
timestamp 1636986456
transform 1 0 43148 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_469
timestamp 18001
transform 1 0 44252 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_475
timestamp 18001
transform 1 0 44804 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_477
timestamp 1636986456
transform 1 0 44988 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_489
timestamp 1636986456
transform 1 0 46092 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_501
timestamp 1636986456
transform 1 0 47196 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_513
timestamp 1636986456
transform 1 0 48300 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_525
timestamp 18001
transform 1 0 49404 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_531
timestamp 18001
transform 1 0 49956 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_533
timestamp 1636986456
transform 1 0 50140 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_545
timestamp 1636986456
transform 1 0 51244 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_557
timestamp 1636986456
transform 1 0 52348 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_569
timestamp 1636986456
transform 1 0 53452 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_581
timestamp 18001
transform 1 0 54556 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_587
timestamp 18001
transform 1 0 55108 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_589
timestamp 1636986456
transform 1 0 55292 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_601
timestamp 1636986456
transform 1 0 56396 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_613
timestamp 1636986456
transform 1 0 57500 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 1636986456
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_15
timestamp 1636986456
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_27
timestamp 1636986456
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_39
timestamp 1636986456
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_51
timestamp 18001
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_55
timestamp 18001
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_57
timestamp 1636986456
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_69
timestamp 1636986456
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_81
timestamp 1636986456
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_93
timestamp 1636986456
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_105
timestamp 18001
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_111
timestamp 18001
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_113
timestamp 18001
transform 1 0 11500 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_121
timestamp 18001
transform 1 0 12236 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_130
timestamp 18001
transform 1 0 13064 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_142
timestamp 18001
transform 1 0 14168 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_150
timestamp 18001
transform 1 0 14904 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_167
timestamp 18001
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_180
timestamp 1636986456
transform 1 0 17664 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_192
timestamp 1636986456
transform 1 0 18768 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_204
timestamp 18001
transform 1 0 19872 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_214
timestamp 18001
transform 1 0 20792 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_221
timestamp 18001
transform 1 0 21436 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_225
timestamp 18001
transform 1 0 21804 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_243
timestamp 1636986456
transform 1 0 23460 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_255
timestamp 1636986456
transform 1 0 24564 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_267
timestamp 18001
transform 1 0 25668 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_279
timestamp 18001
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_300
timestamp 18001
transform 1 0 28704 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_308
timestamp 18001
transform 1 0 29440 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_320
timestamp 18001
transform 1 0 30544 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_329
timestamp 18001
transform 1 0 31372 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_333
timestamp 18001
transform 1 0 31740 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_365
timestamp 18001
transform 1 0 34684 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_369
timestamp 18001
transform 1 0 35052 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_383
timestamp 18001
transform 1 0 36340 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_414
timestamp 1636986456
transform 1 0 39192 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_426
timestamp 1636986456
transform 1 0 40296 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_438
timestamp 18001
transform 1 0 41400 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_446
timestamp 18001
transform 1 0 42136 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_449
timestamp 1636986456
transform 1 0 42412 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_461
timestamp 1636986456
transform 1 0 43516 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_473
timestamp 1636986456
transform 1 0 44620 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_485
timestamp 1636986456
transform 1 0 45724 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_497
timestamp 18001
transform 1 0 46828 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_503
timestamp 18001
transform 1 0 47380 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_505
timestamp 1636986456
transform 1 0 47564 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_517
timestamp 1636986456
transform 1 0 48668 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_529
timestamp 1636986456
transform 1 0 49772 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_541
timestamp 1636986456
transform 1 0 50876 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_553
timestamp 18001
transform 1 0 51980 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_559
timestamp 18001
transform 1 0 52532 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_561
timestamp 1636986456
transform 1 0 52716 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_573
timestamp 1636986456
transform 1 0 53820 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_585
timestamp 1636986456
transform 1 0 54924 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_597
timestamp 1636986456
transform 1 0 56028 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_609
timestamp 18001
transform 1 0 57132 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_615
timestamp 18001
transform 1 0 57684 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_617
timestamp 18001
transform 1 0 57868 0 -1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 1636986456
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_15
timestamp 1636986456
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 18001
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_29
timestamp 1636986456
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_41
timestamp 1636986456
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_53
timestamp 1636986456
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_65
timestamp 1636986456
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_77
timestamp 18001
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_83
timestamp 18001
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_85
timestamp 1636986456
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_97
timestamp 1636986456
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_109
timestamp 18001
transform 1 0 11132 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_117
timestamp 18001
transform 1 0 11868 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_186
timestamp 18001
transform 1 0 18216 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_194
timestamp 18001
transform 1 0 18952 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_197
timestamp 18001
transform 1 0 19228 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_210
timestamp 18001
transform 1 0 20424 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_220
timestamp 18001
transform 1 0 21344 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_227
timestamp 1636986456
transform 1 0 21988 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_239
timestamp 1636986456
transform 1 0 23092 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_251
timestamp 18001
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_253
timestamp 1636986456
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_265
timestamp 18001
transform 1 0 25484 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_289
timestamp 18001
transform 1 0 27692 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_304
timestamp 18001
transform 1 0 29072 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_329
timestamp 18001
transform 1 0 31372 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_333
timestamp 18001
transform 1 0 31740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_352
timestamp 1636986456
transform 1 0 33488 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_365
timestamp 1636986456
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_377
timestamp 18001
transform 1 0 35788 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_419
timestamp 18001
transform 1 0 39652 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_434
timestamp 1636986456
transform 1 0 41032 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_446
timestamp 1636986456
transform 1 0 42136 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_458
timestamp 1636986456
transform 1 0 43240 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_470
timestamp 18001
transform 1 0 44344 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_477
timestamp 1636986456
transform 1 0 44988 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_489
timestamp 1636986456
transform 1 0 46092 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_501
timestamp 1636986456
transform 1 0 47196 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_513
timestamp 1636986456
transform 1 0 48300 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_525
timestamp 18001
transform 1 0 49404 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_531
timestamp 18001
transform 1 0 49956 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_533
timestamp 1636986456
transform 1 0 50140 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_545
timestamp 1636986456
transform 1 0 51244 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_557
timestamp 1636986456
transform 1 0 52348 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_569
timestamp 1636986456
transform 1 0 53452 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_581
timestamp 18001
transform 1 0 54556 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_587
timestamp 18001
transform 1 0 55108 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_589
timestamp 1636986456
transform 1 0 55292 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_601
timestamp 1636986456
transform 1 0 56396 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_613
timestamp 1636986456
transform 1 0 57500 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_3
timestamp 1636986456
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_15
timestamp 1636986456
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_27
timestamp 1636986456
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_39
timestamp 1636986456
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_51
timestamp 18001
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_55
timestamp 18001
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_57
timestamp 1636986456
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_69
timestamp 1636986456
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_81
timestamp 1636986456
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_93
timestamp 1636986456
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_105
timestamp 18001
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_111
timestamp 18001
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_113
timestamp 1636986456
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_125
timestamp 1636986456
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_137
timestamp 1636986456
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_149
timestamp 18001
transform 1 0 14812 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_163
timestamp 18001
transform 1 0 16100 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_167
timestamp 18001
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_189
timestamp 18001
transform 1 0 18492 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_195
timestamp 18001
transform 1 0 19044 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_225
timestamp 18001
transform 1 0 21804 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_229
timestamp 18001
transform 1 0 22172 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_237
timestamp 18001
transform 1 0 22908 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_258
timestamp 18001
transform 1 0 24840 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_289
timestamp 18001
transform 1 0 27692 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_293
timestamp 18001
transform 1 0 28060 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_305
timestamp 1636986456
transform 1 0 29164 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_317
timestamp 18001
transform 1 0 30268 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_325
timestamp 18001
transform 1 0 31004 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_348
timestamp 1636986456
transform 1 0 33120 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_360
timestamp 1636986456
transform 1 0 34224 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_372
timestamp 18001
transform 1 0 35328 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_407
timestamp 18001
transform 1 0 38548 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_430
timestamp 1636986456
transform 1 0 40664 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_442
timestamp 18001
transform 1 0 41768 0 -1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_449
timestamp 1636986456
transform 1 0 42412 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_461
timestamp 1636986456
transform 1 0 43516 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_473
timestamp 1636986456
transform 1 0 44620 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_485
timestamp 1636986456
transform 1 0 45724 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_497
timestamp 18001
transform 1 0 46828 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_503
timestamp 18001
transform 1 0 47380 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_505
timestamp 1636986456
transform 1 0 47564 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_517
timestamp 1636986456
transform 1 0 48668 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_529
timestamp 1636986456
transform 1 0 49772 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_541
timestamp 1636986456
transform 1 0 50876 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_553
timestamp 18001
transform 1 0 51980 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_559
timestamp 18001
transform 1 0 52532 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_561
timestamp 1636986456
transform 1 0 52716 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_573
timestamp 1636986456
transform 1 0 53820 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_585
timestamp 1636986456
transform 1 0 54924 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_597
timestamp 1636986456
transform 1 0 56028 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_609
timestamp 18001
transform 1 0 57132 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_615
timestamp 18001
transform 1 0 57684 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_617
timestamp 18001
transform 1 0 57868 0 -1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_3
timestamp 1636986456
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_15
timestamp 1636986456
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 18001
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_29
timestamp 1636986456
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_41
timestamp 1636986456
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_53
timestamp 1636986456
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_65
timestamp 1636986456
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_77
timestamp 18001
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_83
timestamp 18001
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_85
timestamp 1636986456
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_97
timestamp 1636986456
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_109
timestamp 1636986456
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_121
timestamp 1636986456
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_133
timestamp 18001
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_139
timestamp 18001
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_141
timestamp 1636986456
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_153
timestamp 1636986456
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_165
timestamp 1636986456
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_185
timestamp 18001
transform 1 0 18124 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_193
timestamp 18001
transform 1 0 18860 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_197
timestamp 1636986456
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_215
timestamp 18001
transform 1 0 20884 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_223
timestamp 18001
transform 1 0 21620 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_249
timestamp 18001
transform 1 0 24012 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_253
timestamp 1636986456
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_265
timestamp 1636986456
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_277
timestamp 18001
transform 1 0 26588 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_283
timestamp 18001
transform 1 0 27140 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_303
timestamp 18001
transform 1 0 28980 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_307
timestamp 18001
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_309
timestamp 1636986456
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_321
timestamp 1636986456
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_333
timestamp 18001
transform 1 0 31740 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_344
timestamp 18001
transform 1 0 32752 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_352
timestamp 1636986456
transform 1 0 33488 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_365
timestamp 18001
transform 1 0 34684 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_371
timestamp 18001
transform 1 0 35236 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_395
timestamp 18001
transform 1 0 37444 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_399
timestamp 18001
transform 1 0 37812 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_421
timestamp 1636986456
transform 1 0 39836 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_433
timestamp 1636986456
transform 1 0 40940 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_445
timestamp 1636986456
transform 1 0 42044 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_457
timestamp 1636986456
transform 1 0 43148 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_469
timestamp 18001
transform 1 0 44252 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_475
timestamp 18001
transform 1 0 44804 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_477
timestamp 1636986456
transform 1 0 44988 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_489
timestamp 1636986456
transform 1 0 46092 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_501
timestamp 1636986456
transform 1 0 47196 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_513
timestamp 1636986456
transform 1 0 48300 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_525
timestamp 18001
transform 1 0 49404 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_531
timestamp 18001
transform 1 0 49956 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_533
timestamp 1636986456
transform 1 0 50140 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_545
timestamp 1636986456
transform 1 0 51244 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_557
timestamp 1636986456
transform 1 0 52348 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_569
timestamp 1636986456
transform 1 0 53452 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_581
timestamp 18001
transform 1 0 54556 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_587
timestamp 18001
transform 1 0 55108 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_589
timestamp 1636986456
transform 1 0 55292 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_601
timestamp 1636986456
transform 1 0 56396 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_613
timestamp 1636986456
transform 1 0 57500 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_3
timestamp 1636986456
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_15
timestamp 1636986456
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_27
timestamp 1636986456
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_39
timestamp 1636986456
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_51
timestamp 18001
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_55
timestamp 18001
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_57
timestamp 1636986456
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_69
timestamp 1636986456
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_81
timestamp 1636986456
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_93
timestamp 1636986456
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_105
timestamp 18001
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_111
timestamp 18001
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_113
timestamp 1636986456
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_125
timestamp 18001
transform 1 0 12604 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_129
timestamp 18001
transform 1 0 12972 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_150
timestamp 1636986456
transform 1 0 14904 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_162
timestamp 18001
transform 1 0 16008 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_169
timestamp 18001
transform 1 0 16652 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_173
timestamp 1636986456
transform 1 0 17020 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_185
timestamp 1636986456
transform 1 0 18124 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_197
timestamp 1636986456
transform 1 0 19228 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_209
timestamp 1636986456
transform 1 0 20332 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_221
timestamp 18001
transform 1 0 21436 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_245
timestamp 1636986456
transform 1 0 23644 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_257
timestamp 1636986456
transform 1 0 24748 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_269
timestamp 18001
transform 1 0 25852 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_277
timestamp 18001
transform 1 0 26588 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_281
timestamp 18001
transform 1 0 26956 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_289
timestamp 18001
transform 1 0 27692 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_308
timestamp 18001
transform 1 0 29440 0 -1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_319
timestamp 1636986456
transform 1 0 30452 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_331
timestamp 18001
transform 1 0 31556 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_335
timestamp 18001
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_337
timestamp 18001
transform 1 0 32108 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_360
timestamp 1636986456
transform 1 0 34224 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_372
timestamp 18001
transform 1 0 35328 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_380
timestamp 18001
transform 1 0 36064 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_393
timestamp 18001
transform 1 0 37260 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_399
timestamp 1636986456
transform 1 0 37812 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_411
timestamp 1636986456
transform 1 0 38916 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_423
timestamp 18001
transform 1 0 40020 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_429
timestamp 18001
transform 1 0 40572 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_438
timestamp 18001
transform 1 0 41400 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_446
timestamp 18001
transform 1 0 42136 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_449
timestamp 1636986456
transform 1 0 42412 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_461
timestamp 1636986456
transform 1 0 43516 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_473
timestamp 1636986456
transform 1 0 44620 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_485
timestamp 1636986456
transform 1 0 45724 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_497
timestamp 18001
transform 1 0 46828 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_503
timestamp 18001
transform 1 0 47380 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_505
timestamp 1636986456
transform 1 0 47564 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_517
timestamp 1636986456
transform 1 0 48668 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_529
timestamp 1636986456
transform 1 0 49772 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_541
timestamp 1636986456
transform 1 0 50876 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_553
timestamp 18001
transform 1 0 51980 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_559
timestamp 18001
transform 1 0 52532 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_561
timestamp 1636986456
transform 1 0 52716 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_573
timestamp 1636986456
transform 1 0 53820 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_585
timestamp 1636986456
transform 1 0 54924 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_597
timestamp 1636986456
transform 1 0 56028 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_609
timestamp 18001
transform 1 0 57132 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_615
timestamp 18001
transform 1 0 57684 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_617
timestamp 18001
transform 1 0 57868 0 -1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_3
timestamp 1636986456
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_15
timestamp 1636986456
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_27
timestamp 18001
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_29
timestamp 1636986456
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_41
timestamp 1636986456
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_53
timestamp 1636986456
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_65
timestamp 1636986456
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_77
timestamp 18001
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_83
timestamp 18001
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_85
timestamp 1636986456
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_97
timestamp 1636986456
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_109
timestamp 18001
transform 1 0 11132 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_117
timestamp 18001
transform 1 0 11868 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_148
timestamp 1636986456
transform 1 0 14720 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_160
timestamp 18001
transform 1 0 15824 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_194
timestamp 18001
transform 1 0 18952 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_197
timestamp 18001
transform 1 0 19228 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_203
timestamp 18001
transform 1 0 19780 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_211
timestamp 1636986456
transform 1 0 20516 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_223
timestamp 18001
transform 1 0 21620 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_241
timestamp 18001
transform 1 0 23276 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_249
timestamp 18001
transform 1 0 24012 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_253
timestamp 1636986456
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_265
timestamp 18001
transform 1 0 25484 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_275
timestamp 18001
transform 1 0 26404 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_286
timestamp 18001
transform 1 0 27416 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_301
timestamp 18001
transform 1 0 28796 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_307
timestamp 18001
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_309
timestamp 18001
transform 1 0 29532 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_322
timestamp 18001
transform 1 0 30728 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_329
timestamp 18001
transform 1 0 31372 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_335
timestamp 18001
transform 1 0 31924 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_352
timestamp 1636986456
transform 1 0 33488 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_365
timestamp 18001
transform 1 0 34684 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_369
timestamp 18001
transform 1 0 35052 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_379
timestamp 18001
transform 1 0 35972 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_393
timestamp 18001
transform 1 0 37260 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_399
timestamp 18001
transform 1 0 37812 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_405
timestamp 18001
transform 1 0 38364 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_421
timestamp 18001
transform 1 0 39836 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_445
timestamp 1636986456
transform 1 0 42044 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_457
timestamp 1636986456
transform 1 0 43148 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_469
timestamp 18001
transform 1 0 44252 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_475
timestamp 18001
transform 1 0 44804 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_477
timestamp 1636986456
transform 1 0 44988 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_489
timestamp 1636986456
transform 1 0 46092 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_501
timestamp 1636986456
transform 1 0 47196 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_513
timestamp 1636986456
transform 1 0 48300 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_525
timestamp 18001
transform 1 0 49404 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_531
timestamp 18001
transform 1 0 49956 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_533
timestamp 1636986456
transform 1 0 50140 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_545
timestamp 1636986456
transform 1 0 51244 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_557
timestamp 1636986456
transform 1 0 52348 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_569
timestamp 1636986456
transform 1 0 53452 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_581
timestamp 18001
transform 1 0 54556 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_587
timestamp 18001
transform 1 0 55108 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_589
timestamp 1636986456
transform 1 0 55292 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_601
timestamp 1636986456
transform 1 0 56396 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_613
timestamp 1636986456
transform 1 0 57500 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_3
timestamp 1636986456
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_15
timestamp 1636986456
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_27
timestamp 1636986456
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_39
timestamp 1636986456
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_51
timestamp 18001
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_55
timestamp 18001
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_57
timestamp 1636986456
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_69
timestamp 1636986456
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_81
timestamp 1636986456
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_93
timestamp 1636986456
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_105
timestamp 18001
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_111
timestamp 18001
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_113
timestamp 1636986456
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_125
timestamp 18001
transform 1 0 12604 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_148
timestamp 1636986456
transform 1 0 14720 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_160
timestamp 18001
transform 1 0 15824 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_176
timestamp 18001
transform 1 0 17296 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_216
timestamp 18001
transform 1 0 20976 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_225
timestamp 18001
transform 1 0 21804 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_247
timestamp 1636986456
transform 1 0 23828 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_289
timestamp 18001
transform 1 0 27692 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_293
timestamp 18001
transform 1 0 28060 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_311
timestamp 18001
transform 1 0 29716 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_319
timestamp 18001
transform 1 0 30452 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_330
timestamp 18001
transform 1 0 31464 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_337
timestamp 18001
transform 1 0 32108 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_348
timestamp 1636986456
transform 1 0 33120 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_360
timestamp 18001
transform 1 0 34224 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_386
timestamp 18001
transform 1 0 36616 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_404
timestamp 18001
transform 1 0 38272 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_410
timestamp 18001
transform 1 0 38824 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_414
timestamp 18001
transform 1 0 39192 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_418
timestamp 1636986456
transform 1 0 39560 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_430
timestamp 1636986456
transform 1 0 40664 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_442
timestamp 18001
transform 1 0 41768 0 -1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_449
timestamp 1636986456
transform 1 0 42412 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_461
timestamp 1636986456
transform 1 0 43516 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_473
timestamp 1636986456
transform 1 0 44620 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_485
timestamp 1636986456
transform 1 0 45724 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_497
timestamp 18001
transform 1 0 46828 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_503
timestamp 18001
transform 1 0 47380 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_505
timestamp 1636986456
transform 1 0 47564 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_517
timestamp 1636986456
transform 1 0 48668 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_529
timestamp 1636986456
transform 1 0 49772 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_541
timestamp 1636986456
transform 1 0 50876 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_553
timestamp 18001
transform 1 0 51980 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_559
timestamp 18001
transform 1 0 52532 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_561
timestamp 1636986456
transform 1 0 52716 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_573
timestamp 1636986456
transform 1 0 53820 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_585
timestamp 1636986456
transform 1 0 54924 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_597
timestamp 1636986456
transform 1 0 56028 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_609
timestamp 18001
transform 1 0 57132 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_615
timestamp 18001
transform 1 0 57684 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_617
timestamp 18001
transform 1 0 57868 0 -1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_3
timestamp 1636986456
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_15
timestamp 1636986456
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_27
timestamp 18001
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_29
timestamp 1636986456
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_41
timestamp 1636986456
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_53
timestamp 1636986456
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_65
timestamp 1636986456
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_77
timestamp 18001
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_83
timestamp 18001
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_85
timestamp 1636986456
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_97
timestamp 1636986456
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_109
timestamp 1636986456
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_128
timestamp 1636986456
transform 1 0 12880 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_145
timestamp 18001
transform 1 0 14444 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_161
timestamp 18001
transform 1 0 15916 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_177
timestamp 1636986456
transform 1 0 17388 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_193
timestamp 18001
transform 1 0 18860 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_197
timestamp 18001
transform 1 0 19228 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_211
timestamp 1636986456
transform 1 0 20516 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_223
timestamp 18001
transform 1 0 21620 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_253
timestamp 1636986456
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_265
timestamp 1636986456
transform 1 0 25484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_277
timestamp 18001
transform 1 0 26588 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_285
timestamp 18001
transform 1 0 27324 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_299
timestamp 18001
transform 1 0 28612 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_305
timestamp 18001
transform 1 0 29164 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_309
timestamp 18001
transform 1 0 29532 0 1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_323
timestamp 1636986456
transform 1 0 30820 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_335
timestamp 18001
transform 1 0 31924 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_344
timestamp 1636986456
transform 1 0 32752 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_356
timestamp 18001
transform 1 0 33856 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_365
timestamp 18001
transform 1 0 34684 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_374
timestamp 1636986456
transform 1 0 35512 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_386
timestamp 1636986456
transform 1 0 36616 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_398
timestamp 18001
transform 1 0 37720 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_411
timestamp 18001
transform 1 0 38916 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_419
timestamp 18001
transform 1 0 39652 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_429
timestamp 1636986456
transform 1 0 40572 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_441
timestamp 1636986456
transform 1 0 41676 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_453
timestamp 1636986456
transform 1 0 42780 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_465
timestamp 18001
transform 1 0 43884 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_473
timestamp 18001
transform 1 0 44620 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_477
timestamp 1636986456
transform 1 0 44988 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_489
timestamp 1636986456
transform 1 0 46092 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_501
timestamp 1636986456
transform 1 0 47196 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_513
timestamp 1636986456
transform 1 0 48300 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_525
timestamp 18001
transform 1 0 49404 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_531
timestamp 18001
transform 1 0 49956 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_533
timestamp 1636986456
transform 1 0 50140 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_545
timestamp 1636986456
transform 1 0 51244 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_557
timestamp 1636986456
transform 1 0 52348 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_569
timestamp 1636986456
transform 1 0 53452 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_581
timestamp 18001
transform 1 0 54556 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_587
timestamp 18001
transform 1 0 55108 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_589
timestamp 1636986456
transform 1 0 55292 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_601
timestamp 1636986456
transform 1 0 56396 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_613
timestamp 1636986456
transform 1 0 57500 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_3
timestamp 1636986456
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_15
timestamp 1636986456
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_27
timestamp 1636986456
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_39
timestamp 1636986456
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_51
timestamp 18001
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_55
timestamp 18001
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_57
timestamp 1636986456
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_69
timestamp 1636986456
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_81
timestamp 1636986456
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_93
timestamp 1636986456
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_105
timestamp 18001
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_111
timestamp 18001
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_113
timestamp 18001
transform 1 0 11500 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_119
timestamp 18001
transform 1 0 12052 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_153
timestamp 1636986456
transform 1 0 15180 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_165
timestamp 18001
transform 1 0 16284 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_169
timestamp 1636986456
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_181
timestamp 1636986456
transform 1 0 17756 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_193
timestamp 18001
transform 1 0 18860 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_219
timestamp 18001
transform 1 0 21252 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_223
timestamp 18001
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_225
timestamp 18001
transform 1 0 21804 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_229
timestamp 18001
transform 1 0 22172 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_238
timestamp 1636986456
transform 1 0 23000 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_250
timestamp 1636986456
transform 1 0 24104 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_262
timestamp 1636986456
transform 1 0 25208 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_274
timestamp 18001
transform 1 0 26312 0 -1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_288
timestamp 1636986456
transform 1 0 27600 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_300
timestamp 18001
transform 1 0 28704 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_308
timestamp 18001
transform 1 0 29440 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_317
timestamp 18001
transform 1 0 30268 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_329
timestamp 18001
transform 1 0 31372 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_335
timestamp 18001
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_337
timestamp 18001
transform 1 0 32108 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_356
timestamp 1636986456
transform 1 0 33856 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_376
timestamp 18001
transform 1 0 35696 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_388
timestamp 18001
transform 1 0 36800 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_393
timestamp 18001
transform 1 0 37260 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_425
timestamp 1636986456
transform 1 0 40204 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_437
timestamp 18001
transform 1 0 41308 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_445
timestamp 18001
transform 1 0 42044 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_449
timestamp 18001
transform 1 0 42412 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_470
timestamp 1636986456
transform 1 0 44344 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_482
timestamp 1636986456
transform 1 0 45448 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_494
timestamp 18001
transform 1 0 46552 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_502
timestamp 18001
transform 1 0 47288 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_505
timestamp 1636986456
transform 1 0 47564 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_517
timestamp 1636986456
transform 1 0 48668 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_529
timestamp 1636986456
transform 1 0 49772 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_541
timestamp 1636986456
transform 1 0 50876 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_553
timestamp 18001
transform 1 0 51980 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_559
timestamp 18001
transform 1 0 52532 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_561
timestamp 1636986456
transform 1 0 52716 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_573
timestamp 1636986456
transform 1 0 53820 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_585
timestamp 1636986456
transform 1 0 54924 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_597
timestamp 1636986456
transform 1 0 56028 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_609
timestamp 18001
transform 1 0 57132 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_615
timestamp 18001
transform 1 0 57684 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_617
timestamp 18001
transform 1 0 57868 0 -1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_3
timestamp 1636986456
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_15
timestamp 1636986456
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_27
timestamp 18001
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_29
timestamp 1636986456
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_41
timestamp 1636986456
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_53
timestamp 1636986456
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_65
timestamp 1636986456
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_77
timestamp 18001
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_83
timestamp 18001
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_85
timestamp 1636986456
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_97
timestamp 1636986456
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_109
timestamp 18001
transform 1 0 11132 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_117
timestamp 18001
transform 1 0 11868 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_152
timestamp 18001
transform 1 0 15088 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_193
timestamp 18001
transform 1 0 18860 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_236
timestamp 1636986456
transform 1 0 22816 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_248
timestamp 18001
transform 1 0 23920 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_253
timestamp 18001
transform 1 0 24380 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_286
timestamp 18001
transform 1 0 27416 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_293
timestamp 18001
transform 1 0 28060 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_307
timestamp 18001
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_323
timestamp 18001
transform 1 0 30820 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_334
timestamp 18001
transform 1 0 31832 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_342
timestamp 18001
transform 1 0 32568 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_361
timestamp 18001
transform 1 0 34316 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_365
timestamp 18001
transform 1 0 34684 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_382
timestamp 1636986456
transform 1 0 36248 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_394
timestamp 1636986456
transform 1 0 37352 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_406
timestamp 18001
transform 1 0 38456 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_415
timestamp 18001
transform 1 0 39284 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_419
timestamp 18001
transform 1 0 39652 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_436
timestamp 18001
transform 1 0 41216 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_440
timestamp 18001
transform 1 0 41584 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_461
timestamp 1636986456
transform 1 0 43516 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_473
timestamp 18001
transform 1 0 44620 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_477
timestamp 1636986456
transform 1 0 44988 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_489
timestamp 18001
transform 1 0 46092 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_498
timestamp 1636986456
transform 1 0 46920 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_510
timestamp 1636986456
transform 1 0 48024 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_522
timestamp 18001
transform 1 0 49128 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_530
timestamp 18001
transform 1 0 49864 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_533
timestamp 1636986456
transform 1 0 50140 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_545
timestamp 1636986456
transform 1 0 51244 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_557
timestamp 1636986456
transform 1 0 52348 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_569
timestamp 1636986456
transform 1 0 53452 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_581
timestamp 18001
transform 1 0 54556 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_587
timestamp 18001
transform 1 0 55108 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_589
timestamp 1636986456
transform 1 0 55292 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_601
timestamp 1636986456
transform 1 0 56396 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_613
timestamp 1636986456
transform 1 0 57500 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_3
timestamp 1636986456
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_15
timestamp 1636986456
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_27
timestamp 1636986456
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_39
timestamp 1636986456
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_51
timestamp 18001
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_55
timestamp 18001
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_57
timestamp 1636986456
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_69
timestamp 1636986456
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_81
timestamp 1636986456
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_93
timestamp 1636986456
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_105
timestamp 18001
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_111
timestamp 18001
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_113
timestamp 1636986456
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_125
timestamp 1636986456
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_137
timestamp 1636986456
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_149
timestamp 18001
transform 1 0 14812 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_164
timestamp 18001
transform 1 0 16192 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_169
timestamp 18001
transform 1 0 16652 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_191
timestamp 18001
transform 1 0 18676 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_199
timestamp 18001
transform 1 0 19412 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_204
timestamp 18001
transform 1 0 19872 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_218
timestamp 18001
transform 1 0 21160 0 -1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_225
timestamp 1636986456
transform 1 0 21804 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_237
timestamp 18001
transform 1 0 22908 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_245
timestamp 18001
transform 1 0 23644 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_281
timestamp 18001
transform 1 0 26956 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_293
timestamp 18001
transform 1 0 28060 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_297
timestamp 18001
transform 1 0 28428 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_305
timestamp 18001
transform 1 0 29164 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_311
timestamp 1636986456
transform 1 0 29716 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_323
timestamp 1636986456
transform 1 0 30820 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_335
timestamp 18001
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_343
timestamp 18001
transform 1 0 32660 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_353
timestamp 1636986456
transform 1 0 33580 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_365
timestamp 1636986456
transform 1 0 34684 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_377
timestamp 18001
transform 1 0 35788 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_383
timestamp 18001
transform 1 0 36340 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_391
timestamp 18001
transform 1 0 37076 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_398
timestamp 18001
transform 1 0 37720 0 -1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_418
timestamp 1636986456
transform 1 0 39560 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_430
timestamp 1636986456
transform 1 0 40664 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_442
timestamp 18001
transform 1 0 41768 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_458
timestamp 18001
transform 1 0 43240 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_470
timestamp 18001
transform 1 0 44344 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_478
timestamp 18001
transform 1 0 45080 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_499
timestamp 18001
transform 1 0 47012 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_503
timestamp 18001
transform 1 0 47380 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_505
timestamp 1636986456
transform 1 0 47564 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_517
timestamp 18001
transform 1 0 48668 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_538
timestamp 1636986456
transform 1 0 50600 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_550
timestamp 18001
transform 1 0 51704 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_558
timestamp 18001
transform 1 0 52440 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_561
timestamp 1636986456
transform 1 0 52716 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_573
timestamp 1636986456
transform 1 0 53820 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_585
timestamp 1636986456
transform 1 0 54924 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_597
timestamp 1636986456
transform 1 0 56028 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_609
timestamp 18001
transform 1 0 57132 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_615
timestamp 18001
transform 1 0 57684 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_617
timestamp 18001
transform 1 0 57868 0 -1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_3
timestamp 1636986456
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_15
timestamp 1636986456
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_27
timestamp 18001
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_29
timestamp 1636986456
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_41
timestamp 1636986456
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_53
timestamp 1636986456
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_65
timestamp 1636986456
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_77
timestamp 18001
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_83
timestamp 18001
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_85
timestamp 1636986456
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_97
timestamp 1636986456
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_109
timestamp 18001
transform 1 0 11132 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_117
timestamp 18001
transform 1 0 11868 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_138
timestamp 18001
transform 1 0 13800 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_141
timestamp 18001
transform 1 0 14076 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_147
timestamp 18001
transform 1 0 14628 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_211
timestamp 1636986456
transform 1 0 20516 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_223
timestamp 1636986456
transform 1 0 21620 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_235
timestamp 18001
transform 1 0 22724 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_243
timestamp 18001
transform 1 0 23460 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_253
timestamp 18001
transform 1 0 24380 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_266
timestamp 18001
transform 1 0 25576 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_270
timestamp 18001
transform 1 0 25944 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_281
timestamp 1636986456
transform 1 0 26956 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_293
timestamp 1636986456
transform 1 0 28060 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_305
timestamp 18001
transform 1 0 29164 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_316
timestamp 18001
transform 1 0 30176 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_320
timestamp 18001
transform 1 0 30544 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_327
timestamp 18001
transform 1 0 31188 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_341
timestamp 18001
transform 1 0 32476 0 1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_349
timestamp 1636986456
transform 1 0 33212 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_361
timestamp 18001
transform 1 0 34316 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_365
timestamp 1636986456
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_377
timestamp 18001
transform 1 0 35788 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_401
timestamp 18001
transform 1 0 37996 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_409
timestamp 18001
transform 1 0 38732 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_421
timestamp 18001
transform 1 0 39836 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_436
timestamp 18001
transform 1 0 41216 0 1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_448
timestamp 1636986456
transform 1 0 42320 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_460
timestamp 1636986456
transform 1 0 43424 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_472
timestamp 18001
transform 1 0 44528 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_477
timestamp 18001
transform 1 0 44988 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_555
timestamp 1636986456
transform 1 0 52164 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_567
timestamp 1636986456
transform 1 0 53268 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_579
timestamp 18001
transform 1 0 54372 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_587
timestamp 18001
transform 1 0 55108 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_611
timestamp 1636986456
transform 1 0 57316 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_623
timestamp 18001
transform 1 0 58420 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_3
timestamp 1636986456
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_15
timestamp 1636986456
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_27
timestamp 1636986456
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_39
timestamp 1636986456
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_51
timestamp 18001
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_55
timestamp 18001
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_57
timestamp 1636986456
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_69
timestamp 1636986456
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_81
timestamp 1636986456
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_93
timestamp 1636986456
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_105
timestamp 18001
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_111
timestamp 18001
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_113
timestamp 1636986456
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_125
timestamp 18001
transform 1 0 12604 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_148
timestamp 18001
transform 1 0 14720 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_162
timestamp 18001
transform 1 0 16008 0 -1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_169
timestamp 1636986456
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_181
timestamp 18001
transform 1 0 17756 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_209
timestamp 1636986456
transform 1 0 20332 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_221
timestamp 18001
transform 1 0 21436 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_245
timestamp 18001
transform 1 0 23644 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_281
timestamp 1636986456
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_293
timestamp 18001
transform 1 0 28060 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_327
timestamp 18001
transform 1 0 31188 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_335
timestamp 18001
transform 1 0 31924 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_340
timestamp 18001
transform 1 0 32384 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_366
timestamp 18001
transform 1 0 34776 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_374
timestamp 18001
transform 1 0 35512 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_383
timestamp 18001
transform 1 0 36340 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_391
timestamp 18001
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_393
timestamp 1636986456
transform 1 0 37260 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_405
timestamp 18001
transform 1 0 38364 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_476
timestamp 18001
transform 1 0 44896 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_484
timestamp 18001
transform 1 0 45632 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_503
timestamp 18001
transform 1 0 47380 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_515
timestamp 18001
transform 1 0 48484 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_571
timestamp 1636986456
transform 1 0 53636 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_583
timestamp 1636986456
transform 1 0 54740 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_595
timestamp 1636986456
transform 1 0 55844 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_607
timestamp 18001
transform 1 0 56948 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_615
timestamp 18001
transform 1 0 57684 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_617
timestamp 18001
transform 1 0 57868 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_8
timestamp 1636986456
transform 1 0 1840 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_20
timestamp 18001
transform 1 0 2944 0 1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_29
timestamp 1636986456
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_41
timestamp 1636986456
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_53
timestamp 1636986456
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_65
timestamp 1636986456
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_77
timestamp 18001
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_83
timestamp 18001
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_85
timestamp 1636986456
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_97
timestamp 1636986456
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_109
timestamp 18001
transform 1 0 11132 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_117
timestamp 18001
transform 1 0 11868 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_130
timestamp 18001
transform 1 0 13064 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_176
timestamp 1636986456
transform 1 0 17296 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_217
timestamp 18001
transform 1 0 21068 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_249
timestamp 18001
transform 1 0 24012 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_287
timestamp 18001
transform 1 0 27508 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_327
timestamp 1636986456
transform 1 0 31188 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_339
timestamp 18001
transform 1 0 32292 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_363
timestamp 18001
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_393
timestamp 1636986456
transform 1 0 37260 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_405
timestamp 1636986456
transform 1 0 38364 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_417
timestamp 18001
transform 1 0 39468 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_421
timestamp 18001
transform 1 0 39836 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_452
timestamp 18001
transform 1 0 42688 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_470
timestamp 18001
transform 1 0 44344 0 1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_477
timestamp 1636986456
transform 1 0 44988 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_489
timestamp 18001
transform 1 0 46092 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_508
timestamp 18001
transform 1 0 47840 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_533
timestamp 18001
transform 1 0 50140 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_541
timestamp 18001
transform 1 0 50876 0 1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_567
timestamp 1636986456
transform 1 0 53268 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_579
timestamp 18001
transform 1 0 54372 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_587
timestamp 18001
transform 1 0 55108 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_589
timestamp 1636986456
transform 1 0 55292 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_601
timestamp 1636986456
transform 1 0 56396 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_613
timestamp 1636986456
transform 1 0 57500 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_3
timestamp 1636986456
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_15
timestamp 1636986456
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_27
timestamp 1636986456
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_39
timestamp 1636986456
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_51
timestamp 18001
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_55
timestamp 18001
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_57
timestamp 1636986456
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_69
timestamp 1636986456
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_81
timestamp 1636986456
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_93
timestamp 1636986456
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_105
timestamp 18001
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_111
timestamp 18001
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_113
timestamp 1636986456
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_149
timestamp 18001
transform 1 0 14812 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_158
timestamp 18001
transform 1 0 15640 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_166
timestamp 18001
transform 1 0 16376 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_169
timestamp 1636986456
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_181
timestamp 18001
transform 1 0 17756 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_216
timestamp 18001
transform 1 0 20976 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_225
timestamp 18001
transform 1 0 21804 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_237
timestamp 18001
transform 1 0 22908 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_276
timestamp 18001
transform 1 0 26496 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_281
timestamp 1636986456
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_293
timestamp 1636986456
transform 1 0 28060 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_305
timestamp 18001
transform 1 0 29164 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_313
timestamp 18001
transform 1 0 29900 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_337
timestamp 18001
transform 1 0 32108 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_345
timestamp 18001
transform 1 0 32844 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_354
timestamp 18001
transform 1 0 33672 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_362
timestamp 18001
transform 1 0 34408 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_365
timestamp 1636986456
transform 1 0 34684 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_377
timestamp 18001
transform 1 0 35788 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_383
timestamp 18001
transform 1 0 36340 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_388
timestamp 18001
transform 1 0 36800 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_393
timestamp 18001
transform 1 0 37260 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_397
timestamp 18001
transform 1 0 37628 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_407
timestamp 18001
transform 1 0 38548 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_420
timestamp 1636986456
transform 1 0 39744 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_432
timestamp 1636986456
transform 1 0 40848 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_444
timestamp 18001
transform 1 0 41952 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_449
timestamp 18001
transform 1 0 42412 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_477
timestamp 1636986456
transform 1 0 44988 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_489
timestamp 18001
transform 1 0 46092 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_503
timestamp 18001
transform 1 0 47380 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_505
timestamp 18001
transform 1 0 47564 0 -1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_533
timestamp 1636986456
transform 1 0 50140 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_545
timestamp 18001
transform 1 0 51244 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_559
timestamp 18001
transform 1 0 52532 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_563
timestamp 18001
transform 1 0 52900 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_584
timestamp 18001
transform 1 0 54832 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_605
timestamp 18001
transform 1 0 56764 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_613
timestamp 18001
transform 1 0 57500 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_617
timestamp 18001
transform 1 0 57868 0 -1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_3
timestamp 1636986456
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_15
timestamp 1636986456
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_27
timestamp 18001
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_29
timestamp 1636986456
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_41
timestamp 1636986456
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_53
timestamp 1636986456
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_65
timestamp 1636986456
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_77
timestamp 18001
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_83
timestamp 18001
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_85
timestamp 1636986456
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_97
timestamp 1636986456
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_109
timestamp 1636986456
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_121
timestamp 18001
transform 1 0 12236 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_129
timestamp 18001
transform 1 0 12972 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_135
timestamp 18001
transform 1 0 13524 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_139
timestamp 18001
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_149
timestamp 1636986456
transform 1 0 14812 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_161
timestamp 1636986456
transform 1 0 15916 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_173
timestamp 1636986456
transform 1 0 17020 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_185
timestamp 18001
transform 1 0 18124 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_193
timestamp 18001
transform 1 0 18860 0 1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_209
timestamp 1636986456
transform 1 0 20332 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_221
timestamp 18001
transform 1 0 21436 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_233
timestamp 18001
transform 1 0 22540 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_259
timestamp 18001
transform 1 0 24932 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_263
timestamp 18001
transform 1 0 25300 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_270
timestamp 18001
transform 1 0 25944 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_278
timestamp 18001
transform 1 0 26680 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_284
timestamp 1636986456
transform 1 0 27232 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_296
timestamp 1636986456
transform 1 0 28336 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_309
timestamp 18001
transform 1 0 29532 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_329
timestamp 18001
transform 1 0 31372 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_339
timestamp 18001
transform 1 0 32292 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_349
timestamp 1636986456
transform 1 0 33212 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_361
timestamp 18001
transform 1 0 34316 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_365
timestamp 18001
transform 1 0 34684 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_419
timestamp 18001
transform 1 0 39652 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_421
timestamp 18001
transform 1 0 39836 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_433
timestamp 1636986456
transform 1 0 40940 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_445
timestamp 18001
transform 1 0 42044 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_456
timestamp 18001
transform 1 0 43056 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_460
timestamp 18001
transform 1 0 43424 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_468
timestamp 18001
transform 1 0 44160 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_477
timestamp 18001
transform 1 0 44988 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_483
timestamp 18001
transform 1 0 45540 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_504
timestamp 18001
transform 1 0 47472 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_508
timestamp 18001
transform 1 0 47840 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_513
timestamp 18001
transform 1 0 48300 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_522
timestamp 18001
transform 1 0 49128 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_530
timestamp 18001
transform 1 0 49864 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_541
timestamp 18001
transform 1 0 50876 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_545
timestamp 18001
transform 1 0 51244 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_576
timestamp 18001
transform 1 0 54096 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_587
timestamp 18001
transform 1 0 55108 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_610
timestamp 1636986456
transform 1 0 57224 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_622
timestamp 18001
transform 1 0 58328 0 1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_3
timestamp 1636986456
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_15
timestamp 1636986456
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_27
timestamp 1636986456
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_39
timestamp 1636986456
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_51
timestamp 18001
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_55
timestamp 18001
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_57
timestamp 1636986456
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_69
timestamp 1636986456
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_81
timestamp 1636986456
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_93
timestamp 1636986456
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_105
timestamp 18001
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_111
timestamp 18001
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_113
timestamp 1636986456
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_125
timestamp 1636986456
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_137
timestamp 1636986456
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_149
timestamp 1636986456
transform 1 0 14812 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_161
timestamp 18001
transform 1 0 15916 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_167
timestamp 18001
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_169
timestamp 1636986456
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_181
timestamp 1636986456
transform 1 0 17756 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_193
timestamp 18001
transform 1 0 18860 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_205
timestamp 1636986456
transform 1 0 19964 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_217
timestamp 18001
transform 1 0 21068 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_233
timestamp 18001
transform 1 0 22540 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_247
timestamp 18001
transform 1 0 23828 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_260
timestamp 18001
transform 1 0 25024 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_267
timestamp 18001
transform 1 0 25668 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_281
timestamp 18001
transform 1 0 26956 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_296
timestamp 18001
transform 1 0 28336 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_304
timestamp 18001
transform 1 0 29072 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_333
timestamp 18001
transform 1 0 31740 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_337
timestamp 18001
transform 1 0 32108 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_351
timestamp 18001
transform 1 0 33396 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_373
timestamp 18001
transform 1 0 35420 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_383
timestamp 18001
transform 1 0 36340 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_391
timestamp 18001
transform 1 0 37076 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_395
timestamp 18001
transform 1 0 37444 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_422
timestamp 18001
transform 1 0 39928 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_443
timestamp 18001
transform 1 0 41860 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_447
timestamp 18001
transform 1 0 42228 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_449
timestamp 18001
transform 1 0 42412 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_478
timestamp 1636986456
transform 1 0 45080 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_490
timestamp 18001
transform 1 0 46184 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_498
timestamp 18001
transform 1 0 46920 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_538
timestamp 1636986456
transform 1 0 50600 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_550
timestamp 18001
transform 1 0 51704 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_558
timestamp 18001
transform 1 0 52440 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_569
timestamp 18001
transform 1 0 53452 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_593
timestamp 18001
transform 1 0 55660 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_617
timestamp 18001
transform 1 0 57868 0 -1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_3
timestamp 1636986456
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_15
timestamp 1636986456
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_27
timestamp 18001
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_29
timestamp 1636986456
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_41
timestamp 1636986456
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_53
timestamp 1636986456
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_65
timestamp 1636986456
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_77
timestamp 18001
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_83
timestamp 18001
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_85
timestamp 1636986456
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_97
timestamp 1636986456
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_109
timestamp 1636986456
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_121
timestamp 1636986456
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_133
timestamp 18001
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_139
timestamp 18001
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_141
timestamp 1636986456
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_153
timestamp 1636986456
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_165
timestamp 18001
transform 1 0 16284 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_195
timestamp 18001
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_205
timestamp 18001
transform 1 0 19964 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_251
timestamp 18001
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_319
timestamp 18001
transform 1 0 30452 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_348
timestamp 1636986456
transform 1 0 33120 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_360
timestamp 18001
transform 1 0 34224 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_365
timestamp 18001
transform 1 0 34684 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_437
timestamp 18001
transform 1 0 41308 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_446
timestamp 18001
transform 1 0 42136 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_450
timestamp 18001
transform 1 0 42504 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_471
timestamp 18001
transform 1 0 44436 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_475
timestamp 18001
transform 1 0 44804 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_477
timestamp 18001
transform 1 0 44988 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_483
timestamp 18001
transform 1 0 45540 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_488
timestamp 18001
transform 1 0 46000 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_505
timestamp 18001
transform 1 0 47564 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_533
timestamp 1636986456
transform 1 0 50140 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_545
timestamp 1636986456
transform 1 0 51244 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_557
timestamp 1636986456
transform 1 0 52348 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_569
timestamp 18001
transform 1 0 53452 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_614
timestamp 18001
transform 1 0 57592 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_622
timestamp 18001
transform 1 0 58328 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_3
timestamp 1636986456
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_15
timestamp 1636986456
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_27
timestamp 1636986456
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_39
timestamp 1636986456
transform 1 0 4692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_51
timestamp 18001
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_55
timestamp 18001
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_57
timestamp 1636986456
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_69
timestamp 1636986456
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_81
timestamp 1636986456
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_93
timestamp 1636986456
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_105
timestamp 18001
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_111
timestamp 18001
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_113
timestamp 1636986456
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_125
timestamp 1636986456
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_137
timestamp 1636986456
transform 1 0 13708 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_149
timestamp 1636986456
transform 1 0 14812 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_161
timestamp 18001
transform 1 0 15916 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_167
timestamp 18001
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_169
timestamp 18001
transform 1 0 16652 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_207
timestamp 1636986456
transform 1 0 20148 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_219
timestamp 18001
transform 1 0 21252 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_223
timestamp 18001
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_225
timestamp 1636986456
transform 1 0 21804 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_243
timestamp 18001
transform 1 0 23460 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_277
timestamp 18001
transform 1 0 26588 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_283
timestamp 18001
transform 1 0 27140 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_291
timestamp 1636986456
transform 1 0 27876 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_303
timestamp 18001
transform 1 0 28980 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_317
timestamp 18001
transform 1 0 30268 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_343
timestamp 18001
transform 1 0 32660 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_351
timestamp 18001
transform 1 0 33396 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_383
timestamp 18001
transform 1 0 36340 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_389
timestamp 18001
transform 1 0 36892 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_399
timestamp 18001
transform 1 0 37812 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_407
timestamp 18001
transform 1 0 38548 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_440
timestamp 18001
transform 1 0 41584 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_496
timestamp 18001
transform 1 0 46736 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_502
timestamp 18001
transform 1 0 47288 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_518
timestamp 18001
transform 1 0 48760 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_527
timestamp 18001
transform 1 0 49588 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_545
timestamp 18001
transform 1 0 51244 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_556
timestamp 18001
transform 1 0 52256 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_568
timestamp 18001
transform 1 0 53360 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_617
timestamp 18001
transform 1 0 57868 0 -1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_3
timestamp 1636986456
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_15
timestamp 1636986456
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_27
timestamp 18001
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_29
timestamp 1636986456
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_41
timestamp 1636986456
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_53
timestamp 1636986456
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_65
timestamp 1636986456
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_77
timestamp 18001
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_83
timestamp 18001
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_85
timestamp 1636986456
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_97
timestamp 1636986456
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_109
timestamp 1636986456
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_121
timestamp 1636986456
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_133
timestamp 18001
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_139
timestamp 18001
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_141
timestamp 1636986456
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_153
timestamp 1636986456
transform 1 0 15180 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_165
timestamp 18001
transform 1 0 16284 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_180
timestamp 1636986456
transform 1 0 17664 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_192
timestamp 18001
transform 1 0 18768 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_197
timestamp 1636986456
transform 1 0 19228 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_209
timestamp 1636986456
transform 1 0 20332 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_221
timestamp 1636986456
transform 1 0 21436 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_233
timestamp 1636986456
transform 1 0 22540 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_245
timestamp 18001
transform 1 0 23644 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_251
timestamp 18001
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_253
timestamp 18001
transform 1 0 24380 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_258
timestamp 18001
transform 1 0 24840 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_266
timestamp 18001
transform 1 0 25576 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_276
timestamp 1636986456
transform 1 0 26496 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_288
timestamp 1636986456
transform 1 0 27600 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_300
timestamp 18001
transform 1 0 28704 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_309
timestamp 18001
transform 1 0 29532 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_321
timestamp 18001
transform 1 0 30636 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_342
timestamp 1636986456
transform 1 0 32568 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_354
timestamp 18001
transform 1 0 33672 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_362
timestamp 18001
transform 1 0 34408 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_372
timestamp 18001
transform 1 0 35328 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_378
timestamp 18001
transform 1 0 35880 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_393
timestamp 1636986456
transform 1 0 37260 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_409
timestamp 18001
transform 1 0 38732 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_419
timestamp 18001
transform 1 0 39652 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_429
timestamp 18001
transform 1 0 40572 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_466
timestamp 18001
transform 1 0 43976 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_474
timestamp 18001
transform 1 0 44712 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_477
timestamp 1636986456
transform 1 0 44988 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_489
timestamp 18001
transform 1 0 46092 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_523
timestamp 18001
transform 1 0 49220 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_531
timestamp 18001
transform 1 0 49956 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_533
timestamp 18001
transform 1 0 50140 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_537
timestamp 18001
transform 1 0 50508 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_587
timestamp 18001
transform 1 0 55108 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_589
timestamp 18001
transform 1 0 55292 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_622
timestamp 18001
transform 1 0 58328 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_3
timestamp 1636986456
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_15
timestamp 1636986456
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_27
timestamp 1636986456
transform 1 0 3588 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_39
timestamp 1636986456
transform 1 0 4692 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_51
timestamp 18001
transform 1 0 5796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_55
timestamp 18001
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_57
timestamp 1636986456
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_69
timestamp 1636986456
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_81
timestamp 1636986456
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_93
timestamp 1636986456
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_105
timestamp 18001
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_111
timestamp 18001
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_113
timestamp 1636986456
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_125
timestamp 1636986456
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_137
timestamp 1636986456
transform 1 0 13708 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_149
timestamp 1636986456
transform 1 0 14812 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_161
timestamp 18001
transform 1 0 15916 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_167
timestamp 18001
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_182
timestamp 18001
transform 1 0 17848 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_212
timestamp 1636986456
transform 1 0 20608 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_225
timestamp 18001
transform 1 0 21804 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_233
timestamp 18001
transform 1 0 22540 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_239
timestamp 18001
transform 1 0 23092 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_247
timestamp 18001
transform 1 0 23828 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_255
timestamp 18001
transform 1 0 24564 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_283
timestamp 18001
transform 1 0 27140 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_291
timestamp 18001
transform 1 0 27876 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_307
timestamp 18001
transform 1 0 29348 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_315
timestamp 18001
transform 1 0 30084 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_335
timestamp 18001
transform 1 0 31924 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_343
timestamp 1636986456
transform 1 0 32660 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_355
timestamp 1636986456
transform 1 0 33764 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_367
timestamp 18001
transform 1 0 34868 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_371
timestamp 18001
transform 1 0 35236 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_393
timestamp 18001
transform 1 0 37260 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_397
timestamp 18001
transform 1 0 37628 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_443
timestamp 18001
transform 1 0 41860 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_447
timestamp 18001
transform 1 0 42228 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_449
timestamp 18001
transform 1 0 42412 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_453
timestamp 18001
transform 1 0 42780 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_456
timestamp 1636986456
transform 1 0 43056 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_468
timestamp 1636986456
transform 1 0 44160 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_480
timestamp 18001
transform 1 0 45264 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_491
timestamp 1636986456
transform 1 0 46276 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_503
timestamp 18001
transform 1 0 47380 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_505
timestamp 1636986456
transform 1 0 47564 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_517
timestamp 1636986456
transform 1 0 48668 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_529
timestamp 18001
transform 1 0 49772 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_538
timestamp 1636986456
transform 1 0 50600 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_550
timestamp 18001
transform 1 0 51704 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_558
timestamp 18001
transform 1 0 52440 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_570
timestamp 18001
transform 1 0 53544 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_580
timestamp 1636986456
transform 1 0 54464 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_592
timestamp 18001
transform 1 0 55568 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_596
timestamp 18001
transform 1 0 55936 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_599
timestamp 18001
transform 1 0 56212 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_613
timestamp 18001
transform 1 0 57500 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_3
timestamp 1636986456
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_15
timestamp 1636986456
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_27
timestamp 18001
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_29
timestamp 1636986456
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_41
timestamp 1636986456
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_53
timestamp 1636986456
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_65
timestamp 1636986456
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_77
timestamp 18001
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_83
timestamp 18001
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_85
timestamp 1636986456
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_97
timestamp 1636986456
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_109
timestamp 1636986456
transform 1 0 11132 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_121
timestamp 1636986456
transform 1 0 12236 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_133
timestamp 18001
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_139
timestamp 18001
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_141
timestamp 1636986456
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_153
timestamp 18001
transform 1 0 15180 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_173
timestamp 18001
transform 1 0 17020 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_197
timestamp 18001
transform 1 0 19228 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_209
timestamp 18001
transform 1 0 20332 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_250
timestamp 18001
transform 1 0 24104 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_253
timestamp 18001
transform 1 0 24380 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_261
timestamp 18001
transform 1 0 25116 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_280
timestamp 18001
transform 1 0 26864 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_309
timestamp 18001
transform 1 0 29532 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_313
timestamp 18001
transform 1 0 29900 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_341
timestamp 1636986456
transform 1 0 32476 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_353
timestamp 18001
transform 1 0 33580 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_365
timestamp 18001
transform 1 0 34684 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_392
timestamp 18001
transform 1 0 37168 0 1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_429
timestamp 1636986456
transform 1 0 40572 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_441
timestamp 1636986456
transform 1 0 41676 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_453
timestamp 1636986456
transform 1 0 42780 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_465
timestamp 18001
transform 1 0 43884 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_473
timestamp 18001
transform 1 0 44620 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_497
timestamp 18001
transform 1 0 46828 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_527
timestamp 18001
transform 1 0 49588 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_531
timestamp 18001
transform 1 0 49956 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_540
timestamp 18001
transform 1 0 50784 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_548
timestamp 18001
transform 1 0 51520 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_555
timestamp 18001
transform 1 0 52164 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_563
timestamp 18001
transform 1 0 52900 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_568
timestamp 1636986456
transform 1 0 53360 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_580
timestamp 18001
transform 1 0 54464 0 1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_589
timestamp 1636986456
transform 1 0 55292 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_601
timestamp 18001
transform 1 0 56396 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_605
timestamp 18001
transform 1 0 56764 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_622
timestamp 18001
transform 1 0 58328 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_3
timestamp 1636986456
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_15
timestamp 1636986456
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_27
timestamp 1636986456
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_39
timestamp 1636986456
transform 1 0 4692 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_51
timestamp 18001
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_55
timestamp 18001
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_57
timestamp 1636986456
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_69
timestamp 1636986456
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_81
timestamp 1636986456
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_93
timestamp 1636986456
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_105
timestamp 18001
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_111
timestamp 18001
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_113
timestamp 1636986456
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_125
timestamp 1636986456
transform 1 0 12604 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_137
timestamp 1636986456
transform 1 0 13708 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_149
timestamp 18001
transform 1 0 14812 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_167
timestamp 18001
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_169
timestamp 1636986456
transform 1 0 16652 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_181
timestamp 18001
transform 1 0 17756 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_189
timestamp 18001
transform 1 0 18492 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_208
timestamp 1636986456
transform 1 0 20240 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_220
timestamp 18001
transform 1 0 21344 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_234
timestamp 18001
transform 1 0 22632 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_245
timestamp 18001
transform 1 0 23644 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_253
timestamp 18001
transform 1 0 24380 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_279
timestamp 18001
transform 1 0 26772 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_283
timestamp 18001
transform 1 0 27140 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_291
timestamp 18001
transform 1 0 27876 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_304
timestamp 1636986456
transform 1 0 29072 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_316
timestamp 18001
transform 1 0 30176 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_331
timestamp 18001
transform 1 0 31556 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_335
timestamp 18001
transform 1 0 31924 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_337
timestamp 1636986456
transform 1 0 32108 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_349
timestamp 18001
transform 1 0 33212 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_357
timestamp 18001
transform 1 0 33948 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_380
timestamp 1636986456
transform 1 0 36064 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_393
timestamp 18001
transform 1 0 37260 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_399
timestamp 18001
transform 1 0 37812 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_407
timestamp 18001
transform 1 0 38548 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_418
timestamp 18001
transform 1 0 39560 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_426
timestamp 18001
transform 1 0 40296 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_444
timestamp 18001
transform 1 0 41952 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_449
timestamp 1636986456
transform 1 0 42412 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_461
timestamp 18001
transform 1 0 43516 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_524
timestamp 18001
transform 1 0 49312 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_556
timestamp 18001
transform 1 0 52256 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_567
timestamp 18001
transform 1 0 53268 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_588
timestamp 1636986456
transform 1 0 55200 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_600
timestamp 18001
transform 1 0 56304 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_613
timestamp 18001
transform 1 0 57500 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_7
timestamp 1636986456
transform 1 0 1748 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_19
timestamp 18001
transform 1 0 2852 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_27
timestamp 18001
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_29
timestamp 1636986456
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_41
timestamp 1636986456
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_53
timestamp 1636986456
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_65
timestamp 1636986456
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_77
timestamp 18001
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_83
timestamp 18001
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_85
timestamp 1636986456
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_97
timestamp 1636986456
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_109
timestamp 1636986456
transform 1 0 11132 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_121
timestamp 1636986456
transform 1 0 12236 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_133
timestamp 18001
transform 1 0 13340 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_139
timestamp 18001
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_141
timestamp 1636986456
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_153
timestamp 1636986456
transform 1 0 15180 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_165
timestamp 1636986456
transform 1 0 16284 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_177
timestamp 1636986456
transform 1 0 17388 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_189
timestamp 18001
transform 1 0 18492 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_195
timestamp 18001
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_197
timestamp 1636986456
transform 1 0 19228 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_209
timestamp 1636986456
transform 1 0 20332 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_221
timestamp 1636986456
transform 1 0 21436 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_233
timestamp 1636986456
transform 1 0 22540 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_245
timestamp 18001
transform 1 0 23644 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_251
timestamp 18001
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_253
timestamp 18001
transform 1 0 24380 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_257
timestamp 18001
transform 1 0 24748 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_287
timestamp 1636986456
transform 1 0 27508 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_299
timestamp 18001
transform 1 0 28612 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_307
timestamp 18001
transform 1 0 29348 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_309
timestamp 18001
transform 1 0 29532 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_325
timestamp 18001
transform 1 0 31004 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_338
timestamp 1636986456
transform 1 0 32200 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_350
timestamp 18001
transform 1 0 33304 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_354
timestamp 18001
transform 1 0 33672 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_390
timestamp 18001
transform 1 0 36984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_419
timestamp 18001
transform 1 0 39652 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_421
timestamp 1636986456
transform 1 0 39836 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_433
timestamp 18001
transform 1 0 40940 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_444
timestamp 1636986456
transform 1 0 41952 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_530
timestamp 18001
transform 1 0 49864 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_533
timestamp 18001
transform 1 0 50140 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_575
timestamp 18001
transform 1 0 54004 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_579
timestamp 18001
transform 1 0 54372 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_609
timestamp 18001
transform 1 0 57132 0 1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_3
timestamp 1636986456
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_15
timestamp 1636986456
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_27
timestamp 1636986456
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_39
timestamp 1636986456
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_51
timestamp 18001
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_55
timestamp 18001
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_57
timestamp 1636986456
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_69
timestamp 1636986456
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_81
timestamp 1636986456
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_93
timestamp 1636986456
transform 1 0 9660 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_105
timestamp 18001
transform 1 0 10764 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_111
timestamp 18001
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_113
timestamp 1636986456
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_125
timestamp 1636986456
transform 1 0 12604 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_137
timestamp 1636986456
transform 1 0 13708 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_149
timestamp 1636986456
transform 1 0 14812 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_161
timestamp 18001
transform 1 0 15916 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_167
timestamp 18001
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_169
timestamp 1636986456
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_181
timestamp 18001
transform 1 0 17756 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_217
timestamp 18001
transform 1 0 21068 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_223
timestamp 18001
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_262
timestamp 18001
transform 1 0 25208 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_276
timestamp 18001
transform 1 0 26496 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_281
timestamp 1636986456
transform 1 0 26956 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_293
timestamp 18001
transform 1 0 28060 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_309
timestamp 18001
transform 1 0 29532 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_330
timestamp 18001
transform 1 0 31464 0 -1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_337
timestamp 1636986456
transform 1 0 32108 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_349
timestamp 18001
transform 1 0 33212 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_390
timestamp 18001
transform 1 0 36984 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_393
timestamp 1636986456
transform 1 0 37260 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_405
timestamp 18001
transform 1 0 38364 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_420
timestamp 18001
transform 1 0 39744 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_463
timestamp 18001
transform 1 0 43700 0 -1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_485
timestamp 1636986456
transform 1 0 45724 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_497
timestamp 18001
transform 1 0 46828 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_503
timestamp 18001
transform 1 0 47380 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_535
timestamp 1636986456
transform 1 0 50324 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_547
timestamp 1636986456
transform 1 0 51428 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_559
timestamp 18001
transform 1 0 52532 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_561
timestamp 18001
transform 1 0 52716 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_567
timestamp 18001
transform 1 0 53268 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_575
timestamp 1636986456
transform 1 0 54004 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_593
timestamp 18001
transform 1 0 55660 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_606
timestamp 18001
transform 1 0 56856 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_614
timestamp 18001
transform 1 0 57592 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_617
timestamp 18001
transform 1 0 57868 0 -1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_3
timestamp 1636986456
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_15
timestamp 1636986456
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_27
timestamp 18001
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_29
timestamp 1636986456
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_41
timestamp 1636986456
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_53
timestamp 1636986456
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_65
timestamp 1636986456
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_77
timestamp 18001
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_83
timestamp 18001
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_85
timestamp 1636986456
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_97
timestamp 1636986456
transform 1 0 10028 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_109
timestamp 1636986456
transform 1 0 11132 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_121
timestamp 1636986456
transform 1 0 12236 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_133
timestamp 18001
transform 1 0 13340 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_139
timestamp 18001
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_141
timestamp 1636986456
transform 1 0 14076 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_153
timestamp 1636986456
transform 1 0 15180 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_165
timestamp 1636986456
transform 1 0 16284 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_177
timestamp 1636986456
transform 1 0 17388 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_217
timestamp 18001
transform 1 0 21068 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_268
timestamp 18001
transform 1 0 25760 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_283
timestamp 18001
transform 1 0 27140 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_287
timestamp 18001
transform 1 0 27508 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_316
timestamp 18001
transform 1 0 30176 0 1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_348
timestamp 1636986456
transform 1 0 33120 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_360
timestamp 18001
transform 1 0 34224 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_365
timestamp 18001
transform 1 0 34684 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_368
timestamp 18001
transform 1 0 34960 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_376
timestamp 18001
transform 1 0 35696 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_389
timestamp 18001
transform 1 0 36892 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_397
timestamp 18001
transform 1 0 37628 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_429
timestamp 18001
transform 1 0 40572 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_458
timestamp 18001
transform 1 0 43240 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_464
timestamp 18001
transform 1 0 43792 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_475
timestamp 18001
transform 1 0 44804 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_488
timestamp 18001
transform 1 0 46000 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_492
timestamp 18001
transform 1 0 46368 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_513
timestamp 18001
transform 1 0 48300 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_547
timestamp 18001
transform 1 0 51428 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_559
timestamp 1636986456
transform 1 0 52532 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_571
timestamp 1636986456
transform 1 0 53636 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_583
timestamp 18001
transform 1 0 54740 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_589
timestamp 18001
transform 1 0 55292 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_620
timestamp 18001
transform 1 0 58144 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_624
timestamp 18001
transform 1 0 58512 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_3
timestamp 1636986456
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_15
timestamp 1636986456
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_27
timestamp 1636986456
transform 1 0 3588 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_39
timestamp 1636986456
transform 1 0 4692 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_51
timestamp 18001
transform 1 0 5796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_55
timestamp 18001
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_57
timestamp 1636986456
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_69
timestamp 1636986456
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_81
timestamp 1636986456
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_93
timestamp 1636986456
transform 1 0 9660 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_105
timestamp 18001
transform 1 0 10764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_111
timestamp 18001
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_113
timestamp 1636986456
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_125
timestamp 1636986456
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_137
timestamp 1636986456
transform 1 0 13708 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_149
timestamp 1636986456
transform 1 0 14812 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_161
timestamp 18001
transform 1 0 15916 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_167
timestamp 18001
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_169
timestamp 1636986456
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_181
timestamp 1636986456
transform 1 0 17756 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_216
timestamp 18001
transform 1 0 20976 0 -1 21760
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_225
timestamp 1636986456
transform 1 0 21804 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_237
timestamp 18001
transform 1 0 22908 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_241
timestamp 18001
transform 1 0 23276 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_260
timestamp 18001
transform 1 0 25024 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_327
timestamp 18001
transform 1 0 31188 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_348
timestamp 18001
transform 1 0 33120 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_356
timestamp 18001
transform 1 0 33856 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_387
timestamp 18001
transform 1 0 36708 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_391
timestamp 18001
transform 1 0 37076 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_393
timestamp 1636986456
transform 1 0 37260 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_405
timestamp 1636986456
transform 1 0 38364 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_417
timestamp 1636986456
transform 1 0 39468 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_429
timestamp 18001
transform 1 0 40572 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_437
timestamp 18001
transform 1 0 41308 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_449
timestamp 1636986456
transform 1 0 42412 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_461
timestamp 18001
transform 1 0 43516 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_497
timestamp 18001
transform 1 0 46828 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_501
timestamp 18001
transform 1 0 47196 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_533
timestamp 18001
transform 1 0 50140 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_595
timestamp 18001
transform 1 0 55844 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_602
timestamp 18001
transform 1 0 56488 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_614
timestamp 18001
transform 1 0 57592 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_3
timestamp 1636986456
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_15
timestamp 1636986456
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_27
timestamp 18001
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_29
timestamp 1636986456
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_41
timestamp 1636986456
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_53
timestamp 1636986456
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_65
timestamp 1636986456
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_77
timestamp 18001
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_83
timestamp 18001
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_85
timestamp 1636986456
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_97
timestamp 1636986456
transform 1 0 10028 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_109
timestamp 1636986456
transform 1 0 11132 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_121
timestamp 1636986456
transform 1 0 12236 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_133
timestamp 18001
transform 1 0 13340 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_139
timestamp 18001
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_141
timestamp 1636986456
transform 1 0 14076 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_153
timestamp 1636986456
transform 1 0 15180 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_165
timestamp 1636986456
transform 1 0 16284 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_177
timestamp 1636986456
transform 1 0 17388 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_189
timestamp 18001
transform 1 0 18492 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_197
timestamp 18001
transform 1 0 19228 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_201
timestamp 18001
transform 1 0 19596 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_210
timestamp 1636986456
transform 1 0 20424 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_222
timestamp 1636986456
transform 1 0 21528 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_234
timestamp 18001
transform 1 0 22632 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_242
timestamp 18001
transform 1 0 23368 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_248
timestamp 18001
transform 1 0 23920 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_253
timestamp 1636986456
transform 1 0 24380 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_265
timestamp 18001
transform 1 0 25484 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_294
timestamp 1636986456
transform 1 0 28152 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_306
timestamp 18001
transform 1 0 29256 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_313
timestamp 1636986456
transform 1 0 29900 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_325
timestamp 18001
transform 1 0 31004 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_354
timestamp 18001
transform 1 0 33672 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_362
timestamp 18001
transform 1 0 34408 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_365
timestamp 18001
transform 1 0 34684 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_402
timestamp 1636986456
transform 1 0 38088 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_414
timestamp 18001
transform 1 0 39192 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_421
timestamp 18001
transform 1 0 39836 0 1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_450
timestamp 1636986456
transform 1 0 42504 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_462
timestamp 1636986456
transform 1 0 43608 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_474
timestamp 18001
transform 1 0 44712 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_482
timestamp 1636986456
transform 1 0 45448 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_494
timestamp 18001
transform 1 0 46552 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_502
timestamp 18001
transform 1 0 47288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_530
timestamp 18001
transform 1 0 49864 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_533
timestamp 18001
transform 1 0 50140 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_542
timestamp 1636986456
transform 1 0 50968 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_566
timestamp 18001
transform 1 0 53176 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_576
timestamp 1636986456
transform 1 0 54096 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_595
timestamp 18001
transform 1 0 55844 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_603
timestamp 18001
transform 1 0 56580 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_622
timestamp 18001
transform 1 0 58328 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_3
timestamp 1636986456
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_15
timestamp 1636986456
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_27
timestamp 1636986456
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_39
timestamp 1636986456
transform 1 0 4692 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_51
timestamp 18001
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_55
timestamp 18001
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_57
timestamp 1636986456
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_69
timestamp 1636986456
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_81
timestamp 1636986456
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_93
timestamp 1636986456
transform 1 0 9660 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_105
timestamp 18001
transform 1 0 10764 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_111
timestamp 18001
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_113
timestamp 1636986456
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_125
timestamp 1636986456
transform 1 0 12604 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_137
timestamp 1636986456
transform 1 0 13708 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_149
timestamp 1636986456
transform 1 0 14812 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_161
timestamp 18001
transform 1 0 15916 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_167
timestamp 18001
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_169
timestamp 1636986456
transform 1 0 16652 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_181
timestamp 18001
transform 1 0 17756 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_200
timestamp 18001
transform 1 0 19504 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_211
timestamp 1636986456
transform 1 0 20516 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_223
timestamp 18001
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_245
timestamp 1636986456
transform 1 0 23644 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_257
timestamp 18001
transform 1 0 24748 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_265
timestamp 18001
transform 1 0 25484 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_275
timestamp 18001
transform 1 0 26404 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_279
timestamp 18001
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_281
timestamp 1636986456
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_302
timestamp 1636986456
transform 1 0 28888 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_314
timestamp 1636986456
transform 1 0 29992 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_326
timestamp 18001
transform 1 0 31096 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_334
timestamp 18001
transform 1 0 31832 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_348
timestamp 1636986456
transform 1 0 33120 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_360
timestamp 18001
transform 1 0 34224 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_366
timestamp 18001
transform 1 0 34776 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_389
timestamp 18001
transform 1 0 36892 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_393
timestamp 18001
transform 1 0 37260 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_397
timestamp 18001
transform 1 0 37628 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_406
timestamp 18001
transform 1 0 38456 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_412
timestamp 18001
transform 1 0 39008 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_423
timestamp 18001
transform 1 0 40020 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_431
timestamp 18001
transform 1 0 40756 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_444
timestamp 18001
transform 1 0 41952 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_458
timestamp 18001
transform 1 0 43240 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_466
timestamp 18001
transform 1 0 43976 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_487
timestamp 1636986456
transform 1 0 45908 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_499
timestamp 18001
transform 1 0 47012 0 -1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_528
timestamp 1636986456
transform 1 0 49680 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_540
timestamp 1636986456
transform 1 0 50784 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_552
timestamp 18001
transform 1 0 51888 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_578
timestamp 18001
transform 1 0 54280 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_599
timestamp 1636986456
transform 1 0 56212 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_611
timestamp 18001
transform 1 0 57316 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_615
timestamp 18001
transform 1 0 57684 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_617
timestamp 18001
transform 1 0 57868 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_3
timestamp 1636986456
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_15
timestamp 1636986456
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_27
timestamp 18001
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_29
timestamp 1636986456
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_41
timestamp 1636986456
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_53
timestamp 1636986456
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_65
timestamp 1636986456
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_77
timestamp 18001
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_83
timestamp 18001
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_85
timestamp 1636986456
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_97
timestamp 1636986456
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_109
timestamp 1636986456
transform 1 0 11132 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_121
timestamp 1636986456
transform 1 0 12236 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_133
timestamp 18001
transform 1 0 13340 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_139
timestamp 18001
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_141
timestamp 1636986456
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_153
timestamp 1636986456
transform 1 0 15180 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_165
timestamp 1636986456
transform 1 0 16284 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_177
timestamp 18001
transform 1 0 17388 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_217
timestamp 18001
transform 1 0 21068 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_248
timestamp 18001
transform 1 0 23920 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_253
timestamp 1636986456
transform 1 0 24380 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_265
timestamp 18001
transform 1 0 25484 0 1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_275
timestamp 1636986456
transform 1 0 26404 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_309
timestamp 18001
transform 1 0 29532 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_317
timestamp 18001
transform 1 0 30268 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_347
timestamp 1636986456
transform 1 0 33028 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_359
timestamp 18001
transform 1 0 34132 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_363
timestamp 18001
transform 1 0 34500 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_365
timestamp 18001
transform 1 0 34684 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_388
timestamp 1636986456
transform 1 0 36800 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_400
timestamp 18001
transform 1 0 37904 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_430
timestamp 18001
transform 1 0 40664 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_447
timestamp 18001
transform 1 0 42228 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_467
timestamp 18001
transform 1 0 44068 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_493
timestamp 18001
transform 1 0 46460 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_517
timestamp 18001
transform 1 0 48668 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_527
timestamp 18001
transform 1 0 49588 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_531
timestamp 18001
transform 1 0 49956 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_533
timestamp 18001
transform 1 0 50140 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_542
timestamp 18001
transform 1 0 50968 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_550
timestamp 18001
transform 1 0 51704 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_572
timestamp 18001
transform 1 0 53728 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_589
timestamp 18001
transform 1 0 55292 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_613
timestamp 1636986456
transform 1 0 57500 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_3
timestamp 1636986456
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_15
timestamp 1636986456
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_27
timestamp 1636986456
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_39
timestamp 1636986456
transform 1 0 4692 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_51
timestamp 18001
transform 1 0 5796 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_55
timestamp 18001
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_57
timestamp 1636986456
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_69
timestamp 1636986456
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_81
timestamp 1636986456
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_93
timestamp 1636986456
transform 1 0 9660 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_105
timestamp 18001
transform 1 0 10764 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_111
timestamp 18001
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_113
timestamp 1636986456
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_125
timestamp 1636986456
transform 1 0 12604 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_137
timestamp 1636986456
transform 1 0 13708 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_149
timestamp 1636986456
transform 1 0 14812 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_161
timestamp 18001
transform 1 0 15916 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_167
timestamp 18001
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_169
timestamp 1636986456
transform 1 0 16652 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_181
timestamp 18001
transform 1 0 17756 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_185
timestamp 18001
transform 1 0 18124 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_213
timestamp 18001
transform 1 0 20700 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_225
timestamp 18001
transform 1 0 21804 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_240
timestamp 18001
transform 1 0 23184 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_250
timestamp 18001
transform 1 0 24104 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_279
timestamp 18001
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_285
timestamp 18001
transform 1 0 27324 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_305
timestamp 1636986456
transform 1 0 29164 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_317
timestamp 1636986456
transform 1 0 30268 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_329
timestamp 18001
transform 1 0 31372 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_335
timestamp 18001
transform 1 0 31924 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_344
timestamp 18001
transform 1 0 32752 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_350
timestamp 18001
transform 1 0 33304 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_356
timestamp 18001
transform 1 0 33856 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_367
timestamp 18001
transform 1 0 34868 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_393
timestamp 18001
transform 1 0 37260 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_401
timestamp 18001
transform 1 0 37996 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_431
timestamp 1636986456
transform 1 0 40756 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_443
timestamp 18001
transform 1 0 41860 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_447
timestamp 18001
transform 1 0 42228 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_469
timestamp 18001
transform 1 0 44252 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_487
timestamp 18001
transform 1 0 45908 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_491
timestamp 18001
transform 1 0 46276 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_500
timestamp 18001
transform 1 0 47104 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_503
timestamp 18001
transform 1 0 47380 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_521
timestamp 18001
transform 1 0 49036 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_556
timestamp 18001
transform 1 0 52256 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_566
timestamp 18001
transform 1 0 53176 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_572
timestamp 18001
transform 1 0 53728 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_605
timestamp 18001
transform 1 0 56764 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_615
timestamp 18001
transform 1 0 57684 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_617
timestamp 18001
transform 1 0 57868 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_3
timestamp 1636986456
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_15
timestamp 1636986456
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_27
timestamp 18001
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_29
timestamp 1636986456
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_41
timestamp 1636986456
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_53
timestamp 1636986456
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_65
timestamp 1636986456
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_77
timestamp 18001
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_83
timestamp 18001
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_85
timestamp 1636986456
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_97
timestamp 1636986456
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_109
timestamp 1636986456
transform 1 0 11132 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_121
timestamp 1636986456
transform 1 0 12236 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_133
timestamp 18001
transform 1 0 13340 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_139
timestamp 18001
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_141
timestamp 1636986456
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_153
timestamp 1636986456
transform 1 0 15180 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_165
timestamp 1636986456
transform 1 0 16284 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_177
timestamp 1636986456
transform 1 0 17388 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_189
timestamp 18001
transform 1 0 18492 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_195
timestamp 18001
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_204
timestamp 1636986456
transform 1 0 19872 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_216
timestamp 1636986456
transform 1 0 20976 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_228
timestamp 18001
transform 1 0 22080 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_243
timestamp 18001
transform 1 0 23460 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_251
timestamp 18001
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_253
timestamp 18001
transform 1 0 24380 0 1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_279
timestamp 1636986456
transform 1 0 26772 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_291
timestamp 18001
transform 1 0 27876 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_304
timestamp 18001
transform 1 0 29072 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_309
timestamp 18001
transform 1 0 29532 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_346
timestamp 18001
transform 1 0 32936 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_392
timestamp 1636986456
transform 1 0 37168 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_404
timestamp 18001
transform 1 0 38272 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_408
timestamp 18001
transform 1 0 38640 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_411
timestamp 18001
transform 1 0 38916 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_417
timestamp 18001
transform 1 0 39468 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_432
timestamp 18001
transform 1 0 40848 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_440
timestamp 18001
transform 1 0 41584 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_446
timestamp 18001
transform 1 0 42136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_469
timestamp 18001
transform 1 0 44252 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_473
timestamp 18001
transform 1 0 44620 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_477
timestamp 18001
transform 1 0 44988 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_485
timestamp 18001
transform 1 0 45724 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_515
timestamp 18001
transform 1 0 48484 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_526
timestamp 18001
transform 1 0 49496 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_533
timestamp 18001
transform 1 0 50140 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_546
timestamp 18001
transform 1 0 51336 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_557
timestamp 18001
transform 1 0 52348 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_565
timestamp 18001
transform 1 0 53084 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_582
timestamp 18001
transform 1 0 54648 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_589
timestamp 18001
transform 1 0 55292 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_593
timestamp 18001
transform 1 0 55660 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_596
timestamp 18001
transform 1 0 55936 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_604
timestamp 18001
transform 1 0 56672 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_615
timestamp 18001
transform 1 0 57684 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_623
timestamp 18001
transform 1 0 58420 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_3
timestamp 1636986456
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_15
timestamp 1636986456
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_27
timestamp 1636986456
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_39
timestamp 1636986456
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_51
timestamp 18001
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_55
timestamp 18001
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_57
timestamp 1636986456
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_69
timestamp 1636986456
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_81
timestamp 1636986456
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_93
timestamp 1636986456
transform 1 0 9660 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_105
timestamp 18001
transform 1 0 10764 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_111
timestamp 18001
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_113
timestamp 1636986456
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_125
timestamp 1636986456
transform 1 0 12604 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_137
timestamp 1636986456
transform 1 0 13708 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_149
timestamp 1636986456
transform 1 0 14812 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_161
timestamp 18001
transform 1 0 15916 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_167
timestamp 18001
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_169
timestamp 1636986456
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_181
timestamp 18001
transform 1 0 17756 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_212
timestamp 18001
transform 1 0 20608 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_220
timestamp 18001
transform 1 0 21344 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_245
timestamp 1636986456
transform 1 0 23644 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_277
timestamp 18001
transform 1 0 26588 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_281
timestamp 18001
transform 1 0 26956 0 -1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_315
timestamp 1636986456
transform 1 0 30084 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_327
timestamp 18001
transform 1 0 31188 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_344
timestamp 1636986456
transform 1 0 32752 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_356
timestamp 18001
transform 1 0 33856 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_364
timestamp 18001
transform 1 0 34592 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_381
timestamp 18001
transform 1 0 36156 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_389
timestamp 18001
transform 1 0 36892 0 -1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_404
timestamp 1636986456
transform 1 0 38272 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_416
timestamp 18001
transform 1 0 39376 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_437
timestamp 18001
transform 1 0 41308 0 -1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_466
timestamp 1636986456
transform 1 0 43976 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_478
timestamp 18001
transform 1 0 45080 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_484
timestamp 18001
transform 1 0 45632 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_503
timestamp 18001
transform 1 0 47380 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_507
timestamp 18001
transform 1 0 47748 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_515
timestamp 18001
transform 1 0 48484 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_519
timestamp 18001
transform 1 0 48852 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_540
timestamp 1636986456
transform 1 0 50784 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_552
timestamp 18001
transform 1 0 51888 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_561
timestamp 18001
transform 1 0 52716 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_570
timestamp 1636986456
transform 1 0 53544 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_582
timestamp 18001
transform 1 0 54648 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_617
timestamp 18001
transform 1 0 57868 0 -1 25024
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_3
timestamp 1636986456
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_15
timestamp 1636986456
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_27
timestamp 18001
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_29
timestamp 1636986456
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_41
timestamp 1636986456
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_53
timestamp 1636986456
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_65
timestamp 1636986456
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_77
timestamp 18001
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_83
timestamp 18001
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_85
timestamp 1636986456
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_97
timestamp 1636986456
transform 1 0 10028 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_109
timestamp 1636986456
transform 1 0 11132 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_121
timestamp 1636986456
transform 1 0 12236 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_133
timestamp 18001
transform 1 0 13340 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_139
timestamp 18001
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_141
timestamp 1636986456
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_153
timestamp 1636986456
transform 1 0 15180 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_165
timestamp 18001
transform 1 0 16284 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_173
timestamp 18001
transform 1 0 17020 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_197
timestamp 18001
transform 1 0 19228 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_212
timestamp 18001
transform 1 0 20608 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_251
timestamp 18001
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_253
timestamp 1636986456
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_265
timestamp 18001
transform 1 0 25484 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_280
timestamp 1636986456
transform 1 0 26864 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_292
timestamp 18001
transform 1 0 27968 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_307
timestamp 18001
transform 1 0 29348 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_311
timestamp 1636986456
transform 1 0 29716 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_323
timestamp 18001
transform 1 0 30820 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_354
timestamp 18001
transform 1 0 33672 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_362
timestamp 18001
transform 1 0 34408 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_397
timestamp 18001
transform 1 0 37628 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_418
timestamp 18001
transform 1 0 39560 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_429
timestamp 18001
transform 1 0 40572 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_472
timestamp 18001
transform 1 0 44528 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_477
timestamp 18001
transform 1 0 44988 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_483
timestamp 18001
transform 1 0 45540 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_520
timestamp 18001
transform 1 0 48944 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_543
timestamp 18001
transform 1 0 51060 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_583
timestamp 18001
transform 1 0 54740 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_587
timestamp 18001
transform 1 0 55108 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_603
timestamp 18001
transform 1 0 56580 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_622
timestamp 18001
transform 1 0 58328 0 1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_3
timestamp 1636986456
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_15
timestamp 1636986456
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_27
timestamp 1636986456
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_39
timestamp 1636986456
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_51
timestamp 18001
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_55
timestamp 18001
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_57
timestamp 1636986456
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_69
timestamp 1636986456
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_81
timestamp 1636986456
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_93
timestamp 1636986456
transform 1 0 9660 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_105
timestamp 18001
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_111
timestamp 18001
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_113
timestamp 1636986456
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_125
timestamp 1636986456
transform 1 0 12604 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_137
timestamp 1636986456
transform 1 0 13708 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_149
timestamp 1636986456
transform 1 0 14812 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_161
timestamp 18001
transform 1 0 15916 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_167
timestamp 18001
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_169
timestamp 1636986456
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_181
timestamp 1636986456
transform 1 0 17756 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_200
timestamp 1636986456
transform 1 0 19504 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_212
timestamp 1636986456
transform 1 0 20608 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_225
timestamp 18001
transform 1 0 21804 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_248
timestamp 18001
transform 1 0 23920 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_266
timestamp 18001
transform 1 0 25576 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_270
timestamp 18001
transform 1 0 25944 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_278
timestamp 18001
transform 1 0 26680 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_281
timestamp 18001
transform 1 0 26956 0 -1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_316
timestamp 1636986456
transform 1 0 30176 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_328
timestamp 18001
transform 1 0 31280 0 -1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_344
timestamp 1636986456
transform 1 0 32752 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_356
timestamp 1636986456
transform 1 0 33856 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_368
timestamp 18001
transform 1 0 34960 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_381
timestamp 18001
transform 1 0 36156 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_389
timestamp 18001
transform 1 0 36892 0 -1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_393
timestamp 1636986456
transform 1 0 37260 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_405
timestamp 18001
transform 1 0 38364 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_411
timestamp 18001
transform 1 0 38916 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_426
timestamp 1636986456
transform 1 0 40296 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_438
timestamp 18001
transform 1 0 41400 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_446
timestamp 18001
transform 1 0 42136 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_449
timestamp 18001
transform 1 0 42412 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_473
timestamp 18001
transform 1 0 44620 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_481
timestamp 18001
transform 1 0 45356 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_503
timestamp 18001
transform 1 0 47380 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_520
timestamp 18001
transform 1 0 48944 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_528
timestamp 18001
transform 1 0 49680 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_537
timestamp 18001
transform 1 0 50508 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_545
timestamp 18001
transform 1 0 51244 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_556
timestamp 18001
transform 1 0 52256 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_569
timestamp 18001
transform 1 0 53452 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_577
timestamp 18001
transform 1 0 54188 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_600
timestamp 18001
transform 1 0 56304 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_614
timestamp 18001
transform 1 0 57592 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_3
timestamp 1636986456
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_15
timestamp 1636986456
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_27
timestamp 18001
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_29
timestamp 1636986456
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_41
timestamp 1636986456
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_53
timestamp 1636986456
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_65
timestamp 1636986456
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_77
timestamp 18001
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_83
timestamp 18001
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_85
timestamp 1636986456
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_97
timestamp 1636986456
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_109
timestamp 1636986456
transform 1 0 11132 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_121
timestamp 1636986456
transform 1 0 12236 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_133
timestamp 18001
transform 1 0 13340 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_139
timestamp 18001
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_141
timestamp 1636986456
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_153
timestamp 1636986456
transform 1 0 15180 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_165
timestamp 1636986456
transform 1 0 16284 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_177
timestamp 1636986456
transform 1 0 17388 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_189
timestamp 18001
transform 1 0 18492 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_195
timestamp 18001
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_197
timestamp 1636986456
transform 1 0 19228 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_209
timestamp 1636986456
transform 1 0 20332 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_221
timestamp 1636986456
transform 1 0 21436 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_233
timestamp 18001
transform 1 0 22540 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_236
timestamp 1636986456
transform 1 0 22816 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_248
timestamp 18001
transform 1 0 23920 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_259
timestamp 18001
transform 1 0 24932 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_283
timestamp 18001
transform 1 0 27140 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_294
timestamp 18001
transform 1 0 28152 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_305
timestamp 18001
transform 1 0 29164 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_309
timestamp 18001
transform 1 0 29532 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_318
timestamp 1636986456
transform 1 0 30360 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_330
timestamp 18001
transform 1 0 31464 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_338
timestamp 18001
transform 1 0 32200 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_346
timestamp 1636986456
transform 1 0 32936 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_358
timestamp 18001
transform 1 0 34040 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_365
timestamp 18001
transform 1 0 34684 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_388
timestamp 1636986456
transform 1 0 36800 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_400
timestamp 18001
transform 1 0 37904 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_408
timestamp 18001
transform 1 0 38640 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_421
timestamp 18001
transform 1 0 39836 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_437
timestamp 1636986456
transform 1 0 41308 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_449
timestamp 1636986456
transform 1 0 42412 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_461
timestamp 1636986456
transform 1 0 43516 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_473
timestamp 18001
transform 1 0 44620 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_477
timestamp 18001
transform 1 0 44988 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_485
timestamp 18001
transform 1 0 45724 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_514
timestamp 18001
transform 1 0 48392 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_522
timestamp 18001
transform 1 0 49128 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_541
timestamp 1636986456
transform 1 0 50876 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_553
timestamp 18001
transform 1 0 51980 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_557
timestamp 18001
transform 1 0 52348 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_564
timestamp 18001
transform 1 0 52992 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_578
timestamp 18001
transform 1 0 54280 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_586
timestamp 18001
transform 1 0 55016 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_589
timestamp 1636986456
transform 1 0 55292 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_601
timestamp 1636986456
transform 1 0 56396 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_613
timestamp 18001
transform 1 0 57500 0 1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_3
timestamp 1636986456
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_15
timestamp 1636986456
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_27
timestamp 1636986456
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_39
timestamp 1636986456
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_51
timestamp 18001
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_55
timestamp 18001
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_57
timestamp 1636986456
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_69
timestamp 1636986456
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_81
timestamp 1636986456
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_93
timestamp 1636986456
transform 1 0 9660 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_105
timestamp 18001
transform 1 0 10764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_111
timestamp 18001
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_113
timestamp 1636986456
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_125
timestamp 1636986456
transform 1 0 12604 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_137
timestamp 1636986456
transform 1 0 13708 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_149
timestamp 1636986456
transform 1 0 14812 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_161
timestamp 18001
transform 1 0 15916 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_167
timestamp 18001
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_169
timestamp 1636986456
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_181
timestamp 1636986456
transform 1 0 17756 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_193
timestamp 1636986456
transform 1 0 18860 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_205
timestamp 1636986456
transform 1 0 19964 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_217
timestamp 18001
transform 1 0 21068 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_223
timestamp 18001
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_225
timestamp 1636986456
transform 1 0 21804 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_237
timestamp 18001
transform 1 0 22908 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_281
timestamp 18001
transform 1 0 26956 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_305
timestamp 1636986456
transform 1 0 29164 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_317
timestamp 1636986456
transform 1 0 30268 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_329
timestamp 18001
transform 1 0 31372 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_335
timestamp 18001
transform 1 0 31924 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_358
timestamp 18001
transform 1 0 34040 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_362
timestamp 18001
transform 1 0 34408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_391
timestamp 18001
transform 1 0 37076 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_393
timestamp 1636986456
transform 1 0 37260 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_405
timestamp 1636986456
transform 1 0 38364 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_417
timestamp 18001
transform 1 0 39468 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_421
timestamp 18001
transform 1 0 39836 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_427
timestamp 18001
transform 1 0 40388 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_440
timestamp 18001
transform 1 0 41584 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_449
timestamp 18001
transform 1 0 42412 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_455
timestamp 18001
transform 1 0 42964 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_466
timestamp 1636986456
transform 1 0 43976 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_478
timestamp 1636986456
transform 1 0 45080 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_490
timestamp 18001
transform 1 0 46184 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_496
timestamp 18001
transform 1 0 46736 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_507
timestamp 18001
transform 1 0 47748 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_545
timestamp 1636986456
transform 1 0 51244 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_557
timestamp 18001
transform 1 0 52348 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_581
timestamp 1636986456
transform 1 0 54556 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_593
timestamp 1636986456
transform 1 0 55660 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_605
timestamp 18001
transform 1 0 56764 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_613
timestamp 18001
transform 1 0 57500 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_617
timestamp 18001
transform 1 0 57868 0 -1 27200
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_3
timestamp 1636986456
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_15
timestamp 1636986456
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_27
timestamp 18001
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_29
timestamp 1636986456
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_41
timestamp 1636986456
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_53
timestamp 1636986456
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_65
timestamp 1636986456
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_77
timestamp 18001
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_83
timestamp 18001
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_85
timestamp 1636986456
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_97
timestamp 1636986456
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_109
timestamp 1636986456
transform 1 0 11132 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_121
timestamp 1636986456
transform 1 0 12236 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_133
timestamp 18001
transform 1 0 13340 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_139
timestamp 18001
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_141
timestamp 1636986456
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_153
timestamp 1636986456
transform 1 0 15180 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_165
timestamp 1636986456
transform 1 0 16284 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_177
timestamp 1636986456
transform 1 0 17388 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_189
timestamp 18001
transform 1 0 18492 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_195
timestamp 18001
transform 1 0 19044 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_197
timestamp 1636986456
transform 1 0 19228 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_209
timestamp 1636986456
transform 1 0 20332 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_221
timestamp 1636986456
transform 1 0 21436 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_233
timestamp 1636986456
transform 1 0 22540 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_245
timestamp 18001
transform 1 0 23644 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_251
timestamp 18001
transform 1 0 24196 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_253
timestamp 1636986456
transform 1 0 24380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_265
timestamp 1636986456
transform 1 0 25484 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_277
timestamp 1636986456
transform 1 0 26588 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_289
timestamp 1636986456
transform 1 0 27692 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_301
timestamp 18001
transform 1 0 28796 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_305
timestamp 18001
transform 1 0 29164 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_362
timestamp 18001
transform 1 0 34408 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_386
timestamp 18001
transform 1 0 36616 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_394
timestamp 18001
transform 1 0 37352 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_430
timestamp 18001
transform 1 0 40664 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_443
timestamp 18001
transform 1 0 41860 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_452
timestamp 18001
transform 1 0 42688 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_475
timestamp 18001
transform 1 0 44804 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_477
timestamp 1636986456
transform 1 0 44988 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_489
timestamp 18001
transform 1 0 46092 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_515
timestamp 18001
transform 1 0 48484 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_523
timestamp 18001
transform 1 0 49220 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_561
timestamp 1636986456
transform 1 0 52716 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_573
timestamp 1636986456
transform 1 0 53820 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_585
timestamp 18001
transform 1 0 54924 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_589
timestamp 1636986456
transform 1 0 55292 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_601
timestamp 1636986456
transform 1 0 56396 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_613
timestamp 1636986456
transform 1 0 57500 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_3
timestamp 1636986456
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_15
timestamp 1636986456
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_27
timestamp 1636986456
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_39
timestamp 1636986456
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_51
timestamp 18001
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_55
timestamp 18001
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_57
timestamp 1636986456
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_69
timestamp 1636986456
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_81
timestamp 1636986456
transform 1 0 8556 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_93
timestamp 1636986456
transform 1 0 9660 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_105
timestamp 18001
transform 1 0 10764 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_111
timestamp 18001
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_113
timestamp 1636986456
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_125
timestamp 1636986456
transform 1 0 12604 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_137
timestamp 1636986456
transform 1 0 13708 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_149
timestamp 1636986456
transform 1 0 14812 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_161
timestamp 18001
transform 1 0 15916 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_167
timestamp 18001
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_169
timestamp 1636986456
transform 1 0 16652 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_181
timestamp 1636986456
transform 1 0 17756 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_193
timestamp 1636986456
transform 1 0 18860 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_205
timestamp 1636986456
transform 1 0 19964 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_217
timestamp 18001
transform 1 0 21068 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_223
timestamp 18001
transform 1 0 21620 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_225
timestamp 1636986456
transform 1 0 21804 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_237
timestamp 1636986456
transform 1 0 22908 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_249
timestamp 1636986456
transform 1 0 24012 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_261
timestamp 1636986456
transform 1 0 25116 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_273
timestamp 18001
transform 1 0 26220 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_279
timestamp 18001
transform 1 0 26772 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_281
timestamp 1636986456
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_293
timestamp 18001
transform 1 0 28060 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_315
timestamp 1636986456
transform 1 0 30084 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_327
timestamp 18001
transform 1 0 31188 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_335
timestamp 18001
transform 1 0 31924 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_337
timestamp 1636986456
transform 1 0 32108 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_349
timestamp 1636986456
transform 1 0 33212 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_361
timestamp 1636986456
transform 1 0 34316 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_373
timestamp 1636986456
transform 1 0 35420 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_385
timestamp 18001
transform 1 0 36524 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_389
timestamp 18001
transform 1 0 36892 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_402
timestamp 1636986456
transform 1 0 38088 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_414
timestamp 18001
transform 1 0 39192 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_422
timestamp 18001
transform 1 0 39928 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_430
timestamp 1636986456
transform 1 0 40664 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_442
timestamp 18001
transform 1 0 41768 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_482
timestamp 18001
transform 1 0 45448 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_490
timestamp 18001
transform 1 0 46184 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_502
timestamp 18001
transform 1 0 47288 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_509
timestamp 1636986456
transform 1 0 47932 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_521
timestamp 18001
transform 1 0 49036 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_531
timestamp 18001
transform 1 0 49956 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_545
timestamp 1636986456
transform 1 0 51244 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_557
timestamp 18001
transform 1 0 52348 0 -1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_561
timestamp 1636986456
transform 1 0 52716 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_573
timestamp 1636986456
transform 1 0 53820 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_585
timestamp 1636986456
transform 1 0 54924 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_597
timestamp 1636986456
transform 1 0 56028 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_609
timestamp 18001
transform 1 0 57132 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_615
timestamp 18001
transform 1 0 57684 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_617
timestamp 18001
transform 1 0 57868 0 -1 28288
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_3
timestamp 1636986456
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_15
timestamp 1636986456
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_27
timestamp 18001
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_29
timestamp 1636986456
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_41
timestamp 1636986456
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_53
timestamp 1636986456
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_65
timestamp 1636986456
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_77
timestamp 18001
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_83
timestamp 18001
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_85
timestamp 1636986456
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_97
timestamp 1636986456
transform 1 0 10028 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_109
timestamp 1636986456
transform 1 0 11132 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_121
timestamp 1636986456
transform 1 0 12236 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_133
timestamp 18001
transform 1 0 13340 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_139
timestamp 18001
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_141
timestamp 1636986456
transform 1 0 14076 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_153
timestamp 1636986456
transform 1 0 15180 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_165
timestamp 1636986456
transform 1 0 16284 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_177
timestamp 1636986456
transform 1 0 17388 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_189
timestamp 18001
transform 1 0 18492 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_195
timestamp 18001
transform 1 0 19044 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_197
timestamp 1636986456
transform 1 0 19228 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_209
timestamp 1636986456
transform 1 0 20332 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_221
timestamp 1636986456
transform 1 0 21436 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_233
timestamp 1636986456
transform 1 0 22540 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_245
timestamp 18001
transform 1 0 23644 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_251
timestamp 18001
transform 1 0 24196 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_253
timestamp 1636986456
transform 1 0 24380 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_265
timestamp 18001
transform 1 0 25484 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_286
timestamp 1636986456
transform 1 0 27416 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_48_298
timestamp 18001
transform 1 0 28520 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_306
timestamp 18001
transform 1 0 29256 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_322
timestamp 1636986456
transform 1 0 30728 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_48_334
timestamp 18001
transform 1 0 31832 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_342
timestamp 18001
transform 1 0 32568 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_349
timestamp 1636986456
transform 1 0 33212 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_48_361
timestamp 18001
transform 1 0 34316 0 1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_365
timestamp 1636986456
transform 1 0 34684 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_377
timestamp 18001
transform 1 0 35788 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_48_402
timestamp 18001
transform 1 0 38088 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_412
timestamp 18001
transform 1 0 39008 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_421
timestamp 18001
transform 1 0 39836 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_430
timestamp 1636986456
transform 1 0 40664 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_442
timestamp 18001
transform 1 0 41768 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_450
timestamp 18001
transform 1 0 42504 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_475
timestamp 18001
transform 1 0 44804 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_482
timestamp 18001
transform 1 0 45448 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_487
timestamp 1636986456
transform 1 0 45908 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_499
timestamp 1636986456
transform 1 0 47012 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_511
timestamp 1636986456
transform 1 0 48116 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_523
timestamp 18001
transform 1 0 49220 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_531
timestamp 18001
transform 1 0 49956 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_533
timestamp 18001
transform 1 0 50140 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_543
timestamp 1636986456
transform 1 0 51060 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_555
timestamp 1636986456
transform 1 0 52164 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_567
timestamp 1636986456
transform 1 0 53268 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_579
timestamp 18001
transform 1 0 54372 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_587
timestamp 18001
transform 1 0 55108 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_589
timestamp 1636986456
transform 1 0 55292 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_601
timestamp 1636986456
transform 1 0 56396 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_613
timestamp 1636986456
transform 1 0 57500 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_3
timestamp 1636986456
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_15
timestamp 1636986456
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_27
timestamp 1636986456
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_39
timestamp 1636986456
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_51
timestamp 18001
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_55
timestamp 18001
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_57
timestamp 1636986456
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_69
timestamp 1636986456
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_81
timestamp 1636986456
transform 1 0 8556 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_93
timestamp 1636986456
transform 1 0 9660 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_105
timestamp 18001
transform 1 0 10764 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_111
timestamp 18001
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_113
timestamp 1636986456
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_125
timestamp 1636986456
transform 1 0 12604 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_137
timestamp 1636986456
transform 1 0 13708 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_149
timestamp 1636986456
transform 1 0 14812 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_161
timestamp 18001
transform 1 0 15916 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_167
timestamp 18001
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_169
timestamp 1636986456
transform 1 0 16652 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_181
timestamp 1636986456
transform 1 0 17756 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_193
timestamp 1636986456
transform 1 0 18860 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_205
timestamp 1636986456
transform 1 0 19964 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_217
timestamp 18001
transform 1 0 21068 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_223
timestamp 18001
transform 1 0 21620 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_225
timestamp 1636986456
transform 1 0 21804 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_237
timestamp 1636986456
transform 1 0 22908 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_249
timestamp 1636986456
transform 1 0 24012 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_261
timestamp 18001
transform 1 0 25116 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_269
timestamp 18001
transform 1 0 25852 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_277
timestamp 18001
transform 1 0 26588 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_320
timestamp 1636986456
transform 1 0 30544 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_332
timestamp 18001
transform 1 0 31648 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_377
timestamp 1636986456
transform 1 0 35788 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_389
timestamp 18001
transform 1 0 36892 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_393
timestamp 18001
transform 1 0 37260 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_417
timestamp 18001
transform 1 0 39468 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_421
timestamp 18001
transform 1 0 39836 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_443
timestamp 18001
transform 1 0 41860 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_447
timestamp 18001
transform 1 0 42228 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_449
timestamp 18001
transform 1 0 42412 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_453
timestamp 18001
transform 1 0 42780 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_470
timestamp 1636986456
transform 1 0 44344 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_482
timestamp 18001
transform 1 0 45448 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_494
timestamp 18001
transform 1 0 46552 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_502
timestamp 18001
transform 1 0 47288 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_505
timestamp 1636986456
transform 1 0 47564 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_517
timestamp 1636986456
transform 1 0 48668 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_529
timestamp 1636986456
transform 1 0 49772 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_541
timestamp 1636986456
transform 1 0 50876 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_553
timestamp 18001
transform 1 0 51980 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_559
timestamp 18001
transform 1 0 52532 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_561
timestamp 1636986456
transform 1 0 52716 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_573
timestamp 1636986456
transform 1 0 53820 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_585
timestamp 1636986456
transform 1 0 54924 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_597
timestamp 1636986456
transform 1 0 56028 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_609
timestamp 18001
transform 1 0 57132 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_615
timestamp 18001
transform 1 0 57684 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_617
timestamp 18001
transform 1 0 57868 0 -1 29376
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_3
timestamp 1636986456
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_15
timestamp 1636986456
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_27
timestamp 18001
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_29
timestamp 1636986456
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_41
timestamp 1636986456
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_53
timestamp 1636986456
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_65
timestamp 1636986456
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_77
timestamp 18001
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_83
timestamp 18001
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_85
timestamp 1636986456
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_97
timestamp 1636986456
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_109
timestamp 1636986456
transform 1 0 11132 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_121
timestamp 1636986456
transform 1 0 12236 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_133
timestamp 18001
transform 1 0 13340 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_139
timestamp 18001
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_141
timestamp 1636986456
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_153
timestamp 1636986456
transform 1 0 15180 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_165
timestamp 1636986456
transform 1 0 16284 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_177
timestamp 1636986456
transform 1 0 17388 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_189
timestamp 18001
transform 1 0 18492 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_195
timestamp 18001
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_197
timestamp 1636986456
transform 1 0 19228 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_209
timestamp 1636986456
transform 1 0 20332 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_221
timestamp 1636986456
transform 1 0 21436 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_240
timestamp 1636986456
transform 1 0 23184 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_261
timestamp 1636986456
transform 1 0 25116 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_273
timestamp 1636986456
transform 1 0 26220 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_285
timestamp 1636986456
transform 1 0 27324 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_297
timestamp 18001
transform 1 0 28428 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_307
timestamp 18001
transform 1 0 29348 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_313
timestamp 1636986456
transform 1 0 29900 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_325
timestamp 1636986456
transform 1 0 31004 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_50_337
timestamp 18001
transform 1 0 32108 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_345
timestamp 18001
transform 1 0 32844 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_353
timestamp 18001
transform 1 0 33580 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_363
timestamp 18001
transform 1 0 34500 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_370
timestamp 1636986456
transform 1 0 35144 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_382
timestamp 18001
transform 1 0 36248 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_50_390
timestamp 18001
transform 1 0 36984 0 1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_404
timestamp 1636986456
transform 1 0 38272 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_416
timestamp 18001
transform 1 0 39376 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_421
timestamp 18001
transform 1 0 39836 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_433
timestamp 1636986456
transform 1 0 40940 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_445
timestamp 18001
transform 1 0 42044 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_453
timestamp 18001
transform 1 0 42780 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_457
timestamp 18001
transform 1 0 43148 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_477
timestamp 18001
transform 1 0 44988 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_506
timestamp 1636986456
transform 1 0 47656 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_518
timestamp 1636986456
transform 1 0 48760 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_530
timestamp 18001
transform 1 0 49864 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_533
timestamp 1636986456
transform 1 0 50140 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_545
timestamp 1636986456
transform 1 0 51244 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_557
timestamp 1636986456
transform 1 0 52348 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_569
timestamp 1636986456
transform 1 0 53452 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_581
timestamp 18001
transform 1 0 54556 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_587
timestamp 18001
transform 1 0 55108 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_589
timestamp 1636986456
transform 1 0 55292 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_601
timestamp 1636986456
transform 1 0 56396 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_613
timestamp 1636986456
transform 1 0 57500 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_3
timestamp 1636986456
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_15
timestamp 1636986456
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_27
timestamp 1636986456
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_39
timestamp 1636986456
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_51
timestamp 18001
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_55
timestamp 18001
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_57
timestamp 1636986456
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_69
timestamp 1636986456
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_81
timestamp 1636986456
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_93
timestamp 1636986456
transform 1 0 9660 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_105
timestamp 18001
transform 1 0 10764 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_111
timestamp 18001
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_113
timestamp 1636986456
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_125
timestamp 1636986456
transform 1 0 12604 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_137
timestamp 1636986456
transform 1 0 13708 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_149
timestamp 1636986456
transform 1 0 14812 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_161
timestamp 18001
transform 1 0 15916 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_167
timestamp 18001
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_169
timestamp 1636986456
transform 1 0 16652 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_51_181
timestamp 18001
transform 1 0 17756 0 -1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_206
timestamp 1636986456
transform 1 0 20056 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_218
timestamp 18001
transform 1 0 21160 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_225
timestamp 18001
transform 1 0 21804 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_253
timestamp 18001
transform 1 0 24380 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_259
timestamp 18001
transform 1 0 24932 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_281
timestamp 1636986456
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_293
timestamp 1636986456
transform 1 0 28060 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_305
timestamp 1636986456
transform 1 0 29164 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_317
timestamp 1636986456
transform 1 0 30268 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_329
timestamp 18001
transform 1 0 31372 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_335
timestamp 18001
transform 1 0 31924 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_337
timestamp 18001
transform 1 0 32108 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_51_347
timestamp 18001
transform 1 0 33028 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_354
timestamp 18001
transform 1 0 33672 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_51_360
timestamp 18001
transform 1 0 34224 0 -1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_365
timestamp 1636986456
transform 1 0 34684 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_377
timestamp 1636986456
transform 1 0 35788 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_51_389
timestamp 18001
transform 1 0 36892 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_393
timestamp 18001
transform 1 0 37260 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_415
timestamp 1636986456
transform 1 0 39284 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_427
timestamp 1636986456
transform 1 0 40388 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_439
timestamp 18001
transform 1 0 41492 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_445
timestamp 18001
transform 1 0 42044 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_476
timestamp 1636986456
transform 1 0 44896 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_488
timestamp 1636986456
transform 1 0 46000 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_500
timestamp 18001
transform 1 0 47104 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_505
timestamp 1636986456
transform 1 0 47564 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_517
timestamp 1636986456
transform 1 0 48668 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_529
timestamp 1636986456
transform 1 0 49772 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_541
timestamp 1636986456
transform 1 0 50876 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_553
timestamp 18001
transform 1 0 51980 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_559
timestamp 18001
transform 1 0 52532 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_561
timestamp 1636986456
transform 1 0 52716 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_573
timestamp 1636986456
transform 1 0 53820 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_585
timestamp 1636986456
transform 1 0 54924 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_597
timestamp 1636986456
transform 1 0 56028 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_609
timestamp 18001
transform 1 0 57132 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_615
timestamp 18001
transform 1 0 57684 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_617
timestamp 18001
transform 1 0 57868 0 -1 30464
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_3
timestamp 1636986456
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_15
timestamp 1636986456
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_27
timestamp 18001
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_29
timestamp 1636986456
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_41
timestamp 1636986456
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_53
timestamp 1636986456
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_65
timestamp 1636986456
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_77
timestamp 18001
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_83
timestamp 18001
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_85
timestamp 1636986456
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_97
timestamp 1636986456
transform 1 0 10028 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_109
timestamp 1636986456
transform 1 0 11132 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_121
timestamp 1636986456
transform 1 0 12236 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_133
timestamp 18001
transform 1 0 13340 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_139
timestamp 18001
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_141
timestamp 1636986456
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52_153
timestamp 18001
transform 1 0 15180 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52_177
timestamp 18001
transform 1 0 17388 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_52_186
timestamp 18001
transform 1 0 18216 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_194
timestamp 18001
transform 1 0 18952 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_200
timestamp 1636986456
transform 1 0 19504 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_212
timestamp 1636986456
transform 1 0 20608 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_224
timestamp 1636986456
transform 1 0 21712 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_240
timestamp 1636986456
transform 1 0 23184 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52_253
timestamp 18001
transform 1 0 24380 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_257
timestamp 18001
transform 1 0 24748 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_290
timestamp 1636986456
transform 1 0 27784 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_302
timestamp 18001
transform 1 0 28888 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_52_309
timestamp 18001
transform 1 0 29532 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_52_322
timestamp 18001
transform 1 0 30728 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_345
timestamp 18001
transform 1 0 32844 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_363
timestamp 18001
transform 1 0 34500 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_52_373
timestamp 18001
transform 1 0 35420 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_381
timestamp 18001
transform 1 0 36156 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52_415
timestamp 18001
transform 1 0 39284 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_419
timestamp 18001
transform 1 0 39652 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_421
timestamp 1636986456
transform 1 0 39836 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_433
timestamp 1636986456
transform 1 0 40940 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_445
timestamp 1636986456
transform 1 0 42044 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_457
timestamp 1636986456
transform 1 0 43148 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_469
timestamp 18001
transform 1 0 44252 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_475
timestamp 18001
transform 1 0 44804 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_477
timestamp 1636986456
transform 1 0 44988 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_489
timestamp 1636986456
transform 1 0 46092 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_501
timestamp 1636986456
transform 1 0 47196 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_513
timestamp 1636986456
transform 1 0 48300 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_525
timestamp 18001
transform 1 0 49404 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_531
timestamp 18001
transform 1 0 49956 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_533
timestamp 1636986456
transform 1 0 50140 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_545
timestamp 1636986456
transform 1 0 51244 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_557
timestamp 1636986456
transform 1 0 52348 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_569
timestamp 1636986456
transform 1 0 53452 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_581
timestamp 18001
transform 1 0 54556 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_587
timestamp 18001
transform 1 0 55108 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_589
timestamp 1636986456
transform 1 0 55292 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_601
timestamp 1636986456
transform 1 0 56396 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_613
timestamp 1636986456
transform 1 0 57500 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_3
timestamp 1636986456
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_15
timestamp 1636986456
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_27
timestamp 1636986456
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_39
timestamp 1636986456
transform 1 0 4692 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_51
timestamp 18001
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_55
timestamp 18001
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_57
timestamp 1636986456
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_69
timestamp 1636986456
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_81
timestamp 1636986456
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_93
timestamp 1636986456
transform 1 0 9660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_105
timestamp 18001
transform 1 0 10764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_111
timestamp 18001
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_113
timestamp 1636986456
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_125
timestamp 1636986456
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53_137
timestamp 18001
transform 1 0 13708 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53_166
timestamp 18001
transform 1 0 16376 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_188
timestamp 18001
transform 1 0 18400 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53_212
timestamp 18001
transform 1 0 20608 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_223
timestamp 18001
transform 1 0 21620 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_241
timestamp 18001
transform 1 0 23276 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_53_248
timestamp 18001
transform 1 0 23920 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_279
timestamp 18001
transform 1 0 26772 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_281
timestamp 1636986456
transform 1 0 26956 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_293
timestamp 18001
transform 1 0 28060 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53_317
timestamp 18001
transform 1 0 30268 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_332
timestamp 18001
transform 1 0 31648 0 -1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_337
timestamp 1636986456
transform 1 0 32108 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_349
timestamp 18001
transform 1 0 33212 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_368
timestamp 1636986456
transform 1 0 34960 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_380
timestamp 18001
transform 1 0 36064 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_384
timestamp 18001
transform 1 0 36432 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_413
timestamp 1636986456
transform 1 0 39100 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_425
timestamp 1636986456
transform 1 0 40204 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_53_437
timestamp 18001
transform 1 0 41308 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53_445
timestamp 18001
transform 1 0 42044 0 -1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_449
timestamp 1636986456
transform 1 0 42412 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_461
timestamp 1636986456
transform 1 0 43516 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_473
timestamp 1636986456
transform 1 0 44620 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_485
timestamp 1636986456
transform 1 0 45724 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_497
timestamp 18001
transform 1 0 46828 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_503
timestamp 18001
transform 1 0 47380 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_505
timestamp 1636986456
transform 1 0 47564 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_517
timestamp 1636986456
transform 1 0 48668 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_529
timestamp 1636986456
transform 1 0 49772 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_541
timestamp 1636986456
transform 1 0 50876 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_553
timestamp 18001
transform 1 0 51980 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_559
timestamp 18001
transform 1 0 52532 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_561
timestamp 1636986456
transform 1 0 52716 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_573
timestamp 1636986456
transform 1 0 53820 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_585
timestamp 1636986456
transform 1 0 54924 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_597
timestamp 1636986456
transform 1 0 56028 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_609
timestamp 18001
transform 1 0 57132 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_615
timestamp 18001
transform 1 0 57684 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_53_617
timestamp 18001
transform 1 0 57868 0 -1 31552
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_3
timestamp 1636986456
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_15
timestamp 1636986456
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_27
timestamp 18001
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_29
timestamp 1636986456
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_41
timestamp 1636986456
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_53
timestamp 1636986456
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_65
timestamp 1636986456
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_77
timestamp 18001
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_83
timestamp 18001
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_85
timestamp 1636986456
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_97
timestamp 1636986456
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_109
timestamp 1636986456
transform 1 0 11132 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_121
timestamp 1636986456
transform 1 0 12236 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_133
timestamp 18001
transform 1 0 13340 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_139
timestamp 18001
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_141
timestamp 1636986456
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_153
timestamp 18001
transform 1 0 15180 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_54_188
timestamp 18001
transform 1 0 18400 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_54_203
timestamp 18001
transform 1 0 19780 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_207
timestamp 18001
transform 1 0 20148 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_54_248
timestamp 18001
transform 1 0 23920 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_54_261
timestamp 18001
transform 1 0 25116 0 1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_275
timestamp 1636986456
transform 1 0 26404 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_287
timestamp 1636986456
transform 1 0 27508 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_54_299
timestamp 18001
transform 1 0 28612 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_303
timestamp 18001
transform 1 0 28980 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_54_342
timestamp 18001
transform 1 0 32568 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_356
timestamp 18001
transform 1 0 33856 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_363
timestamp 18001
transform 1 0 34500 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_365
timestamp 1636986456
transform 1 0 34684 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_377
timestamp 1636986456
transform 1 0 35788 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_389
timestamp 18001
transform 1 0 36892 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_403
timestamp 1636986456
transform 1 0 38180 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_54_415
timestamp 18001
transform 1 0 39284 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_419
timestamp 18001
transform 1 0 39652 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_421
timestamp 1636986456
transform 1 0 39836 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_433
timestamp 1636986456
transform 1 0 40940 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_445
timestamp 1636986456
transform 1 0 42044 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_457
timestamp 1636986456
transform 1 0 43148 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_469
timestamp 18001
transform 1 0 44252 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_475
timestamp 18001
transform 1 0 44804 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_477
timestamp 1636986456
transform 1 0 44988 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_489
timestamp 1636986456
transform 1 0 46092 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_501
timestamp 1636986456
transform 1 0 47196 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_513
timestamp 1636986456
transform 1 0 48300 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_525
timestamp 18001
transform 1 0 49404 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_531
timestamp 18001
transform 1 0 49956 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_533
timestamp 1636986456
transform 1 0 50140 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_545
timestamp 1636986456
transform 1 0 51244 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_557
timestamp 1636986456
transform 1 0 52348 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_569
timestamp 1636986456
transform 1 0 53452 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_581
timestamp 18001
transform 1 0 54556 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_587
timestamp 18001
transform 1 0 55108 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_589
timestamp 1636986456
transform 1 0 55292 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_601
timestamp 1636986456
transform 1 0 56396 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_613
timestamp 1636986456
transform 1 0 57500 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_3
timestamp 1636986456
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_15
timestamp 1636986456
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_27
timestamp 1636986456
transform 1 0 3588 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_39
timestamp 1636986456
transform 1 0 4692 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_55_51
timestamp 18001
transform 1 0 5796 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_55
timestamp 18001
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_57
timestamp 1636986456
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_69
timestamp 1636986456
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_81
timestamp 1636986456
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_93
timestamp 1636986456
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_105
timestamp 18001
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_111
timestamp 18001
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_113
timestamp 1636986456
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_125
timestamp 1636986456
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_137
timestamp 1636986456
transform 1 0 13708 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_149
timestamp 1636986456
transform 1 0 14812 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_184
timestamp 1636986456
transform 1 0 18032 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_196
timestamp 1636986456
transform 1 0 19136 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_208
timestamp 1636986456
transform 1 0 20240 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_55_220
timestamp 18001
transform 1 0 21344 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_225
timestamp 1636986456
transform 1 0 21804 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_237
timestamp 1636986456
transform 1 0 22908 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_249
timestamp 1636986456
transform 1 0 24012 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_261
timestamp 1636986456
transform 1 0 25116 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_286
timestamp 1636986456
transform 1 0 27416 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_298
timestamp 1636986456
transform 1 0 28520 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_55_310
timestamp 18001
transform 1 0 29624 0 -1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_322
timestamp 1636986456
transform 1 0 30728 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_55_334
timestamp 18001
transform 1 0 31832 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_55_337
timestamp 18001
transform 1 0 32108 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_55_345
timestamp 18001
transform 1 0 32844 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_55_371
timestamp 18001
transform 1 0 35236 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_379
timestamp 18001
transform 1 0 35972 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_391
timestamp 18001
transform 1 0 37076 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_393
timestamp 1636986456
transform 1 0 37260 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_405
timestamp 1636986456
transform 1 0 38364 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_417
timestamp 1636986456
transform 1 0 39468 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_429
timestamp 1636986456
transform 1 0 40572 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_441
timestamp 18001
transform 1 0 41676 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_447
timestamp 18001
transform 1 0 42228 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_449
timestamp 1636986456
transform 1 0 42412 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_461
timestamp 1636986456
transform 1 0 43516 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_473
timestamp 1636986456
transform 1 0 44620 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_485
timestamp 1636986456
transform 1 0 45724 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_497
timestamp 18001
transform 1 0 46828 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_503
timestamp 18001
transform 1 0 47380 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_505
timestamp 1636986456
transform 1 0 47564 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_517
timestamp 1636986456
transform 1 0 48668 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_529
timestamp 1636986456
transform 1 0 49772 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_541
timestamp 1636986456
transform 1 0 50876 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_553
timestamp 18001
transform 1 0 51980 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_559
timestamp 18001
transform 1 0 52532 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_561
timestamp 1636986456
transform 1 0 52716 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_573
timestamp 1636986456
transform 1 0 53820 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_585
timestamp 1636986456
transform 1 0 54924 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_597
timestamp 1636986456
transform 1 0 56028 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_609
timestamp 18001
transform 1 0 57132 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_615
timestamp 18001
transform 1 0 57684 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_55_617
timestamp 18001
transform 1 0 57868 0 -1 32640
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_3
timestamp 1636986456
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_15
timestamp 1636986456
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_27
timestamp 18001
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_29
timestamp 1636986456
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_41
timestamp 1636986456
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_53
timestamp 1636986456
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_65
timestamp 1636986456
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_77
timestamp 18001
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_83
timestamp 18001
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_85
timestamp 1636986456
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_97
timestamp 1636986456
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_109
timestamp 1636986456
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_121
timestamp 1636986456
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_133
timestamp 18001
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_139
timestamp 18001
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_56_141
timestamp 18001
transform 1 0 14076 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_56_164
timestamp 18001
transform 1 0 16192 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_56_174
timestamp 18001
transform 1 0 17112 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_178
timestamp 18001
transform 1 0 17480 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_56_192
timestamp 18001
transform 1 0 18768 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_56_205
timestamp 18001
transform 1 0 19964 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_213
timestamp 18001
transform 1 0 20700 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_234
timestamp 18001
transform 1 0 22632 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_56_243
timestamp 18001
transform 1 0 23460 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_251
timestamp 18001
transform 1 0 24196 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_56_262
timestamp 18001
transform 1 0 25208 0 1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_291
timestamp 1636986456
transform 1 0 27876 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_56_303
timestamp 18001
transform 1 0 28980 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_307
timestamp 18001
transform 1 0 29348 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_56_309
timestamp 18001
transform 1 0 29532 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_317
timestamp 18001
transform 1 0 30268 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_325
timestamp 1636986456
transform 1 0 31004 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_337
timestamp 1636986456
transform 1 0 32108 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_365
timestamp 1636986456
transform 1 0 34684 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_404
timestamp 1636986456
transform 1 0 38272 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_56_416
timestamp 18001
transform 1 0 39376 0 1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_421
timestamp 1636986456
transform 1 0 39836 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_433
timestamp 1636986456
transform 1 0 40940 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_445
timestamp 1636986456
transform 1 0 42044 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_457
timestamp 1636986456
transform 1 0 43148 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_469
timestamp 18001
transform 1 0 44252 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_475
timestamp 18001
transform 1 0 44804 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_477
timestamp 1636986456
transform 1 0 44988 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_489
timestamp 1636986456
transform 1 0 46092 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_501
timestamp 1636986456
transform 1 0 47196 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_513
timestamp 1636986456
transform 1 0 48300 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_525
timestamp 18001
transform 1 0 49404 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_531
timestamp 18001
transform 1 0 49956 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_533
timestamp 1636986456
transform 1 0 50140 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_545
timestamp 1636986456
transform 1 0 51244 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_557
timestamp 1636986456
transform 1 0 52348 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_569
timestamp 1636986456
transform 1 0 53452 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_581
timestamp 18001
transform 1 0 54556 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_587
timestamp 18001
transform 1 0 55108 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_589
timestamp 1636986456
transform 1 0 55292 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_601
timestamp 1636986456
transform 1 0 56396 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_613
timestamp 1636986456
transform 1 0 57500 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_3
timestamp 1636986456
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_15
timestamp 1636986456
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_27
timestamp 1636986456
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_39
timestamp 1636986456
transform 1 0 4692 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57_51
timestamp 18001
transform 1 0 5796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_55
timestamp 18001
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_57
timestamp 1636986456
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_69
timestamp 1636986456
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_81
timestamp 1636986456
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_93
timestamp 1636986456
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_105
timestamp 18001
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_111
timestamp 18001
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_113
timestamp 1636986456
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_125
timestamp 1636986456
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_137
timestamp 1636986456
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_149
timestamp 1636986456
transform 1 0 14812 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_161
timestamp 18001
transform 1 0 15916 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_167
timestamp 18001
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_57_169
timestamp 18001
transform 1 0 16652 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57_195
timestamp 18001
transform 1 0 19044 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_203
timestamp 18001
transform 1 0 19780 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_231
timestamp 18001
transform 1 0 22356 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57_245
timestamp 18001
transform 1 0 23644 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57_258
timestamp 18001
transform 1 0 24840 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_286
timestamp 1636986456
transform 1 0 27416 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_298
timestamp 18001
transform 1 0 28520 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_330
timestamp 18001
transform 1 0 31464 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_337
timestamp 18001
transform 1 0 32108 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_343
timestamp 18001
transform 1 0 32660 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_359
timestamp 1636986456
transform 1 0 34132 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_371
timestamp 1636986456
transform 1 0 35236 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57_383
timestamp 18001
transform 1 0 36340 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_413
timestamp 1636986456
transform 1 0 39100 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_425
timestamp 1636986456
transform 1 0 40204 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57_437
timestamp 18001
transform 1 0 41308 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_57_445
timestamp 18001
transform 1 0 42044 0 -1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_449
timestamp 1636986456
transform 1 0 42412 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_461
timestamp 1636986456
transform 1 0 43516 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_473
timestamp 1636986456
transform 1 0 44620 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_485
timestamp 1636986456
transform 1 0 45724 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_497
timestamp 18001
transform 1 0 46828 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_503
timestamp 18001
transform 1 0 47380 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_505
timestamp 1636986456
transform 1 0 47564 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_517
timestamp 1636986456
transform 1 0 48668 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_529
timestamp 1636986456
transform 1 0 49772 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_541
timestamp 1636986456
transform 1 0 50876 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_553
timestamp 18001
transform 1 0 51980 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_559
timestamp 18001
transform 1 0 52532 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_561
timestamp 1636986456
transform 1 0 52716 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_573
timestamp 1636986456
transform 1 0 53820 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_585
timestamp 1636986456
transform 1 0 54924 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_597
timestamp 1636986456
transform 1 0 56028 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_609
timestamp 18001
transform 1 0 57132 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_615
timestamp 18001
transform 1 0 57684 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57_617
timestamp 18001
transform 1 0 57868 0 -1 33728
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_3
timestamp 1636986456
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_15
timestamp 1636986456
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_27
timestamp 18001
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_29
timestamp 1636986456
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_41
timestamp 1636986456
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_53
timestamp 1636986456
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_65
timestamp 1636986456
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_77
timestamp 18001
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_83
timestamp 18001
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_85
timestamp 1636986456
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_97
timestamp 1636986456
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_109
timestamp 1636986456
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_121
timestamp 1636986456
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_133
timestamp 18001
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_139
timestamp 18001
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_141
timestamp 1636986456
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_153
timestamp 1636986456
transform 1 0 15180 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_165
timestamp 1636986456
transform 1 0 16284 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58_177
timestamp 18001
transform 1 0 17388 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_58_186
timestamp 18001
transform 1 0 18216 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58_194
timestamp 18001
transform 1 0 18952 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_58_197
timestamp 18001
transform 1 0 19228 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_58_205
timestamp 18001
transform 1 0 19964 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58_220
timestamp 18001
transform 1 0 21344 0 1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_227
timestamp 1636986456
transform 1 0 21988 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_58_239
timestamp 18001
transform 1 0 23092 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_247
timestamp 18001
transform 1 0 23828 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_58_253
timestamp 18001
transform 1 0 24380 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_273
timestamp 18001
transform 1 0 26220 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_278
timestamp 18001
transform 1 0 26680 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_287
timestamp 1636986456
transform 1 0 27508 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_58_299
timestamp 18001
transform 1 0 28612 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_307
timestamp 18001
transform 1 0 29348 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_58_309
timestamp 18001
transform 1 0 29532 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_58_317
timestamp 18001
transform 1 0 30268 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_58_327
timestamp 18001
transform 1 0 31188 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_350
timestamp 18001
transform 1 0 33304 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_363
timestamp 18001
transform 1 0 34500 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_365
timestamp 1636986456
transform 1 0 34684 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_377
timestamp 1636986456
transform 1 0 35788 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58_389
timestamp 18001
transform 1 0 36892 0 1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_393
timestamp 1636986456
transform 1 0 37260 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_405
timestamp 1636986456
transform 1 0 38364 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_58_417
timestamp 18001
transform 1 0 39468 0 1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_421
timestamp 1636986456
transform 1 0 39836 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_433
timestamp 1636986456
transform 1 0 40940 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_445
timestamp 1636986456
transform 1 0 42044 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_457
timestamp 1636986456
transform 1 0 43148 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_469
timestamp 18001
transform 1 0 44252 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_475
timestamp 18001
transform 1 0 44804 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_477
timestamp 1636986456
transform 1 0 44988 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_489
timestamp 1636986456
transform 1 0 46092 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_501
timestamp 1636986456
transform 1 0 47196 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_513
timestamp 1636986456
transform 1 0 48300 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_525
timestamp 18001
transform 1 0 49404 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_531
timestamp 18001
transform 1 0 49956 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_533
timestamp 1636986456
transform 1 0 50140 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_545
timestamp 1636986456
transform 1 0 51244 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_557
timestamp 1636986456
transform 1 0 52348 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_569
timestamp 1636986456
transform 1 0 53452 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_581
timestamp 18001
transform 1 0 54556 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_587
timestamp 18001
transform 1 0 55108 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_589
timestamp 1636986456
transform 1 0 55292 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_601
timestamp 1636986456
transform 1 0 56396 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_613
timestamp 1636986456
transform 1 0 57500 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_3
timestamp 1636986456
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_15
timestamp 1636986456
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_27
timestamp 1636986456
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_39
timestamp 1636986456
transform 1 0 4692 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_59_51
timestamp 18001
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_55
timestamp 18001
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_57
timestamp 1636986456
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_69
timestamp 1636986456
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_81
timestamp 1636986456
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_93
timestamp 1636986456
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_105
timestamp 18001
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_111
timestamp 18001
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_113
timestamp 1636986456
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_125
timestamp 1636986456
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_137
timestamp 1636986456
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_149
timestamp 1636986456
transform 1 0 14812 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_161
timestamp 18001
transform 1 0 15916 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_167
timestamp 18001
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_196
timestamp 1636986456
transform 1 0 19136 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_59_208
timestamp 18001
transform 1 0 20240 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_216
timestamp 18001
transform 1 0 20976 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_59_220
timestamp 18001
transform 1 0 21344 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_59_225
timestamp 18001
transform 1 0 21804 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_233
timestamp 18001
transform 1 0 22540 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_59_236
timestamp 18001
transform 1 0 22816 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_59_267
timestamp 18001
transform 1 0 25668 0 -1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_286
timestamp 1636986456
transform 1 0 27416 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_298
timestamp 1636986456
transform 1 0 28520 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_310
timestamp 18001
transform 1 0 29624 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_59_337
timestamp 18001
transform 1 0 32108 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_345
timestamp 18001
transform 1 0 32844 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_367
timestamp 1636986456
transform 1 0 34868 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_379
timestamp 1636986456
transform 1 0 35972 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_391
timestamp 18001
transform 1 0 37076 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_393
timestamp 1636986456
transform 1 0 37260 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_405
timestamp 1636986456
transform 1 0 38364 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_417
timestamp 1636986456
transform 1 0 39468 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_429
timestamp 1636986456
transform 1 0 40572 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_441
timestamp 18001
transform 1 0 41676 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_447
timestamp 18001
transform 1 0 42228 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_449
timestamp 1636986456
transform 1 0 42412 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_461
timestamp 1636986456
transform 1 0 43516 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_473
timestamp 1636986456
transform 1 0 44620 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_485
timestamp 1636986456
transform 1 0 45724 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_497
timestamp 18001
transform 1 0 46828 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_503
timestamp 18001
transform 1 0 47380 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_505
timestamp 1636986456
transform 1 0 47564 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_517
timestamp 1636986456
transform 1 0 48668 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_529
timestamp 1636986456
transform 1 0 49772 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_541
timestamp 1636986456
transform 1 0 50876 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_553
timestamp 18001
transform 1 0 51980 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_559
timestamp 18001
transform 1 0 52532 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_561
timestamp 1636986456
transform 1 0 52716 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_573
timestamp 1636986456
transform 1 0 53820 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_585
timestamp 1636986456
transform 1 0 54924 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_597
timestamp 1636986456
transform 1 0 56028 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_609
timestamp 18001
transform 1 0 57132 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_615
timestamp 18001
transform 1 0 57684 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_59_617
timestamp 18001
transform 1 0 57868 0 -1 34816
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_3
timestamp 1636986456
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_15
timestamp 1636986456
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_27
timestamp 18001
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_29
timestamp 1636986456
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_41
timestamp 1636986456
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_53
timestamp 1636986456
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_65
timestamp 1636986456
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_77
timestamp 18001
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_83
timestamp 18001
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_85
timestamp 1636986456
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_97
timestamp 1636986456
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_109
timestamp 1636986456
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_121
timestamp 1636986456
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_133
timestamp 18001
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_139
timestamp 18001
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_141
timestamp 1636986456
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_153
timestamp 1636986456
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_165
timestamp 1636986456
transform 1 0 16284 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_177
timestamp 18001
transform 1 0 17388 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_60_191
timestamp 18001
transform 1 0 18676 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_195
timestamp 18001
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_197
timestamp 1636986456
transform 1 0 19228 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_209
timestamp 1636986456
transform 1 0 20332 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_60_221
timestamp 18001
transform 1 0 21436 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_234
timestamp 18001
transform 1 0 22632 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_245
timestamp 18001
transform 1 0 23644 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_251
timestamp 18001
transform 1 0 24196 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_253
timestamp 18001
transform 1 0 24380 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_307
timestamp 18001
transform 1 0 29348 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_309
timestamp 1636986456
transform 1 0 29532 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_60_321
timestamp 18001
transform 1 0 30636 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_60_328
timestamp 18001
transform 1 0 31280 0 1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_335
timestamp 1636986456
transform 1 0 31924 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_347
timestamp 1636986456
transform 1 0 33028 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_60_359
timestamp 18001
transform 1 0 34132 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_363
timestamp 18001
transform 1 0 34500 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_365
timestamp 1636986456
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_377
timestamp 1636986456
transform 1 0 35788 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_389
timestamp 1636986456
transform 1 0 36892 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_401
timestamp 1636986456
transform 1 0 37996 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_413
timestamp 18001
transform 1 0 39100 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_419
timestamp 18001
transform 1 0 39652 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_421
timestamp 1636986456
transform 1 0 39836 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_433
timestamp 1636986456
transform 1 0 40940 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_445
timestamp 1636986456
transform 1 0 42044 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_457
timestamp 1636986456
transform 1 0 43148 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_469
timestamp 18001
transform 1 0 44252 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_475
timestamp 18001
transform 1 0 44804 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_477
timestamp 1636986456
transform 1 0 44988 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_489
timestamp 1636986456
transform 1 0 46092 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_501
timestamp 1636986456
transform 1 0 47196 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_513
timestamp 1636986456
transform 1 0 48300 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_525
timestamp 18001
transform 1 0 49404 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_531
timestamp 18001
transform 1 0 49956 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_533
timestamp 1636986456
transform 1 0 50140 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_545
timestamp 1636986456
transform 1 0 51244 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_557
timestamp 1636986456
transform 1 0 52348 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_569
timestamp 1636986456
transform 1 0 53452 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_581
timestamp 18001
transform 1 0 54556 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_587
timestamp 18001
transform 1 0 55108 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_589
timestamp 1636986456
transform 1 0 55292 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_601
timestamp 1636986456
transform 1 0 56396 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_613
timestamp 1636986456
transform 1 0 57500 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_3
timestamp 1636986456
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_15
timestamp 1636986456
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_27
timestamp 1636986456
transform 1 0 3588 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_39
timestamp 1636986456
transform 1 0 4692 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_61_51
timestamp 18001
transform 1 0 5796 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_55
timestamp 18001
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_57
timestamp 1636986456
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_69
timestamp 1636986456
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_81
timestamp 1636986456
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_93
timestamp 1636986456
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_105
timestamp 18001
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_111
timestamp 18001
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_113
timestamp 1636986456
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_125
timestamp 1636986456
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_137
timestamp 1636986456
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_149
timestamp 1636986456
transform 1 0 14812 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_161
timestamp 18001
transform 1 0 15916 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_167
timestamp 18001
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_169
timestamp 1636986456
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_181
timestamp 1636986456
transform 1 0 17756 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_193
timestamp 1636986456
transform 1 0 18860 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_205
timestamp 1636986456
transform 1 0 19964 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_217
timestamp 18001
transform 1 0 21068 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_223
timestamp 18001
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_61_251
timestamp 18001
transform 1 0 24196 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_259
timestamp 18001
transform 1 0 24932 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_281
timestamp 1636986456
transform 1 0 26956 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_61_293
timestamp 18001
transform 1 0 28060 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_297
timestamp 18001
transform 1 0 28428 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_314
timestamp 1636986456
transform 1 0 29992 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_61_326
timestamp 18001
transform 1 0 31096 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_61_334
timestamp 18001
transform 1 0 31832 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_337
timestamp 1636986456
transform 1 0 32108 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_349
timestamp 1636986456
transform 1 0 33212 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_361
timestamp 1636986456
transform 1 0 34316 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_373
timestamp 1636986456
transform 1 0 35420 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_385
timestamp 18001
transform 1 0 36524 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_391
timestamp 18001
transform 1 0 37076 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_393
timestamp 1636986456
transform 1 0 37260 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_405
timestamp 1636986456
transform 1 0 38364 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_417
timestamp 1636986456
transform 1 0 39468 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_429
timestamp 1636986456
transform 1 0 40572 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_441
timestamp 18001
transform 1 0 41676 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_447
timestamp 18001
transform 1 0 42228 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_449
timestamp 1636986456
transform 1 0 42412 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_461
timestamp 1636986456
transform 1 0 43516 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_473
timestamp 1636986456
transform 1 0 44620 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_485
timestamp 1636986456
transform 1 0 45724 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_497
timestamp 18001
transform 1 0 46828 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_503
timestamp 18001
transform 1 0 47380 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_505
timestamp 1636986456
transform 1 0 47564 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_517
timestamp 1636986456
transform 1 0 48668 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_529
timestamp 1636986456
transform 1 0 49772 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_541
timestamp 1636986456
transform 1 0 50876 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_553
timestamp 18001
transform 1 0 51980 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_559
timestamp 18001
transform 1 0 52532 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_561
timestamp 1636986456
transform 1 0 52716 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_573
timestamp 1636986456
transform 1 0 53820 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_585
timestamp 1636986456
transform 1 0 54924 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_597
timestamp 1636986456
transform 1 0 56028 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_609
timestamp 18001
transform 1 0 57132 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_615
timestamp 18001
transform 1 0 57684 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_61_617
timestamp 18001
transform 1 0 57868 0 -1 35904
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_3
timestamp 1636986456
transform 1 0 1380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_15
timestamp 1636986456
transform 1 0 2484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_27
timestamp 18001
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_29
timestamp 1636986456
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_41
timestamp 1636986456
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_53
timestamp 1636986456
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_65
timestamp 1636986456
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_77
timestamp 18001
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_83
timestamp 18001
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_85
timestamp 1636986456
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_97
timestamp 1636986456
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_109
timestamp 1636986456
transform 1 0 11132 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_121
timestamp 1636986456
transform 1 0 12236 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_133
timestamp 18001
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_139
timestamp 18001
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_141
timestamp 1636986456
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_153
timestamp 1636986456
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_165
timestamp 1636986456
transform 1 0 16284 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_177
timestamp 1636986456
transform 1 0 17388 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_189
timestamp 18001
transform 1 0 18492 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_195
timestamp 18001
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_197
timestamp 1636986456
transform 1 0 19228 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_209
timestamp 1636986456
transform 1 0 20332 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_221
timestamp 1636986456
transform 1 0 21436 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_62_233
timestamp 18001
transform 1 0 22540 0 1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_264
timestamp 1636986456
transform 1 0 25392 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_276
timestamp 1636986456
transform 1 0 26496 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_288
timestamp 1636986456
transform 1 0 27600 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_318
timestamp 1636986456
transform 1 0 30360 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_330
timestamp 18001
transform 1 0 31464 0 1 35904
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_339
timestamp 1636986456
transform 1 0 32292 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_351
timestamp 1636986456
transform 1 0 33396 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_363
timestamp 18001
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_365
timestamp 18001
transform 1 0 34684 0 1 35904
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_374
timestamp 1636986456
transform 1 0 35512 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_386
timestamp 18001
transform 1 0 36616 0 1 35904
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_395
timestamp 1636986456
transform 1 0 37444 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_407
timestamp 1636986456
transform 1 0 38548 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_419
timestamp 18001
transform 1 0 39652 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_421
timestamp 1636986456
transform 1 0 39836 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_433
timestamp 1636986456
transform 1 0 40940 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_62_445
timestamp 18001
transform 1 0 42044 0 1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_451
timestamp 1636986456
transform 1 0 42596 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_463
timestamp 1636986456
transform 1 0 43700 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_475
timestamp 18001
transform 1 0 44804 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_477
timestamp 1636986456
transform 1 0 44988 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_489
timestamp 18001
transform 1 0 46092 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_493
timestamp 1636986456
transform 1 0 46460 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_505
timestamp 1636986456
transform 1 0 47564 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_517
timestamp 1636986456
transform 1 0 48668 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_62_529
timestamp 18001
transform 1 0 49772 0 1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_533
timestamp 1636986456
transform 1 0 50140 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_545
timestamp 1636986456
transform 1 0 51244 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_557
timestamp 1636986456
transform 1 0 52348 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_569
timestamp 1636986456
transform 1 0 53452 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_581
timestamp 18001
transform 1 0 54556 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_587
timestamp 18001
transform 1 0 55108 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_589
timestamp 1636986456
transform 1 0 55292 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_601
timestamp 1636986456
transform 1 0 56396 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_613
timestamp 1636986456
transform 1 0 57500 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_3
timestamp 1636986456
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_15
timestamp 1636986456
transform 1 0 2484 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_27
timestamp 1636986456
transform 1 0 3588 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_39
timestamp 1636986456
transform 1 0 4692 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_63_51
timestamp 18001
transform 1 0 5796 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_55
timestamp 18001
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_57
timestamp 1636986456
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_69
timestamp 1636986456
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_81
timestamp 1636986456
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_93
timestamp 1636986456
transform 1 0 9660 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_105
timestamp 18001
transform 1 0 10764 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_111
timestamp 18001
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_113
timestamp 1636986456
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_125
timestamp 1636986456
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_137
timestamp 1636986456
transform 1 0 13708 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_149
timestamp 1636986456
transform 1 0 14812 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_161
timestamp 18001
transform 1 0 15916 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_167
timestamp 18001
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_169
timestamp 1636986456
transform 1 0 16652 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_181
timestamp 1636986456
transform 1 0 17756 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_193
timestamp 1636986456
transform 1 0 18860 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_205
timestamp 1636986456
transform 1 0 19964 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_217
timestamp 18001
transform 1 0 21068 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_223
timestamp 18001
transform 1 0 21620 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_225
timestamp 1636986456
transform 1 0 21804 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_237
timestamp 1636986456
transform 1 0 22908 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_63_249
timestamp 18001
transform 1 0 24012 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_253
timestamp 18001
transform 1 0 24380 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_265
timestamp 18001
transform 1 0 25484 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_63_273
timestamp 18001
transform 1 0 26220 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_63_285
timestamp 18001
transform 1 0 27324 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_294
timestamp 18001
transform 1 0 28152 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_321
timestamp 18001
transform 1 0 30636 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_63_341
timestamp 18001
transform 1 0 32476 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_63_375
timestamp 18001
transform 1 0 35604 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_391
timestamp 18001
transform 1 0 37076 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_63_397
timestamp 18001
transform 1 0 37628 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_63_453
timestamp 18001
transform 1 0 42780 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_494
timestamp 18001
transform 1 0 46552 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_503
timestamp 18001
transform 1 0 47380 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_511
timestamp 1636986456
transform 1 0 48116 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_523
timestamp 1636986456
transform 1 0 49220 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_535
timestamp 1636986456
transform 1 0 50324 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_547
timestamp 1636986456
transform 1 0 51428 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_559
timestamp 18001
transform 1 0 52532 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_561
timestamp 1636986456
transform 1 0 52716 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_573
timestamp 1636986456
transform 1 0 53820 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_585
timestamp 1636986456
transform 1 0 54924 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_597
timestamp 1636986456
transform 1 0 56028 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_609
timestamp 18001
transform 1 0 57132 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_615
timestamp 18001
transform 1 0 57684 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_63_617
timestamp 18001
transform 1 0 57868 0 -1 36992
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_3
timestamp 1636986456
transform 1 0 1380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_15
timestamp 1636986456
transform 1 0 2484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_27
timestamp 18001
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_29
timestamp 1636986456
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_41
timestamp 1636986456
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_53
timestamp 18001
transform 1 0 5980 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_57
timestamp 1636986456
transform 1 0 6348 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_69
timestamp 1636986456
transform 1 0 7452 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_81
timestamp 18001
transform 1 0 8556 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_85
timestamp 1636986456
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_97
timestamp 1636986456
transform 1 0 10028 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_109
timestamp 18001
transform 1 0 11132 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_113
timestamp 1636986456
transform 1 0 11500 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_125
timestamp 1636986456
transform 1 0 12604 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_137
timestamp 18001
transform 1 0 13708 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_141
timestamp 1636986456
transform 1 0 14076 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_153
timestamp 1636986456
transform 1 0 15180 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_165
timestamp 18001
transform 1 0 16284 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_169
timestamp 1636986456
transform 1 0 16652 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_181
timestamp 1636986456
transform 1 0 17756 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_193
timestamp 18001
transform 1 0 18860 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_197
timestamp 1636986456
transform 1 0 19228 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_209
timestamp 1636986456
transform 1 0 20332 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_221
timestamp 18001
transform 1 0 21436 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_64_225
timestamp 18001
transform 1 0 21804 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_233
timestamp 18001
transform 1 0 22540 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_240
timestamp 18001
transform 1 0 23184 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_64_247
timestamp 18001
transform 1 0 23828 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_251
timestamp 18001
transform 1 0 24196 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_253
timestamp 1636986456
transform 1 0 24380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_265
timestamp 1636986456
transform 1 0 25484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_277
timestamp 18001
transform 1 0 26588 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_64_287
timestamp 18001
transform 1 0 27508 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_64_295
timestamp 18001
transform 1 0 28244 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_64_303
timestamp 18001
transform 1 0 28980 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_307
timestamp 18001
transform 1 0 29348 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_309
timestamp 1636986456
transform 1 0 29532 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_321
timestamp 1636986456
transform 1 0 30636 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_333
timestamp 18001
transform 1 0 31740 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_337
timestamp 1636986456
transform 1 0 32108 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_349
timestamp 1636986456
transform 1 0 33212 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_361
timestamp 18001
transform 1 0 34316 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_365
timestamp 1636986456
transform 1 0 34684 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_377
timestamp 1636986456
transform 1 0 35788 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_389
timestamp 18001
transform 1 0 36892 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_393
timestamp 1636986456
transform 1 0 37260 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_405
timestamp 1636986456
transform 1 0 38364 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_417
timestamp 18001
transform 1 0 39468 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_421
timestamp 1636986456
transform 1 0 39836 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_433
timestamp 1636986456
transform 1 0 40940 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_445
timestamp 18001
transform 1 0 42044 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_449
timestamp 1636986456
transform 1 0 42412 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_461
timestamp 1636986456
transform 1 0 43516 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_473
timestamp 18001
transform 1 0 44620 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_477
timestamp 1636986456
transform 1 0 44988 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_489
timestamp 1636986456
transform 1 0 46092 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_501
timestamp 18001
transform 1 0 47196 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_505
timestamp 1636986456
transform 1 0 47564 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_517
timestamp 1636986456
transform 1 0 48668 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_529
timestamp 18001
transform 1 0 49772 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_533
timestamp 1636986456
transform 1 0 50140 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_545
timestamp 1636986456
transform 1 0 51244 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_557
timestamp 18001
transform 1 0 52348 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_561
timestamp 1636986456
transform 1 0 52716 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_573
timestamp 1636986456
transform 1 0 53820 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_585
timestamp 18001
transform 1 0 54924 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_589
timestamp 1636986456
transform 1 0 55292 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_601
timestamp 1636986456
transform 1 0 56396 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_613
timestamp 18001
transform 1 0 57500 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_64_617
timestamp 18001
transform 1 0 57868 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1
timestamp 18001
transform 1 0 34132 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 18001
transform -1 0 16008 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 18001
transform -1 0 37444 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 18001
transform 1 0 36340 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 18001
transform -1 0 26496 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 18001
transform -1 0 57684 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 18001
transform -1 0 41400 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 18001
transform -1 0 58604 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 18001
transform -1 0 58604 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 18001
transform -1 0 58604 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 18001
transform -1 0 58604 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp 18001
transform -1 0 14812 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp 18001
transform 1 0 22540 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold14
timestamp 18001
transform -1 0 25116 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold15
timestamp 18001
transform -1 0 23460 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold16
timestamp 18001
transform -1 0 21344 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold17
timestamp 18001
transform 1 0 22356 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold18
timestamp 18001
transform -1 0 25668 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold19
timestamp 18001
transform -1 0 14720 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold20
timestamp 18001
transform 1 0 25576 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold21
timestamp 18001
transform -1 0 23184 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold22
timestamp 18001
transform -1 0 25116 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold23
timestamp 18001
transform -1 0 17572 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold24
timestamp 18001
transform -1 0 21620 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold25
timestamp 18001
transform -1 0 17388 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold26
timestamp 18001
transform -1 0 25116 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold27
timestamp 18001
transform 1 0 24656 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold28
timestamp 18001
transform 1 0 15640 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold29
timestamp 18001
transform -1 0 27692 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold30
timestamp 18001
transform -1 0 34684 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold31
timestamp 18001
transform -1 0 20976 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold32
timestamp 18001
transform -1 0 31372 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold33
timestamp 18001
transform -1 0 27692 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold34
timestamp 18001
transform -1 0 17112 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold35
timestamp 18001
transform -1 0 35420 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold36
timestamp 18001
transform -1 0 14812 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold37
timestamp 18001
transform -1 0 29900 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold38
timestamp 18001
transform 1 0 27692 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold39
timestamp 18001
transform -1 0 32660 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold40
timestamp 18001
transform -1 0 25760 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold41
timestamp 18001
transform 1 0 25392 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold42
timestamp 18001
transform -1 0 17388 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold43
timestamp 18001
transform 1 0 17388 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold44
timestamp 18001
transform -1 0 19964 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold45
timestamp 18001
transform -1 0 19964 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold46
timestamp 18001
transform -1 0 18308 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold47
timestamp 18001
transform 1 0 24840 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold48
timestamp 18001
transform -1 0 30084 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold49
timestamp 18001
transform -1 0 27508 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold50
timestamp 18001
transform -1 0 40572 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold51
timestamp 18001
transform -1 0 21160 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold52
timestamp 18001
transform -1 0 14812 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold53
timestamp 18001
transform 1 0 17388 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold54
timestamp 18001
transform -1 0 23644 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold55
timestamp 18001
transform -1 0 49036 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold56
timestamp 18001
transform -1 0 23000 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold57
timestamp 18001
transform -1 0 27048 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold58
timestamp 18001
transform -1 0 14812 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold59
timestamp 18001
transform -1 0 46828 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold60
timestamp 18001
transform -1 0 14168 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold61
timestamp 18001
transform -1 0 15548 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold62
timestamp 18001
transform 1 0 52716 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold63
timestamp 18001
transform 1 0 28796 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold64
timestamp 18001
transform -1 0 18676 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold65
timestamp 18001
transform -1 0 40756 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold66
timestamp 18001
transform 1 0 15364 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold67
timestamp 18001
transform -1 0 20608 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold68
timestamp 18001
transform -1 0 22908 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold69
timestamp 18001
transform -1 0 39652 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold70
timestamp 18001
transform -1 0 52348 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold71
timestamp 18001
transform 1 0 20608 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold72
timestamp 18001
transform -1 0 37812 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold73
timestamp 18001
transform 1 0 37996 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold74
timestamp 18001
transform -1 0 48208 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold75
timestamp 18001
transform -1 0 20056 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold76
timestamp 18001
transform -1 0 44344 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold77
timestamp 18001
transform -1 0 31188 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold78
timestamp 18001
transform -1 0 40572 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold79
timestamp 18001
transform -1 0 52716 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold80
timestamp 18001
transform -1 0 48300 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold81
timestamp 18001
transform -1 0 14720 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold82
timestamp 18001
transform -1 0 13984 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold83
timestamp 18001
transform -1 0 53544 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold84
timestamp 18001
transform -1 0 25116 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold85
timestamp 18001
transform 1 0 44252 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold86
timestamp 18001
transform 1 0 30544 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold87
timestamp 18001
transform -1 0 50140 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold88
timestamp 18001
transform -1 0 30360 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold89
timestamp 18001
transform -1 0 54096 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold90
timestamp 18001
transform -1 0 48852 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold91
timestamp 18001
transform 1 0 47564 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold92
timestamp 18001
transform -1 0 51428 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold93
timestamp 18001
transform -1 0 48300 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold94
timestamp 18001
transform 1 0 50232 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold95
timestamp 18001
transform -1 0 39376 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold96
timestamp 18001
transform -1 0 51060 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold97
timestamp 18001
transform -1 0 50876 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold98
timestamp 18001
transform -1 0 46000 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold99
timestamp 18001
transform -1 0 52256 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold100
timestamp 18001
transform -1 0 32292 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold101
timestamp 18001
transform 1 0 47932 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold102
timestamp 18001
transform -1 0 42136 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold103
timestamp 18001
transform -1 0 52256 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold104
timestamp 18001
transform -1 0 23920 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold105
timestamp 18001
transform -1 0 31188 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold106
timestamp 18001
transform -1 0 55108 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold107
timestamp 18001
transform -1 0 27140 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold108
timestamp 18001
transform -1 0 46460 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold109
timestamp 18001
transform 1 0 55292 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold110
timestamp 18001
transform -1 0 54280 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold111
timestamp 18001
transform -1 0 48300 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold112
timestamp 18001
transform -1 0 46276 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold113
timestamp 18001
transform 1 0 31004 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold114
timestamp 18001
transform -1 0 54464 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold115
timestamp 18001
transform 1 0 22540 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold116
timestamp 18001
transform -1 0 22540 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 18001
transform 1 0 19412 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input2
timestamp 18001
transform 1 0 29164 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input3
timestamp 18001
transform 1 0 28428 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input4
timestamp 18001
transform -1 0 31004 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input5
timestamp 18001
transform -1 0 31280 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input6
timestamp 18001
transform 1 0 1380 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output7
timestamp 18001
transform 1 0 58236 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output8
timestamp 18001
transform -1 0 23184 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output9
timestamp 18001
transform -1 0 23828 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output10
timestamp 18001
transform 1 0 58236 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output11
timestamp 18001
transform 1 0 58236 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output12
timestamp 18001
transform -1 0 28980 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output13
timestamp 18001
transform 1 0 57868 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output14
timestamp 18001
transform -1 0 1748 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output15
timestamp 18001
transform 1 0 58236 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output16
timestamp 18001
transform -1 0 27508 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output17
timestamp 18001
transform 1 0 58236 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output18
timestamp 18001
transform -1 0 21068 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output19
timestamp 18001
transform -1 0 21712 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output20
timestamp 18001
transform -1 0 23644 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output21
timestamp 18001
transform -1 0 23092 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_65
timestamp 18001
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 18001
transform -1 0 58880 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_66
timestamp 18001
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 18001
transform -1 0 58880 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_67
timestamp 18001
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 18001
transform -1 0 58880 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_68
timestamp 18001
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 18001
transform -1 0 58880 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_69
timestamp 18001
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 18001
transform -1 0 58880 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_70
timestamp 18001
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 18001
transform -1 0 58880 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_71
timestamp 18001
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 18001
transform -1 0 58880 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_72
timestamp 18001
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 18001
transform -1 0 58880 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_73
timestamp 18001
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 18001
transform -1 0 58880 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_74
timestamp 18001
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 18001
transform -1 0 58880 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_75
timestamp 18001
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 18001
transform -1 0 58880 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_76
timestamp 18001
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 18001
transform -1 0 58880 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_77
timestamp 18001
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 18001
transform -1 0 58880 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_78
timestamp 18001
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 18001
transform -1 0 58880 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_79
timestamp 18001
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 18001
transform -1 0 58880 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_80
timestamp 18001
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 18001
transform -1 0 58880 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_81
timestamp 18001
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 18001
transform -1 0 58880 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_82
timestamp 18001
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 18001
transform -1 0 58880 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_83
timestamp 18001
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 18001
transform -1 0 58880 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_84
timestamp 18001
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 18001
transform -1 0 58880 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_85
timestamp 18001
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp 18001
transform -1 0 58880 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_86
timestamp 18001
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp 18001
transform -1 0 58880 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_87
timestamp 18001
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp 18001
transform -1 0 58880 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_88
timestamp 18001
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp 18001
transform -1 0 58880 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_89
timestamp 18001
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp 18001
transform -1 0 58880 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_90
timestamp 18001
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp 18001
transform -1 0 58880 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_91
timestamp 18001
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp 18001
transform -1 0 58880 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Left_92
timestamp 18001
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Right_27
timestamp 18001
transform -1 0 58880 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Left_93
timestamp 18001
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Right_28
timestamp 18001
transform -1 0 58880 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Left_94
timestamp 18001
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Right_29
timestamp 18001
transform -1 0 58880 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Left_95
timestamp 18001
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Right_30
timestamp 18001
transform -1 0 58880 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Left_96
timestamp 18001
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Right_31
timestamp 18001
transform -1 0 58880 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Left_97
timestamp 18001
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Right_32
timestamp 18001
transform -1 0 58880 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Left_98
timestamp 18001
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Right_33
timestamp 18001
transform -1 0 58880 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Left_99
timestamp 18001
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Right_34
timestamp 18001
transform -1 0 58880 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Left_100
timestamp 18001
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Right_35
timestamp 18001
transform -1 0 58880 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Left_101
timestamp 18001
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Right_36
timestamp 18001
transform -1 0 58880 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Left_102
timestamp 18001
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Right_37
timestamp 18001
transform -1 0 58880 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Left_103
timestamp 18001
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Right_38
timestamp 18001
transform -1 0 58880 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_Left_104
timestamp 18001
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_Right_39
timestamp 18001
transform -1 0 58880 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_Left_105
timestamp 18001
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_Right_40
timestamp 18001
transform -1 0 58880 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_Left_106
timestamp 18001
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_Right_41
timestamp 18001
transform -1 0 58880 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_Left_107
timestamp 18001
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_Right_42
timestamp 18001
transform -1 0 58880 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_Left_108
timestamp 18001
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_Right_43
timestamp 18001
transform -1 0 58880 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_Left_109
timestamp 18001
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_Right_44
timestamp 18001
transform -1 0 58880 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_Left_110
timestamp 18001
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_Right_45
timestamp 18001
transform -1 0 58880 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_Left_111
timestamp 18001
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_Right_46
timestamp 18001
transform -1 0 58880 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_Left_112
timestamp 18001
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_Right_47
timestamp 18001
transform -1 0 58880 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_Left_113
timestamp 18001
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_Right_48
timestamp 18001
transform -1 0 58880 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_Left_114
timestamp 18001
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_Right_49
timestamp 18001
transform -1 0 58880 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_Left_115
timestamp 18001
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_Right_50
timestamp 18001
transform -1 0 58880 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_Left_116
timestamp 18001
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_Right_51
timestamp 18001
transform -1 0 58880 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_52_Left_117
timestamp 18001
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_52_Right_52
timestamp 18001
transform -1 0 58880 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_53_Left_118
timestamp 18001
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_53_Right_53
timestamp 18001
transform -1 0 58880 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_54_Left_119
timestamp 18001
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_54_Right_54
timestamp 18001
transform -1 0 58880 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_55_Left_120
timestamp 18001
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_55_Right_55
timestamp 18001
transform -1 0 58880 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_56_Left_121
timestamp 18001
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_56_Right_56
timestamp 18001
transform -1 0 58880 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_57_Left_122
timestamp 18001
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_57_Right_57
timestamp 18001
transform -1 0 58880 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_58_Left_123
timestamp 18001
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_58_Right_58
timestamp 18001
transform -1 0 58880 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_59_Left_124
timestamp 18001
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_59_Right_59
timestamp 18001
transform -1 0 58880 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_60_Left_125
timestamp 18001
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_60_Right_60
timestamp 18001
transform -1 0 58880 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_61_Left_126
timestamp 18001
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_61_Right_61
timestamp 18001
transform -1 0 58880 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_62_Left_127
timestamp 18001
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_62_Right_62
timestamp 18001
transform -1 0 58880 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_63_Left_128
timestamp 18001
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_63_Right_63
timestamp 18001
transform -1 0 58880 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_64_Left_129
timestamp 18001
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_64_Right_64
timestamp 18001
transform -1 0 58880 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_130
timestamp 18001
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_131
timestamp 18001
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_132
timestamp 18001
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_133
timestamp 18001
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_134
timestamp 18001
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_135
timestamp 18001
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_136
timestamp 18001
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_137
timestamp 18001
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_138
timestamp 18001
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_139
timestamp 18001
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_140
timestamp 18001
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_141
timestamp 18001
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_142
timestamp 18001
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_143
timestamp 18001
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_144
timestamp 18001
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_145
timestamp 18001
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_146
timestamp 18001
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_147
timestamp 18001
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_148
timestamp 18001
transform 1 0 50048 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_149
timestamp 18001
transform 1 0 52624 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_150
timestamp 18001
transform 1 0 55200 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_151
timestamp 18001
transform 1 0 57776 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_152
timestamp 18001
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_153
timestamp 18001
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_154
timestamp 18001
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_155
timestamp 18001
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_156
timestamp 18001
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_157
timestamp 18001
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_158
timestamp 18001
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_159
timestamp 18001
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_160
timestamp 18001
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_161
timestamp 18001
transform 1 0 52624 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_162
timestamp 18001
transform 1 0 57776 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_163
timestamp 18001
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_164
timestamp 18001
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_165
timestamp 18001
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_166
timestamp 18001
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_167
timestamp 18001
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_168
timestamp 18001
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_169
timestamp 18001
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_170
timestamp 18001
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_171
timestamp 18001
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_172
timestamp 18001
transform 1 0 50048 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_173
timestamp 18001
transform 1 0 55200 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_174
timestamp 18001
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_175
timestamp 18001
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_176
timestamp 18001
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_177
timestamp 18001
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_178
timestamp 18001
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_179
timestamp 18001
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_180
timestamp 18001
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_181
timestamp 18001
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_182
timestamp 18001
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_183
timestamp 18001
transform 1 0 52624 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_184
timestamp 18001
transform 1 0 57776 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_185
timestamp 18001
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_186
timestamp 18001
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_187
timestamp 18001
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_188
timestamp 18001
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_189
timestamp 18001
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_190
timestamp 18001
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_191
timestamp 18001
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_192
timestamp 18001
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_193
timestamp 18001
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_194
timestamp 18001
transform 1 0 50048 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_195
timestamp 18001
transform 1 0 55200 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_196
timestamp 18001
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_197
timestamp 18001
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_198
timestamp 18001
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_199
timestamp 18001
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_200
timestamp 18001
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_201
timestamp 18001
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_202
timestamp 18001
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_203
timestamp 18001
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_204
timestamp 18001
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_205
timestamp 18001
transform 1 0 52624 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_206
timestamp 18001
transform 1 0 57776 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_207
timestamp 18001
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_208
timestamp 18001
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_209
timestamp 18001
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_210
timestamp 18001
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_211
timestamp 18001
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_212
timestamp 18001
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_213
timestamp 18001
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_214
timestamp 18001
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_215
timestamp 18001
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_216
timestamp 18001
transform 1 0 50048 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_217
timestamp 18001
transform 1 0 55200 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_218
timestamp 18001
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_219
timestamp 18001
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_220
timestamp 18001
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_221
timestamp 18001
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_222
timestamp 18001
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_223
timestamp 18001
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_224
timestamp 18001
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_225
timestamp 18001
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_226
timestamp 18001
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_227
timestamp 18001
transform 1 0 52624 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_228
timestamp 18001
transform 1 0 57776 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_229
timestamp 18001
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_230
timestamp 18001
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_231
timestamp 18001
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_232
timestamp 18001
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_233
timestamp 18001
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_234
timestamp 18001
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_235
timestamp 18001
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_236
timestamp 18001
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_237
timestamp 18001
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_238
timestamp 18001
transform 1 0 50048 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_239
timestamp 18001
transform 1 0 55200 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_240
timestamp 18001
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_241
timestamp 18001
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_242
timestamp 18001
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_243
timestamp 18001
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_244
timestamp 18001
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_245
timestamp 18001
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_246
timestamp 18001
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_247
timestamp 18001
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_248
timestamp 18001
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_249
timestamp 18001
transform 1 0 52624 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_250
timestamp 18001
transform 1 0 57776 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_251
timestamp 18001
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_252
timestamp 18001
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_253
timestamp 18001
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_254
timestamp 18001
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_255
timestamp 18001
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_256
timestamp 18001
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_257
timestamp 18001
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_258
timestamp 18001
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_259
timestamp 18001
transform 1 0 44896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_260
timestamp 18001
transform 1 0 50048 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_261
timestamp 18001
transform 1 0 55200 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_262
timestamp 18001
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_263
timestamp 18001
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_264
timestamp 18001
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_265
timestamp 18001
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_266
timestamp 18001
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_267
timestamp 18001
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_268
timestamp 18001
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_269
timestamp 18001
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_270
timestamp 18001
transform 1 0 47472 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_271
timestamp 18001
transform 1 0 52624 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_272
timestamp 18001
transform 1 0 57776 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_273
timestamp 18001
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_274
timestamp 18001
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_275
timestamp 18001
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_276
timestamp 18001
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_277
timestamp 18001
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_278
timestamp 18001
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_279
timestamp 18001
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_280
timestamp 18001
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_281
timestamp 18001
transform 1 0 44896 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_282
timestamp 18001
transform 1 0 50048 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_283
timestamp 18001
transform 1 0 55200 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_284
timestamp 18001
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_285
timestamp 18001
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_286
timestamp 18001
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_287
timestamp 18001
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_288
timestamp 18001
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_289
timestamp 18001
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_290
timestamp 18001
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_291
timestamp 18001
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_292
timestamp 18001
transform 1 0 47472 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_293
timestamp 18001
transform 1 0 52624 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_294
timestamp 18001
transform 1 0 57776 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_295
timestamp 18001
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_296
timestamp 18001
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_297
timestamp 18001
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_298
timestamp 18001
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_299
timestamp 18001
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_300
timestamp 18001
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_301
timestamp 18001
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_302
timestamp 18001
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_303
timestamp 18001
transform 1 0 44896 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_304
timestamp 18001
transform 1 0 50048 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_305
timestamp 18001
transform 1 0 55200 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_306
timestamp 18001
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_307
timestamp 18001
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_308
timestamp 18001
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_309
timestamp 18001
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_310
timestamp 18001
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_311
timestamp 18001
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_312
timestamp 18001
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_313
timestamp 18001
transform 1 0 42320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_314
timestamp 18001
transform 1 0 47472 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_315
timestamp 18001
transform 1 0 52624 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_316
timestamp 18001
transform 1 0 57776 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_317
timestamp 18001
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_318
timestamp 18001
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_319
timestamp 18001
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_320
timestamp 18001
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_321
timestamp 18001
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_322
timestamp 18001
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_323
timestamp 18001
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_324
timestamp 18001
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_325
timestamp 18001
transform 1 0 44896 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_326
timestamp 18001
transform 1 0 50048 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_327
timestamp 18001
transform 1 0 55200 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_328
timestamp 18001
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_329
timestamp 18001
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_330
timestamp 18001
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_331
timestamp 18001
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_332
timestamp 18001
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_333
timestamp 18001
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_334
timestamp 18001
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_335
timestamp 18001
transform 1 0 42320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_336
timestamp 18001
transform 1 0 47472 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_337
timestamp 18001
transform 1 0 52624 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_338
timestamp 18001
transform 1 0 57776 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_339
timestamp 18001
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_340
timestamp 18001
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_341
timestamp 18001
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_342
timestamp 18001
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_343
timestamp 18001
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_344
timestamp 18001
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_345
timestamp 18001
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_346
timestamp 18001
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_347
timestamp 18001
transform 1 0 44896 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_348
timestamp 18001
transform 1 0 50048 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_349
timestamp 18001
transform 1 0 55200 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_350
timestamp 18001
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_351
timestamp 18001
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_352
timestamp 18001
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_353
timestamp 18001
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_354
timestamp 18001
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_355
timestamp 18001
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_356
timestamp 18001
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_357
timestamp 18001
transform 1 0 42320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_358
timestamp 18001
transform 1 0 47472 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_359
timestamp 18001
transform 1 0 52624 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_360
timestamp 18001
transform 1 0 57776 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_361
timestamp 18001
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_362
timestamp 18001
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_363
timestamp 18001
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_364
timestamp 18001
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_365
timestamp 18001
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_366
timestamp 18001
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_367
timestamp 18001
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_368
timestamp 18001
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_369
timestamp 18001
transform 1 0 44896 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_370
timestamp 18001
transform 1 0 50048 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_371
timestamp 18001
transform 1 0 55200 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_372
timestamp 18001
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_373
timestamp 18001
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_374
timestamp 18001
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_375
timestamp 18001
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_376
timestamp 18001
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_377
timestamp 18001
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_378
timestamp 18001
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_379
timestamp 18001
transform 1 0 42320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_380
timestamp 18001
transform 1 0 47472 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_381
timestamp 18001
transform 1 0 52624 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_382
timestamp 18001
transform 1 0 57776 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_383
timestamp 18001
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_384
timestamp 18001
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_385
timestamp 18001
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_386
timestamp 18001
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_387
timestamp 18001
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_388
timestamp 18001
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_389
timestamp 18001
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_390
timestamp 18001
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_391
timestamp 18001
transform 1 0 44896 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_392
timestamp 18001
transform 1 0 50048 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_393
timestamp 18001
transform 1 0 55200 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_394
timestamp 18001
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_395
timestamp 18001
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_396
timestamp 18001
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_397
timestamp 18001
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_398
timestamp 18001
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_399
timestamp 18001
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_400
timestamp 18001
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_401
timestamp 18001
transform 1 0 42320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_402
timestamp 18001
transform 1 0 47472 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_403
timestamp 18001
transform 1 0 52624 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_404
timestamp 18001
transform 1 0 57776 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_405
timestamp 18001
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_406
timestamp 18001
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_407
timestamp 18001
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_408
timestamp 18001
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_409
timestamp 18001
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_410
timestamp 18001
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_411
timestamp 18001
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_412
timestamp 18001
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_413
timestamp 18001
transform 1 0 44896 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_414
timestamp 18001
transform 1 0 50048 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_415
timestamp 18001
transform 1 0 55200 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_416
timestamp 18001
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_417
timestamp 18001
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_418
timestamp 18001
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_419
timestamp 18001
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_420
timestamp 18001
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_421
timestamp 18001
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_422
timestamp 18001
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_423
timestamp 18001
transform 1 0 42320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_424
timestamp 18001
transform 1 0 47472 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_425
timestamp 18001
transform 1 0 52624 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_426
timestamp 18001
transform 1 0 57776 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_427
timestamp 18001
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_428
timestamp 18001
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_429
timestamp 18001
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_430
timestamp 18001
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_431
timestamp 18001
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_432
timestamp 18001
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_433
timestamp 18001
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_434
timestamp 18001
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_435
timestamp 18001
transform 1 0 44896 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_436
timestamp 18001
transform 1 0 50048 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_437
timestamp 18001
transform 1 0 55200 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_438
timestamp 18001
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_439
timestamp 18001
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_440
timestamp 18001
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_441
timestamp 18001
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_442
timestamp 18001
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_443
timestamp 18001
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_444
timestamp 18001
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_445
timestamp 18001
transform 1 0 42320 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_446
timestamp 18001
transform 1 0 47472 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_447
timestamp 18001
transform 1 0 52624 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_448
timestamp 18001
transform 1 0 57776 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_449
timestamp 18001
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_450
timestamp 18001
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_451
timestamp 18001
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_452
timestamp 18001
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_453
timestamp 18001
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_454
timestamp 18001
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_455
timestamp 18001
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_456
timestamp 18001
transform 1 0 39744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_457
timestamp 18001
transform 1 0 44896 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_458
timestamp 18001
transform 1 0 50048 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_459
timestamp 18001
transform 1 0 55200 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_460
timestamp 18001
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_461
timestamp 18001
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_462
timestamp 18001
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_463
timestamp 18001
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_464
timestamp 18001
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_465
timestamp 18001
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_466
timestamp 18001
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_467
timestamp 18001
transform 1 0 42320 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_468
timestamp 18001
transform 1 0 47472 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_469
timestamp 18001
transform 1 0 52624 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_470
timestamp 18001
transform 1 0 57776 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_471
timestamp 18001
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_472
timestamp 18001
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_473
timestamp 18001
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_474
timestamp 18001
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_475
timestamp 18001
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_476
timestamp 18001
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_477
timestamp 18001
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_478
timestamp 18001
transform 1 0 39744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_479
timestamp 18001
transform 1 0 44896 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_480
timestamp 18001
transform 1 0 50048 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_481
timestamp 18001
transform 1 0 55200 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_482
timestamp 18001
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_483
timestamp 18001
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_484
timestamp 18001
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_485
timestamp 18001
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_486
timestamp 18001
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_487
timestamp 18001
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_488
timestamp 18001
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_489
timestamp 18001
transform 1 0 42320 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_490
timestamp 18001
transform 1 0 47472 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_491
timestamp 18001
transform 1 0 52624 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_492
timestamp 18001
transform 1 0 57776 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_493
timestamp 18001
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_494
timestamp 18001
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_495
timestamp 18001
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_496
timestamp 18001
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_497
timestamp 18001
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_498
timestamp 18001
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_499
timestamp 18001
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_500
timestamp 18001
transform 1 0 39744 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_501
timestamp 18001
transform 1 0 44896 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_502
timestamp 18001
transform 1 0 50048 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_503
timestamp 18001
transform 1 0 55200 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_504
timestamp 18001
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_505
timestamp 18001
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_506
timestamp 18001
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_507
timestamp 18001
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_508
timestamp 18001
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_509
timestamp 18001
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_510
timestamp 18001
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_511
timestamp 18001
transform 1 0 42320 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_512
timestamp 18001
transform 1 0 47472 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_513
timestamp 18001
transform 1 0 52624 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_514
timestamp 18001
transform 1 0 57776 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_515
timestamp 18001
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_516
timestamp 18001
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_517
timestamp 18001
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_518
timestamp 18001
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_519
timestamp 18001
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_520
timestamp 18001
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_521
timestamp 18001
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_522
timestamp 18001
transform 1 0 39744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_523
timestamp 18001
transform 1 0 44896 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_524
timestamp 18001
transform 1 0 50048 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_525
timestamp 18001
transform 1 0 55200 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_526
timestamp 18001
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_527
timestamp 18001
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_528
timestamp 18001
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_529
timestamp 18001
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_530
timestamp 18001
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_531
timestamp 18001
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_532
timestamp 18001
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_533
timestamp 18001
transform 1 0 42320 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_534
timestamp 18001
transform 1 0 47472 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_535
timestamp 18001
transform 1 0 52624 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_536
timestamp 18001
transform 1 0 57776 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_537
timestamp 18001
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_538
timestamp 18001
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_539
timestamp 18001
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_540
timestamp 18001
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_541
timestamp 18001
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_542
timestamp 18001
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_543
timestamp 18001
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_544
timestamp 18001
transform 1 0 39744 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_545
timestamp 18001
transform 1 0 44896 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_546
timestamp 18001
transform 1 0 50048 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_547
timestamp 18001
transform 1 0 55200 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_548
timestamp 18001
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_549
timestamp 18001
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_550
timestamp 18001
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_551
timestamp 18001
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_552
timestamp 18001
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_553
timestamp 18001
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_554
timestamp 18001
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_555
timestamp 18001
transform 1 0 42320 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_556
timestamp 18001
transform 1 0 47472 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_557
timestamp 18001
transform 1 0 52624 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_558
timestamp 18001
transform 1 0 57776 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_559
timestamp 18001
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_560
timestamp 18001
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_561
timestamp 18001
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_562
timestamp 18001
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_563
timestamp 18001
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_564
timestamp 18001
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_565
timestamp 18001
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_566
timestamp 18001
transform 1 0 39744 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_567
timestamp 18001
transform 1 0 44896 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_568
timestamp 18001
transform 1 0 50048 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_569
timestamp 18001
transform 1 0 55200 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_570
timestamp 18001
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_571
timestamp 18001
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_572
timestamp 18001
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_573
timestamp 18001
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_574
timestamp 18001
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_575
timestamp 18001
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_576
timestamp 18001
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_577
timestamp 18001
transform 1 0 42320 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_578
timestamp 18001
transform 1 0 47472 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_579
timestamp 18001
transform 1 0 52624 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_580
timestamp 18001
transform 1 0 57776 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_581
timestamp 18001
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_582
timestamp 18001
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_583
timestamp 18001
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_584
timestamp 18001
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_585
timestamp 18001
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_586
timestamp 18001
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_587
timestamp 18001
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_588
timestamp 18001
transform 1 0 39744 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_589
timestamp 18001
transform 1 0 44896 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_590
timestamp 18001
transform 1 0 50048 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_591
timestamp 18001
transform 1 0 55200 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_592
timestamp 18001
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_593
timestamp 18001
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_594
timestamp 18001
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_595
timestamp 18001
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_596
timestamp 18001
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_597
timestamp 18001
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_598
timestamp 18001
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_599
timestamp 18001
transform 1 0 42320 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_600
timestamp 18001
transform 1 0 47472 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_601
timestamp 18001
transform 1 0 52624 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_602
timestamp 18001
transform 1 0 57776 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_603
timestamp 18001
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_604
timestamp 18001
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_605
timestamp 18001
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_606
timestamp 18001
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_607
timestamp 18001
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_608
timestamp 18001
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_609
timestamp 18001
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_610
timestamp 18001
transform 1 0 39744 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_611
timestamp 18001
transform 1 0 44896 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_612
timestamp 18001
transform 1 0 50048 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_613
timestamp 18001
transform 1 0 55200 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_614
timestamp 18001
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_615
timestamp 18001
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_616
timestamp 18001
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_617
timestamp 18001
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_618
timestamp 18001
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_619
timestamp 18001
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_620
timestamp 18001
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_621
timestamp 18001
transform 1 0 42320 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_622
timestamp 18001
transform 1 0 47472 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_623
timestamp 18001
transform 1 0 52624 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_624
timestamp 18001
transform 1 0 57776 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_625
timestamp 18001
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_626
timestamp 18001
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_627
timestamp 18001
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_628
timestamp 18001
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_629
timestamp 18001
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_630
timestamp 18001
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_631
timestamp 18001
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_632
timestamp 18001
transform 1 0 39744 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_633
timestamp 18001
transform 1 0 44896 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_634
timestamp 18001
transform 1 0 50048 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_635
timestamp 18001
transform 1 0 55200 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_636
timestamp 18001
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_637
timestamp 18001
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_638
timestamp 18001
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_639
timestamp 18001
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_640
timestamp 18001
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_641
timestamp 18001
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_642
timestamp 18001
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_643
timestamp 18001
transform 1 0 42320 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_644
timestamp 18001
transform 1 0 47472 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_645
timestamp 18001
transform 1 0 52624 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_646
timestamp 18001
transform 1 0 57776 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_647
timestamp 18001
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_648
timestamp 18001
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_649
timestamp 18001
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_650
timestamp 18001
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_651
timestamp 18001
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_652
timestamp 18001
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_653
timestamp 18001
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_654
timestamp 18001
transform 1 0 39744 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_655
timestamp 18001
transform 1 0 44896 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_656
timestamp 18001
transform 1 0 50048 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_657
timestamp 18001
transform 1 0 55200 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_658
timestamp 18001
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_659
timestamp 18001
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_660
timestamp 18001
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_661
timestamp 18001
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_662
timestamp 18001
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_663
timestamp 18001
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_664
timestamp 18001
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_665
timestamp 18001
transform 1 0 42320 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_666
timestamp 18001
transform 1 0 47472 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_667
timestamp 18001
transform 1 0 52624 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_668
timestamp 18001
transform 1 0 57776 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_669
timestamp 18001
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_670
timestamp 18001
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_671
timestamp 18001
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_672
timestamp 18001
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_673
timestamp 18001
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_674
timestamp 18001
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_675
timestamp 18001
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_676
timestamp 18001
transform 1 0 39744 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_677
timestamp 18001
transform 1 0 44896 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_678
timestamp 18001
transform 1 0 50048 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_679
timestamp 18001
transform 1 0 55200 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_680
timestamp 18001
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_681
timestamp 18001
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_682
timestamp 18001
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_683
timestamp 18001
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_684
timestamp 18001
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_685
timestamp 18001
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_686
timestamp 18001
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_687
timestamp 18001
transform 1 0 42320 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_688
timestamp 18001
transform 1 0 47472 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_689
timestamp 18001
transform 1 0 52624 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_690
timestamp 18001
transform 1 0 57776 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_691
timestamp 18001
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_692
timestamp 18001
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_693
timestamp 18001
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_694
timestamp 18001
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_695
timestamp 18001
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_696
timestamp 18001
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_697
timestamp 18001
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_698
timestamp 18001
transform 1 0 39744 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_699
timestamp 18001
transform 1 0 44896 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_700
timestamp 18001
transform 1 0 50048 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_701
timestamp 18001
transform 1 0 55200 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_702
timestamp 18001
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_703
timestamp 18001
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_704
timestamp 18001
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_705
timestamp 18001
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_706
timestamp 18001
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_707
timestamp 18001
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_708
timestamp 18001
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_709
timestamp 18001
transform 1 0 42320 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_710
timestamp 18001
transform 1 0 47472 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_711
timestamp 18001
transform 1 0 52624 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_712
timestamp 18001
transform 1 0 57776 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_713
timestamp 18001
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_714
timestamp 18001
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_715
timestamp 18001
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_716
timestamp 18001
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_717
timestamp 18001
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_718
timestamp 18001
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_719
timestamp 18001
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_720
timestamp 18001
transform 1 0 39744 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_721
timestamp 18001
transform 1 0 44896 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_722
timestamp 18001
transform 1 0 50048 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_723
timestamp 18001
transform 1 0 55200 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_724
timestamp 18001
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_725
timestamp 18001
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_726
timestamp 18001
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_727
timestamp 18001
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_728
timestamp 18001
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_729
timestamp 18001
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_730
timestamp 18001
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_731
timestamp 18001
transform 1 0 42320 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_732
timestamp 18001
transform 1 0 47472 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_733
timestamp 18001
transform 1 0 52624 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_734
timestamp 18001
transform 1 0 57776 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_735
timestamp 18001
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_736
timestamp 18001
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_737
timestamp 18001
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_738
timestamp 18001
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_739
timestamp 18001
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_740
timestamp 18001
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_741
timestamp 18001
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_742
timestamp 18001
transform 1 0 39744 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_743
timestamp 18001
transform 1 0 44896 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_744
timestamp 18001
transform 1 0 50048 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_745
timestamp 18001
transform 1 0 55200 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_746
timestamp 18001
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_747
timestamp 18001
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_748
timestamp 18001
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_749
timestamp 18001
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_750
timestamp 18001
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_751
timestamp 18001
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_752
timestamp 18001
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_753
timestamp 18001
transform 1 0 42320 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_754
timestamp 18001
transform 1 0 47472 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_755
timestamp 18001
transform 1 0 52624 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_756
timestamp 18001
transform 1 0 57776 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_757
timestamp 18001
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_758
timestamp 18001
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_759
timestamp 18001
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_760
timestamp 18001
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_761
timestamp 18001
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_762
timestamp 18001
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_763
timestamp 18001
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_764
timestamp 18001
transform 1 0 39744 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_765
timestamp 18001
transform 1 0 44896 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_766
timestamp 18001
transform 1 0 50048 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_767
timestamp 18001
transform 1 0 55200 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_768
timestamp 18001
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_769
timestamp 18001
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_770
timestamp 18001
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_771
timestamp 18001
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_772
timestamp 18001
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_773
timestamp 18001
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_774
timestamp 18001
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_775
timestamp 18001
transform 1 0 42320 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_776
timestamp 18001
transform 1 0 47472 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_777
timestamp 18001
transform 1 0 52624 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_778
timestamp 18001
transform 1 0 57776 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_779
timestamp 18001
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_780
timestamp 18001
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_781
timestamp 18001
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_782
timestamp 18001
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_783
timestamp 18001
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_784
timestamp 18001
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_785
timestamp 18001
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_786
timestamp 18001
transform 1 0 39744 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_787
timestamp 18001
transform 1 0 44896 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_788
timestamp 18001
transform 1 0 50048 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_789
timestamp 18001
transform 1 0 55200 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_790
timestamp 18001
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_791
timestamp 18001
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_792
timestamp 18001
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_793
timestamp 18001
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_794
timestamp 18001
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_795
timestamp 18001
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_796
timestamp 18001
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_797
timestamp 18001
transform 1 0 42320 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_798
timestamp 18001
transform 1 0 47472 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_799
timestamp 18001
transform 1 0 52624 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_800
timestamp 18001
transform 1 0 57776 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_801
timestamp 18001
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_802
timestamp 18001
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_803
timestamp 18001
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_804
timestamp 18001
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_805
timestamp 18001
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_806
timestamp 18001
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_807
timestamp 18001
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_808
timestamp 18001
transform 1 0 39744 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_809
timestamp 18001
transform 1 0 44896 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_810
timestamp 18001
transform 1 0 50048 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_811
timestamp 18001
transform 1 0 55200 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_812
timestamp 18001
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_813
timestamp 18001
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_814
timestamp 18001
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_815
timestamp 18001
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_816
timestamp 18001
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_817
timestamp 18001
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_818
timestamp 18001
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_819
timestamp 18001
transform 1 0 42320 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_820
timestamp 18001
transform 1 0 47472 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_821
timestamp 18001
transform 1 0 52624 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_822
timestamp 18001
transform 1 0 57776 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_823
timestamp 18001
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_824
timestamp 18001
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_825
timestamp 18001
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_826
timestamp 18001
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_827
timestamp 18001
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_828
timestamp 18001
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_829
timestamp 18001
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_830
timestamp 18001
transform 1 0 39744 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_831
timestamp 18001
transform 1 0 44896 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_832
timestamp 18001
transform 1 0 50048 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_833
timestamp 18001
transform 1 0 55200 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_834
timestamp 18001
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_835
timestamp 18001
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_836
timestamp 18001
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_837
timestamp 18001
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_838
timestamp 18001
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_839
timestamp 18001
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_840
timestamp 18001
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_841
timestamp 18001
transform 1 0 42320 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_842
timestamp 18001
transform 1 0 47472 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_843
timestamp 18001
transform 1 0 52624 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_844
timestamp 18001
transform 1 0 57776 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_845
timestamp 18001
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_846
timestamp 18001
transform 1 0 6256 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_847
timestamp 18001
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_848
timestamp 18001
transform 1 0 11408 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_849
timestamp 18001
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_850
timestamp 18001
transform 1 0 16560 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_851
timestamp 18001
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_852
timestamp 18001
transform 1 0 21712 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_853
timestamp 18001
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_854
timestamp 18001
transform 1 0 26864 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_855
timestamp 18001
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_856
timestamp 18001
transform 1 0 32016 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_857
timestamp 18001
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_858
timestamp 18001
transform 1 0 37168 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_859
timestamp 18001
transform 1 0 39744 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_860
timestamp 18001
transform 1 0 42320 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_861
timestamp 18001
transform 1 0 44896 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_862
timestamp 18001
transform 1 0 47472 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_863
timestamp 18001
transform 1 0 50048 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_864
timestamp 18001
transform 1 0 52624 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_865
timestamp 18001
transform 1 0 55200 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_866
timestamp 18001
transform 1 0 57776 0 1 36992
box -38 -48 130 592
<< labels >>
flabel metal3 s 59200 8168 60000 8288 0 FreeSans 480 0 0 0 clk
port 0 nsew signal input
flabel metal2 s 19338 0 19394 800 0 FreeSans 224 90 0 0 en
port 1 nsew signal input
flabel metal2 s 18 0 74 800 0 FreeSans 224 90 0 0 gpio_in[0]
port 2 nsew signal input
flabel metal2 s 662 0 718 800 0 FreeSans 224 90 0 0 gpio_in[10]
port 3 nsew signal input
flabel metal2 s 1306 0 1362 800 0 FreeSans 224 90 0 0 gpio_in[11]
port 4 nsew signal input
flabel metal2 s 1950 0 2006 800 0 FreeSans 224 90 0 0 gpio_in[12]
port 5 nsew signal input
flabel metal2 s 2594 0 2650 800 0 FreeSans 224 90 0 0 gpio_in[13]
port 6 nsew signal input
flabel metal2 s 3238 0 3294 800 0 FreeSans 224 90 0 0 gpio_in[14]
port 7 nsew signal input
flabel metal2 s 3882 0 3938 800 0 FreeSans 224 90 0 0 gpio_in[15]
port 8 nsew signal input
flabel metal2 s 4526 0 4582 800 0 FreeSans 224 90 0 0 gpio_in[16]
port 9 nsew signal input
flabel metal2 s 5170 0 5226 800 0 FreeSans 224 90 0 0 gpio_in[17]
port 10 nsew signal input
flabel metal2 s 5814 0 5870 800 0 FreeSans 224 90 0 0 gpio_in[18]
port 11 nsew signal input
flabel metal2 s 6458 0 6514 800 0 FreeSans 224 90 0 0 gpio_in[19]
port 12 nsew signal input
flabel metal2 s 7102 0 7158 800 0 FreeSans 224 90 0 0 gpio_in[1]
port 13 nsew signal input
flabel metal2 s 7746 0 7802 800 0 FreeSans 224 90 0 0 gpio_in[20]
port 14 nsew signal input
flabel metal2 s 8390 0 8446 800 0 FreeSans 224 90 0 0 gpio_in[21]
port 15 nsew signal input
flabel metal2 s 9034 0 9090 800 0 FreeSans 224 90 0 0 gpio_in[22]
port 16 nsew signal input
flabel metal2 s 9678 0 9734 800 0 FreeSans 224 90 0 0 gpio_in[23]
port 17 nsew signal input
flabel metal2 s 10322 0 10378 800 0 FreeSans 224 90 0 0 gpio_in[24]
port 18 nsew signal input
flabel metal2 s 10966 0 11022 800 0 FreeSans 224 90 0 0 gpio_in[25]
port 19 nsew signal input
flabel metal2 s 11610 0 11666 800 0 FreeSans 224 90 0 0 gpio_in[26]
port 20 nsew signal input
flabel metal2 s 12254 0 12310 800 0 FreeSans 224 90 0 0 gpio_in[27]
port 21 nsew signal input
flabel metal2 s 12898 0 12954 800 0 FreeSans 224 90 0 0 gpio_in[28]
port 22 nsew signal input
flabel metal2 s 13542 0 13598 800 0 FreeSans 224 90 0 0 gpio_in[29]
port 23 nsew signal input
flabel metal2 s 14186 0 14242 800 0 FreeSans 224 90 0 0 gpio_in[2]
port 24 nsew signal input
flabel metal2 s 29642 0 29698 800 0 FreeSans 224 90 0 0 gpio_in[30]
port 25 nsew signal input
flabel metal2 s 28998 0 29054 800 0 FreeSans 224 90 0 0 gpio_in[31]
port 26 nsew signal input
flabel metal2 s 30286 0 30342 800 0 FreeSans 224 90 0 0 gpio_in[32]
port 27 nsew signal input
flabel metal2 s 30930 0 30986 800 0 FreeSans 224 90 0 0 gpio_in[33]
port 28 nsew signal input
flabel metal2 s 14830 0 14886 800 0 FreeSans 224 90 0 0 gpio_in[3]
port 29 nsew signal input
flabel metal2 s 15474 0 15530 800 0 FreeSans 224 90 0 0 gpio_in[4]
port 30 nsew signal input
flabel metal2 s 16118 0 16174 800 0 FreeSans 224 90 0 0 gpio_in[5]
port 31 nsew signal input
flabel metal2 s 16762 0 16818 800 0 FreeSans 224 90 0 0 gpio_in[6]
port 32 nsew signal input
flabel metal2 s 17406 0 17462 800 0 FreeSans 224 90 0 0 gpio_in[7]
port 33 nsew signal input
flabel metal2 s 18050 0 18106 800 0 FreeSans 224 90 0 0 gpio_in[8]
port 34 nsew signal input
flabel metal2 s 18694 0 18750 800 0 FreeSans 224 90 0 0 gpio_in[9]
port 35 nsew signal input
flabel metal2 s 45098 0 45154 800 0 FreeSans 224 90 0 0 gpio_oeb[0]
port 36 nsew signal output
flabel metal2 s 43810 0 43866 800 0 FreeSans 224 90 0 0 gpio_oeb[10]
port 37 nsew signal output
flabel metal2 s 43166 0 43222 800 0 FreeSans 224 90 0 0 gpio_oeb[11]
port 38 nsew signal output
flabel metal2 s 38658 0 38714 800 0 FreeSans 224 90 0 0 gpio_oeb[12]
port 39 nsew signal output
flabel metal2 s 40590 0 40646 800 0 FreeSans 224 90 0 0 gpio_oeb[13]
port 40 nsew signal output
flabel metal2 s 47674 39200 47730 40000 0 FreeSans 224 90 0 0 gpio_oeb[14]
port 41 nsew signal output
flabel metal2 s 24490 39200 24546 40000 0 FreeSans 224 90 0 0 gpio_oeb[15]
port 42 nsew signal output
flabel metal2 s 34794 39200 34850 40000 0 FreeSans 224 90 0 0 gpio_oeb[16]
port 43 nsew signal output
flabel metal2 s 47030 39200 47086 40000 0 FreeSans 224 90 0 0 gpio_oeb[17]
port 44 nsew signal output
flabel metal2 s 32218 39200 32274 40000 0 FreeSans 224 90 0 0 gpio_oeb[18]
port 45 nsew signal output
flabel metal2 s 40590 39200 40646 40000 0 FreeSans 224 90 0 0 gpio_oeb[19]
port 46 nsew signal output
flabel metal2 s 41234 0 41290 800 0 FreeSans 224 90 0 0 gpio_oeb[1]
port 47 nsew signal output
flabel metal2 s 36726 39200 36782 40000 0 FreeSans 224 90 0 0 gpio_oeb[20]
port 48 nsew signal output
flabel metal2 s 28998 39200 29054 40000 0 FreeSans 224 90 0 0 gpio_oeb[21]
port 49 nsew signal output
flabel metal2 s 27710 39200 27766 40000 0 FreeSans 224 90 0 0 gpio_oeb[22]
port 50 nsew signal output
flabel metal2 s 25134 39200 25190 40000 0 FreeSans 224 90 0 0 gpio_oeb[23]
port 51 nsew signal output
flabel metal2 s 41234 39200 41290 40000 0 FreeSans 224 90 0 0 gpio_oeb[24]
port 52 nsew signal output
flabel metal2 s 38658 39200 38714 40000 0 FreeSans 224 90 0 0 gpio_oeb[25]
port 53 nsew signal output
flabel metal2 s 35438 39200 35494 40000 0 FreeSans 224 90 0 0 gpio_oeb[26]
port 54 nsew signal output
flabel metal2 s 38014 39200 38070 40000 0 FreeSans 224 90 0 0 gpio_oeb[27]
port 55 nsew signal output
flabel metal2 s 41878 39200 41934 40000 0 FreeSans 224 90 0 0 gpio_oeb[28]
port 56 nsew signal output
flabel metal2 s 27066 39200 27122 40000 0 FreeSans 224 90 0 0 gpio_oeb[29]
port 57 nsew signal output
flabel metal2 s 37370 0 37426 800 0 FreeSans 224 90 0 0 gpio_oeb[2]
port 58 nsew signal output
flabel metal2 s 36726 0 36782 800 0 FreeSans 224 90 0 0 gpio_oeb[30]
port 59 nsew signal output
flabel metal2 s 39302 0 39358 800 0 FreeSans 224 90 0 0 gpio_oeb[31]
port 60 nsew signal output
flabel metal2 s 39946 0 40002 800 0 FreeSans 224 90 0 0 gpio_oeb[32]
port 61 nsew signal output
flabel metal2 s 35438 0 35494 800 0 FreeSans 224 90 0 0 gpio_oeb[33]
port 62 nsew signal output
flabel metal2 s 41878 0 41934 800 0 FreeSans 224 90 0 0 gpio_oeb[3]
port 63 nsew signal output
flabel metal2 s 42522 0 42578 800 0 FreeSans 224 90 0 0 gpio_oeb[4]
port 64 nsew signal output
flabel metal2 s 44454 0 44510 800 0 FreeSans 224 90 0 0 gpio_oeb[5]
port 65 nsew signal output
flabel metal2 s 38014 0 38070 800 0 FreeSans 224 90 0 0 gpio_oeb[6]
port 66 nsew signal output
flabel metal2 s 36082 0 36138 800 0 FreeSans 224 90 0 0 gpio_oeb[7]
port 67 nsew signal output
flabel metal2 s 34794 0 34850 800 0 FreeSans 224 90 0 0 gpio_oeb[8]
port 68 nsew signal output
flabel metal2 s 34150 0 34206 800 0 FreeSans 224 90 0 0 gpio_oeb[9]
port 69 nsew signal output
flabel metal2 s 42522 39200 42578 40000 0 FreeSans 224 90 0 0 gpio_out[0]
port 70 nsew signal output
flabel metal2 s 43166 39200 43222 40000 0 FreeSans 224 90 0 0 gpio_out[10]
port 71 nsew signal output
flabel metal2 s 33506 39200 33562 40000 0 FreeSans 224 90 0 0 gpio_out[11]
port 72 nsew signal output
flabel metal2 s 30930 39200 30986 40000 0 FreeSans 224 90 0 0 gpio_out[12]
port 73 nsew signal output
flabel metal2 s 30286 39200 30342 40000 0 FreeSans 224 90 0 0 gpio_out[13]
port 74 nsew signal output
flabel metal3 s 59200 19728 60000 19848 0 FreeSans 480 0 0 0 gpio_out[14]
port 75 nsew signal output
flabel metal2 s 22558 39200 22614 40000 0 FreeSans 224 90 0 0 gpio_out[15]
port 76 nsew signal output
flabel metal2 s 23202 39200 23258 40000 0 FreeSans 224 90 0 0 gpio_out[16]
port 77 nsew signal output
flabel metal3 s 59200 25848 60000 25968 0 FreeSans 480 0 0 0 gpio_out[17]
port 78 nsew signal output
flabel metal3 s 59200 22448 60000 22568 0 FreeSans 480 0 0 0 gpio_out[18]
port 79 nsew signal output
flabel metal2 s 28354 39200 28410 40000 0 FreeSans 224 90 0 0 gpio_out[19]
port 80 nsew signal output
flabel metal2 s 43810 39200 43866 40000 0 FreeSans 224 90 0 0 gpio_out[1]
port 81 nsew signal output
flabel metal3 s 59200 19048 60000 19168 0 FreeSans 480 0 0 0 gpio_out[20]
port 82 nsew signal output
flabel metal3 s 0 19728 800 19848 0 FreeSans 480 0 0 0 gpio_out[21]
port 83 nsew signal output
flabel metal3 s 59200 23128 60000 23248 0 FreeSans 480 0 0 0 gpio_out[22]
port 84 nsew signal output
flabel metal2 s 39302 39200 39358 40000 0 FreeSans 224 90 0 0 gpio_out[23]
port 85 nsew signal output
flabel metal2 s 26422 39200 26478 40000 0 FreeSans 224 90 0 0 gpio_out[24]
port 86 nsew signal output
flabel metal3 s 59200 13608 60000 13728 0 FreeSans 480 0 0 0 gpio_out[25]
port 87 nsew signal output
flabel metal2 s 20626 0 20682 800 0 FreeSans 224 90 0 0 gpio_out[26]
port 88 nsew signal output
flabel metal2 s 21270 0 21326 800 0 FreeSans 224 90 0 0 gpio_out[27]
port 89 nsew signal output
flabel metal2 s 23202 0 23258 800 0 FreeSans 224 90 0 0 gpio_out[28]
port 90 nsew signal output
flabel metal2 s 22558 0 22614 800 0 FreeSans 224 90 0 0 gpio_out[29]
port 91 nsew signal output
flabel metal2 s 44454 39200 44510 40000 0 FreeSans 224 90 0 0 gpio_out[2]
port 92 nsew signal output
flabel metal2 s 29642 39200 29698 40000 0 FreeSans 224 90 0 0 gpio_out[30]
port 93 nsew signal output
flabel metal2 s 45098 39200 45154 40000 0 FreeSans 224 90 0 0 gpio_out[31]
port 94 nsew signal output
flabel metal2 s 25778 39200 25834 40000 0 FreeSans 224 90 0 0 gpio_out[32]
port 95 nsew signal output
flabel metal2 s 45742 39200 45798 40000 0 FreeSans 224 90 0 0 gpio_out[33]
port 96 nsew signal output
flabel metal2 s 36082 39200 36138 40000 0 FreeSans 224 90 0 0 gpio_out[3]
port 97 nsew signal output
flabel metal2 s 39946 39200 40002 40000 0 FreeSans 224 90 0 0 gpio_out[4]
port 98 nsew signal output
flabel metal2 s 32862 39200 32918 40000 0 FreeSans 224 90 0 0 gpio_out[5]
port 99 nsew signal output
flabel metal2 s 34150 39200 34206 40000 0 FreeSans 224 90 0 0 gpio_out[6]
port 100 nsew signal output
flabel metal2 s 31574 39200 31630 40000 0 FreeSans 224 90 0 0 gpio_out[7]
port 101 nsew signal output
flabel metal2 s 46386 39200 46442 40000 0 FreeSans 224 90 0 0 gpio_out[8]
port 102 nsew signal output
flabel metal2 s 37370 39200 37426 40000 0 FreeSans 224 90 0 0 gpio_out[9]
port 103 nsew signal output
flabel metal3 s 0 14288 800 14408 0 FreeSans 480 0 0 0 nrst
port 104 nsew signal input
flabel metal4 s 4208 2128 4528 37584 0 FreeSans 1920 90 0 0 vccd1
port 105 nsew power bidirectional
flabel metal4 s 34928 2128 35248 37584 0 FreeSans 1920 90 0 0 vccd1
port 105 nsew power bidirectional
flabel metal4 s 4868 2128 5188 37584 0 FreeSans 1920 90 0 0 vssd1
port 106 nsew ground bidirectional
flabel metal4 s 35588 2128 35908 37584 0 FreeSans 1920 90 0 0 vssd1
port 106 nsew ground bidirectional
rlabel metal1 29992 37536 29992 37536 0 vccd1
rlabel metal1 29992 36992 29992 36992 0 vssd1
rlabel metal1 37582 7514 37582 7514 0 _0000_
rlabel metal1 38548 9350 38548 9350 0 _0001_
rlabel metal1 25944 28458 25944 28458 0 _0002_
rlabel metal2 29394 31450 29394 31450 0 _0003_
rlabel metal1 29893 31994 29893 31994 0 _0004_
rlabel metal1 33626 34170 33626 34170 0 _0005_
rlabel metal1 30544 34170 30544 34170 0 _0006_
rlabel metal1 30176 33422 30176 33422 0 _0007_
rlabel metal1 28612 28118 28612 28118 0 _0008_
rlabel metal1 28934 29070 28934 29070 0 _0009_
rlabel metal1 32476 28730 32476 28730 0 _0010_
rlabel metal1 35236 29070 35236 29070 0 _0011_
rlabel metal2 32246 30464 32246 30464 0 _0012_
rlabel metal2 37306 30226 37306 30226 0 _0013_
rlabel metal1 38226 31926 38226 31926 0 _0014_
rlabel metal1 37582 33592 37582 33592 0 _0015_
rlabel metal2 36110 32674 36110 32674 0 _0016_
rlabel metal1 36892 9350 36892 9350 0 _0017_
rlabel metal1 39606 8058 39606 8058 0 _0018_
rlabel metal2 45494 13022 45494 13022 0 _0019_
rlabel metal2 31050 18360 31050 18360 0 _0020_
rlabel metal2 28106 22882 28106 22882 0 _0021_
rlabel metal1 40933 22202 40933 22202 0 _0022_
rlabel metal2 41354 20196 41354 20196 0 _0023_
rlabel metal2 34546 19108 34546 19108 0 _0024_
rlabel metal1 42044 13974 42044 13974 0 _0025_
rlabel metal2 30498 15198 30498 15198 0 _0026_
rlabel metal2 46322 13804 46322 13804 0 _0027_
rlabel metal2 32154 18530 32154 18530 0 _0028_
rlabel metal1 26732 22202 26732 22202 0 _0029_
rlabel metal2 44390 22814 44390 22814 0 _0030_
rlabel metal2 41722 21148 41722 21148 0 _0031_
rlabel metal2 34730 20196 34730 20196 0 _0032_
rlabel metal2 42734 14382 42734 14382 0 _0033_
rlabel metal2 32798 16354 32798 16354 0 _0034_
rlabel metal2 45954 15640 45954 15640 0 _0035_
rlabel metal2 28014 18462 28014 18462 0 _0036_
rlabel metal2 22402 23715 22402 23715 0 _0037_
rlabel metal2 48898 22882 48898 22882 0 _0038_
rlabel metal1 44804 19754 44804 19754 0 _0039_
rlabel metal2 35190 21692 35190 21692 0 _0040_
rlabel metal2 44298 14484 44298 14484 0 _0041_
rlabel metal2 29670 16558 29670 16558 0 _0042_
rlabel via1 48432 14790 48432 14790 0 _0043_
rlabel metal1 26266 17850 26266 17850 0 _0044_
rlabel metal2 22218 22746 22218 22746 0 _0045_
rlabel metal2 45954 25058 45954 25058 0 _0046_
rlabel metal2 45310 18972 45310 18972 0 _0047_
rlabel metal1 37260 22406 37260 22406 0 _0048_
rlabel metal2 43838 16762 43838 16762 0 _0049_
rlabel metal2 27278 16796 27278 16796 0 _0050_
rlabel metal2 49082 13294 49082 13294 0 _0051_
rlabel metal2 22586 18972 22586 18972 0 _0052_
rlabel metal2 18630 22610 18630 22610 0 _0053_
rlabel metal1 45908 25942 45908 25942 0 _0054_
rlabel metal1 48714 18802 48714 18802 0 _0055_
rlabel metal1 36340 23086 36340 23086 0 _0056_
rlabel metal1 42872 16150 42872 16150 0 _0057_
rlabel metal1 22717 16762 22717 16762 0 _0058_
rlabel metal2 51474 13532 51474 13532 0 _0059_
rlabel metal2 21942 18972 21942 18972 0 _0060_
rlabel metal2 18538 23902 18538 23902 0 _0061_
rlabel metal2 46874 26588 46874 26588 0 _0062_
rlabel metal1 50094 18938 50094 18938 0 _0063_
rlabel metal1 35236 24786 35236 24786 0 _0064_
rlabel metal2 40342 16286 40342 16286 0 _0065_
rlabel metal1 21022 16218 21022 16218 0 _0066_
rlabel metal2 51750 14824 51750 14824 0 _0067_
rlabel metal1 19320 18190 19320 18190 0 _0068_
rlabel metal2 18262 25262 18262 25262 0 _0069_
rlabel metal1 49312 27030 49312 27030 0 _0070_
rlabel metal1 51704 18938 51704 18938 0 _0071_
rlabel metal1 36202 26452 36202 26452 0 _0072_
rlabel metal1 37674 15130 37674 15130 0 _0073_
rlabel metal1 18124 17102 18124 17102 0 _0074_
rlabel metal2 53314 15232 53314 15232 0 _0075_
rlabel metal2 17618 18972 17618 18972 0 _0076_
rlabel metal1 18807 25466 18807 25466 0 _0077_
rlabel metal1 50600 27098 50600 27098 0 _0078_
rlabel metal2 53682 19754 53682 19754 0 _0079_
rlabel metal1 34822 26554 34822 26554 0 _0080_
rlabel metal1 35466 15538 35466 15538 0 _0081_
rlabel metal1 17756 16626 17756 16626 0 _0082_
rlabel metal1 56488 15062 56488 15062 0 _0083_
rlabel metal2 18814 20842 18814 20842 0 _0084_
rlabel metal2 22402 24990 22402 24990 0 _0085_
rlabel metal1 52762 26554 52762 26554 0 _0086_
rlabel metal2 55614 19992 55614 19992 0 _0087_
rlabel metal2 32798 27268 32798 27268 0 _0088_
rlabel metal1 34408 16014 34408 16014 0 _0089_
rlabel metal2 18170 15198 18170 15198 0 _0090_
rlabel metal2 56626 15844 56626 15844 0 _0091_
rlabel metal1 19044 20842 19044 20842 0 _0092_
rlabel metal2 22034 25432 22034 25432 0 _0093_
rlabel metal1 52072 25194 52072 25194 0 _0094_
rlabel metal1 57316 20570 57316 20570 0 _0095_
rlabel metal2 30958 27268 30958 27268 0 _0096_
rlabel metal2 33810 17374 33810 17374 0 _0097_
rlabel metal2 20746 14892 20746 14892 0 _0098_
rlabel metal2 56258 17374 56258 17374 0 _0099_
rlabel metal2 22218 20570 22218 20570 0 _0100_
rlabel metal1 23966 26554 23966 26554 0 _0101_
rlabel metal1 56028 25466 56028 25466 0 _0102_
rlabel metal1 55844 21658 55844 21658 0 _0103_
rlabel metal1 32292 25330 32292 25330 0 _0104_
rlabel metal2 36018 18020 36018 18020 0 _0105_
rlabel metal2 21758 14892 21758 14892 0 _0106_
rlabel metal2 54418 17374 54418 17374 0 _0107_
rlabel metal2 23690 20672 23690 20672 0 _0108_
rlabel metal1 25208 26554 25208 26554 0 _0109_
rlabel metal1 56212 24378 56212 24378 0 _0110_
rlabel metal1 52808 21590 52808 21590 0 _0111_
rlabel metal2 31418 24412 31418 24412 0 _0112_
rlabel metal2 41538 17884 41538 17884 0 _0113_
rlabel metal2 22126 14654 22126 14654 0 _0114_
rlabel metal2 52762 17816 52762 17816 0 _0115_
rlabel metal1 27048 21454 27048 21454 0 _0116_
rlabel metal1 27692 25874 27692 25874 0 _0117_
rlabel metal2 54326 23834 54326 23834 0 _0118_
rlabel metal1 50968 21114 50968 21114 0 _0119_
rlabel metal1 32200 23086 32200 23086 0 _0120_
rlabel metal1 38640 18326 38640 18326 0 _0121_
rlabel metal2 26266 14892 26266 14892 0 _0122_
rlabel metal2 50646 17442 50646 17442 0 _0123_
rlabel metal2 29946 20638 29946 20638 0 _0124_
rlabel metal1 28612 25942 28612 25942 0 _0125_
rlabel metal2 50738 23902 50738 23902 0 _0126_
rlabel metal2 47518 21284 47518 21284 0 _0127_
rlabel metal2 32154 22236 32154 22236 0 _0128_
rlabel metal1 37674 19278 37674 19278 0 _0129_
rlabel metal2 25622 13464 25622 13464 0 _0130_
rlabel metal1 47196 17306 47196 17306 0 _0131_
rlabel metal1 29633 21114 29633 21114 0 _0132_
rlabel metal1 27922 24378 27922 24378 0 _0133_
rlabel metal1 53728 22746 53728 22746 0 _0134_
rlabel metal2 45034 21284 45034 21284 0 _0135_
rlabel metal2 31602 21148 31602 21148 0 _0136_
rlabel metal1 38364 20570 38364 20570 0 _0137_
rlabel metal1 25484 12750 25484 12750 0 _0138_
rlabel metal2 25898 10404 25898 10404 0 _0139_
rlabel metal2 36662 6052 36662 6052 0 _0140_
rlabel metal2 37674 29342 37674 29342 0 _0141_
rlabel metal1 36800 28186 36800 28186 0 _0142_
rlabel metal1 39882 27608 39882 27608 0 _0143_
rlabel metal1 43010 30158 43010 30158 0 _0144_
rlabel metal1 46828 29274 46828 29274 0 _0145_
rlabel metal1 46588 27642 46588 27642 0 _0146_
rlabel metal1 25753 6970 25753 6970 0 _0147_
rlabel metal1 25714 8058 25714 8058 0 _0148_
rlabel metal1 28060 5270 28060 5270 0 _0149_
rlabel metal1 27554 5780 27554 5780 0 _0150_
rlabel metal1 29716 7242 29716 7242 0 _0151_
rlabel metal1 32384 6970 32384 6970 0 _0152_
rlabel metal1 30682 5338 30682 5338 0 _0153_
rlabel metal2 33350 5474 33350 5474 0 _0154_
rlabel metal1 40112 9962 40112 9962 0 _0155_
rlabel metal1 23920 33626 23920 33626 0 _0156_
rlabel metal1 25300 35258 25300 35258 0 _0157_
rlabel metal1 27330 35258 27330 35258 0 _0158_
rlabel metal1 27462 32538 27462 32538 0 _0159_
rlabel metal1 25576 33082 25576 33082 0 _0160_
rlabel metal1 21482 32946 21482 32946 0 _0161_
rlabel metal2 20286 33830 20286 33830 0 _0162_
rlabel metal1 17342 34374 17342 34374 0 _0163_
rlabel metal1 15318 32538 15318 32538 0 _0164_
rlabel metal2 18262 33252 18262 33252 0 _0165_
rlabel metal1 14996 31246 14996 31246 0 _0166_
rlabel metal1 17664 30634 17664 30634 0 _0167_
rlabel metal1 18400 30294 18400 30294 0 _0168_
rlabel metal2 20562 31484 20562 31484 0 _0169_
rlabel metal2 22402 31586 22402 31586 0 _0170_
rlabel metal1 22724 29818 22724 29818 0 _0171_
rlabel metal1 26404 30294 26404 30294 0 _0172_
rlabel metal1 26680 30770 26680 30770 0 _0173_
rlabel metal1 42642 12614 42642 12614 0 _0174_
rlabel metal1 29256 13498 29256 13498 0 _0175_
rlabel metal1 27002 11866 27002 11866 0 _0176_
rlabel metal1 32982 14042 32982 14042 0 _0177_
rlabel metal1 41998 12104 41998 12104 0 _0178_
rlabel metal1 35972 14042 35972 14042 0 _0179_
rlabel metal1 39008 13498 39008 13498 0 _0180_
rlabel metal1 29118 14280 29118 14280 0 _0181_
rlabel metal2 55982 23324 55982 23324 0 _0182_
rlabel metal2 20010 4318 20010 4318 0 _0183_
rlabel metal1 20424 3162 20424 3162 0 _0184_
rlabel metal1 23552 3094 23552 3094 0 _0185_
rlabel metal2 23782 3604 23782 3604 0 _0186_
rlabel metal1 57311 18734 57311 18734 0 _0187_
rlabel metal2 21942 35462 21942 35462 0 _0188_
rlabel metal2 23322 35938 23322 35938 0 _0189_
rlabel metal1 57357 25262 57357 25262 0 _0190_
rlabel metal2 57546 21794 57546 21794 0 _0191_
rlabel metal1 28888 35258 28888 35258 0 _0192_
rlabel metal1 57311 17646 57311 17646 0 _0193_
rlabel metal2 16146 19142 16146 19142 0 _0194_
rlabel metal1 18400 31790 18400 31790 0 _0195_
rlabel metal1 16560 31926 16560 31926 0 _0196_
rlabel metal1 20286 31212 20286 31212 0 _0197_
rlabel metal1 18906 30702 18906 30702 0 _0198_
rlabel metal1 21758 31178 21758 31178 0 _0199_
rlabel metal2 22034 31110 22034 31110 0 _0200_
rlabel metal1 25898 31858 25898 31858 0 _0201_
rlabel metal1 25208 31178 25208 31178 0 _0202_
rlabel metal2 32614 9860 32614 9860 0 _0203_
rlabel metal1 32890 10778 32890 10778 0 _0204_
rlabel metal1 35068 11730 35068 11730 0 _0205_
rlabel metal2 27922 10914 27922 10914 0 _0206_
rlabel metal1 32016 10030 32016 10030 0 _0207_
rlabel metal1 32614 9350 32614 9350 0 _0208_
rlabel metal1 28290 11084 28290 11084 0 _0209_
rlabel metal1 31188 10234 31188 10234 0 _0210_
rlabel metal2 34730 9962 34730 9962 0 _0211_
rlabel metal1 36294 10574 36294 10574 0 _0212_
rlabel metal2 34454 10812 34454 10812 0 _0213_
rlabel metal1 36202 10608 36202 10608 0 _0214_
rlabel metal2 38594 10676 38594 10676 0 _0215_
rlabel metal1 35512 11662 35512 11662 0 _0216_
rlabel metal1 32154 11152 32154 11152 0 _0217_
rlabel metal2 39422 11968 39422 11968 0 _0218_
rlabel metal2 35926 10268 35926 10268 0 _0219_
rlabel metal1 39330 11696 39330 11696 0 _0220_
rlabel metal1 32384 12954 32384 12954 0 _0221_
rlabel metal2 37766 13668 37766 13668 0 _0222_
rlabel metal1 33350 11798 33350 11798 0 _0223_
rlabel metal2 34914 11169 34914 11169 0 _0224_
rlabel metal1 37122 11662 37122 11662 0 _0225_
rlabel metal1 38502 11084 38502 11084 0 _0226_
rlabel metal1 39238 12784 39238 12784 0 _0227_
rlabel metal1 37720 13430 37720 13430 0 _0228_
rlabel metal1 34454 10098 34454 10098 0 _0229_
rlabel metal1 35604 13906 35604 13906 0 _0230_
rlabel metal1 39698 13294 39698 13294 0 _0231_
rlabel metal1 39514 12104 39514 12104 0 _0232_
rlabel metal1 39422 11288 39422 11288 0 _0233_
rlabel metal1 35972 11866 35972 11866 0 _0234_
rlabel metal1 34960 11866 34960 11866 0 _0235_
rlabel metal1 35006 12172 35006 12172 0 _0236_
rlabel metal1 35098 10778 35098 10778 0 _0237_
rlabel metal2 35466 11730 35466 11730 0 _0238_
rlabel metal2 42918 12461 42918 12461 0 _0239_
rlabel via2 29762 11747 29762 11747 0 _0240_
rlabel metal1 29118 11628 29118 11628 0 _0241_
rlabel metal1 30084 12614 30084 12614 0 _0242_
rlabel metal2 31510 11900 31510 11900 0 _0243_
rlabel metal1 31832 13158 31832 13158 0 _0244_
rlabel metal1 32706 11254 32706 11254 0 _0245_
rlabel metal2 33718 11084 33718 11084 0 _0246_
rlabel metal1 29578 12342 29578 12342 0 _0247_
rlabel metal2 31786 11492 31786 11492 0 _0248_
rlabel metal2 30498 11322 30498 11322 0 _0249_
rlabel metal1 30452 11322 30452 11322 0 _0250_
rlabel metal1 30774 12104 30774 12104 0 _0251_
rlabel metal1 30038 12410 30038 12410 0 _0252_
rlabel metal2 31142 13124 31142 13124 0 _0253_
rlabel metal1 29854 13260 29854 13260 0 _0254_
rlabel metal1 33028 12750 33028 12750 0 _0255_
rlabel metal1 29716 10234 29716 10234 0 _0256_
rlabel metal1 29302 10676 29302 10676 0 _0257_
rlabel metal1 29946 10778 29946 10778 0 _0258_
rlabel metal1 29026 12750 29026 12750 0 _0259_
rlabel metal1 29256 12682 29256 12682 0 _0260_
rlabel metal1 29302 12410 29302 12410 0 _0261_
rlabel metal1 28152 12818 28152 12818 0 _0262_
rlabel metal1 27876 11118 27876 11118 0 _0263_
rlabel metal1 28428 11322 28428 11322 0 _0264_
rlabel metal2 32614 11900 32614 11900 0 _0265_
rlabel metal1 33120 12614 33120 12614 0 _0266_
rlabel metal2 33534 13396 33534 13396 0 _0267_
rlabel metal1 39514 11220 39514 11220 0 _0268_
rlabel metal1 39330 10778 39330 10778 0 _0269_
rlabel metal2 39146 11492 39146 11492 0 _0270_
rlabel metal1 39698 11730 39698 11730 0 _0271_
rlabel metal1 40296 11866 40296 11866 0 _0272_
rlabel metal1 40388 11594 40388 11594 0 _0273_
rlabel metal2 38594 13464 38594 13464 0 _0274_
rlabel metal1 38916 10710 38916 10710 0 _0275_
rlabel metal1 37076 13158 37076 13158 0 _0276_
rlabel metal2 36478 13600 36478 13600 0 _0277_
rlabel metal2 36294 13702 36294 13702 0 _0278_
rlabel metal2 39238 13056 39238 13056 0 _0279_
rlabel metal1 30406 14382 30406 14382 0 _0280_
rlabel metal1 42182 25398 42182 25398 0 _0281_
rlabel via1 38683 25262 38683 25262 0 _0282_
rlabel metal1 39514 24174 39514 24174 0 _0283_
rlabel metal2 39606 22780 39606 22780 0 _0284_
rlabel metal2 40066 26112 40066 26112 0 _0285_
rlabel metal1 38272 23086 38272 23086 0 _0286_
rlabel via2 39790 22389 39790 22389 0 _0287_
rlabel via1 42926 26010 42926 26010 0 _0288_
rlabel metal1 42734 23086 42734 23086 0 _0289_
rlabel metal1 42458 24174 42458 24174 0 _0290_
rlabel metal2 39974 23477 39974 23477 0 _0291_
rlabel metal1 39928 24786 39928 24786 0 _0292_
rlabel metal1 32614 25704 32614 25704 0 _0293_
rlabel metal1 44850 23222 44850 23222 0 _0294_
rlabel metal2 56718 23341 56718 23341 0 _0295_
rlabel metal2 22954 4318 22954 4318 0 _0296_
rlabel metal2 21206 3706 21206 3706 0 _0297_
rlabel metal1 21482 3026 21482 3026 0 _0298_
rlabel metal2 23506 3910 23506 3910 0 _0299_
rlabel metal1 22770 3162 22770 3162 0 _0300_
rlabel metal1 23000 2482 23000 2482 0 _0301_
rlabel metal3 45494 21964 45494 21964 0 _0302_
rlabel metal1 33994 19822 33994 19822 0 _0303_
rlabel metal1 40250 21046 40250 21046 0 _0304_
rlabel via1 40160 18258 40160 18258 0 _0305_
rlabel metal1 43378 25772 43378 25772 0 _0306_
rlabel metal2 39514 17000 39514 17000 0 _0307_
rlabel metal2 38870 25007 38870 25007 0 _0308_
rlabel metal1 48346 16116 48346 16116 0 _0309_
rlabel metal2 39882 19023 39882 19023 0 _0310_
rlabel metal2 40894 19652 40894 19652 0 _0311_
rlabel metal1 38778 22746 38778 22746 0 _0312_
rlabel metal2 33994 23494 33994 23494 0 _0313_
rlabel metal2 40894 17255 40894 17255 0 _0314_
rlabel metal2 41170 16966 41170 16966 0 _0315_
rlabel metal1 37858 18326 37858 18326 0 _0316_
rlabel metal1 40066 18326 40066 18326 0 _0317_
rlabel metal2 38778 24344 38778 24344 0 _0318_
rlabel metal1 35420 23698 35420 23698 0 _0319_
rlabel metal1 48668 16762 48668 16762 0 _0320_
rlabel metal1 49542 16422 49542 16422 0 _0321_
rlabel metal2 49726 17476 49726 17476 0 _0322_
rlabel metal2 49542 17578 49542 17578 0 _0323_
rlabel metal1 49036 15946 49036 15946 0 _0324_
rlabel metal1 47610 16558 47610 16558 0 _0325_
rlabel metal2 48392 16762 48392 16762 0 _0326_
rlabel metal2 56626 18598 56626 18598 0 _0327_
rlabel metal1 28014 19380 28014 19380 0 _0328_
rlabel metal2 25438 20230 25438 20230 0 _0329_
rlabel metal1 25208 18938 25208 18938 0 _0330_
rlabel metal1 28750 19482 28750 19482 0 _0331_
rlabel metal1 26358 20026 26358 20026 0 _0332_
rlabel metal1 26726 19924 26726 19924 0 _0333_
rlabel metal3 34822 20468 34822 20468 0 _0334_
rlabel metal2 30406 19312 30406 19312 0 _0335_
rlabel metal1 26450 18938 26450 18938 0 _0336_
rlabel metal1 26772 19686 26772 19686 0 _0337_
rlabel metal2 25070 24004 25070 24004 0 _0338_
rlabel metal2 25530 24378 25530 24378 0 _0339_
rlabel metal1 25806 24378 25806 24378 0 _0340_
rlabel metal1 25944 23698 25944 23698 0 _0341_
rlabel metal1 26128 23698 26128 23698 0 _0342_
rlabel metal1 25392 23834 25392 23834 0 _0343_
rlabel metal2 26082 24956 26082 24956 0 _0344_
rlabel metal1 28704 24310 28704 24310 0 _0345_
rlabel metal2 25438 24412 25438 24412 0 _0346_
rlabel metal1 25162 35496 25162 35496 0 _0347_
rlabel metal1 49542 23290 49542 23290 0 _0348_
rlabel metal2 50370 24718 50370 24718 0 _0349_
rlabel metal2 50278 25092 50278 25092 0 _0350_
rlabel metal1 50048 24922 50048 24922 0 _0351_
rlabel via2 41998 25347 41998 25347 0 _0352_
rlabel metal1 48162 25432 48162 25432 0 _0353_
rlabel metal2 50186 25636 50186 25636 0 _0354_
rlabel metal2 45310 23970 45310 23970 0 _0355_
rlabel metal1 49174 24276 49174 24276 0 _0356_
rlabel metal2 48806 24106 48806 24106 0 _0357_
rlabel metal1 49266 24174 49266 24174 0 _0358_
rlabel metal1 49496 24378 49496 24378 0 _0359_
rlabel metal2 56902 25823 56902 25823 0 _0360_
rlabel metal1 44206 21046 44206 21046 0 _0361_
rlabel metal1 48162 20026 48162 20026 0 _0362_
rlabel metal1 48990 20026 48990 20026 0 _0363_
rlabel metal1 47426 20808 47426 20808 0 _0364_
rlabel metal2 49358 20502 49358 20502 0 _0365_
rlabel metal1 49036 20230 49036 20230 0 _0366_
rlabel metal1 49358 20366 49358 20366 0 _0367_
rlabel metal2 47610 20740 47610 20740 0 _0368_
rlabel metal1 49082 20400 49082 20400 0 _0369_
rlabel metal2 56902 20995 56902 20995 0 _0370_
rlabel metal1 29348 35258 29348 35258 0 _0371_
rlabel metal1 35650 23732 35650 23732 0 _0372_
rlabel metal2 35006 24072 35006 24072 0 _0373_
rlabel metal1 37536 24786 37536 24786 0 _0374_
rlabel metal2 37490 24990 37490 24990 0 _0375_
rlabel metal1 37674 24684 37674 24684 0 _0376_
rlabel metal1 38134 24786 38134 24786 0 _0377_
rlabel metal2 34546 24480 34546 24480 0 _0378_
rlabel metal1 33304 23834 33304 23834 0 _0379_
rlabel metal1 34362 24276 34362 24276 0 _0380_
rlabel metal1 34040 20026 34040 20026 0 _0381_
rlabel metal1 34638 21658 34638 21658 0 _0382_
rlabel via2 34086 24395 34086 24395 0 _0383_
rlabel metal1 43056 17306 43056 17306 0 _0384_
rlabel metal1 40986 17748 40986 17748 0 _0385_
rlabel metal1 39790 16422 39790 16422 0 _0386_
rlabel metal2 40710 17986 40710 17986 0 _0387_
rlabel metal1 39560 16762 39560 16762 0 _0388_
rlabel metal2 40618 17476 40618 17476 0 _0389_
rlabel metal2 40066 18054 40066 18054 0 _0390_
rlabel metal2 39882 16898 39882 16898 0 _0391_
rlabel metal1 40526 17578 40526 17578 0 _0392_
rlabel metal2 41170 17561 41170 17561 0 _0393_
rlabel metal2 26818 16252 26818 16252 0 _0394_
rlabel metal2 24426 16762 24426 16762 0 _0395_
rlabel metal2 24978 16694 24978 16694 0 _0396_
rlabel metal1 25254 16422 25254 16422 0 _0397_
rlabel metal1 26956 16558 26956 16558 0 _0398_
rlabel metal1 25806 16694 25806 16694 0 _0399_
rlabel metal2 25898 16864 25898 16864 0 _0400_
rlabel metal1 28106 17034 28106 17034 0 _0401_
rlabel metal1 25392 17170 25392 17170 0 _0402_
rlabel metal2 16790 18020 16790 18020 0 _0403_
rlabel metal1 27692 11050 27692 11050 0 _0404_
rlabel metal1 32982 28526 32982 28526 0 _0405_
rlabel metal1 20838 33898 20838 33898 0 _0406_
rlabel metal1 42734 27982 42734 27982 0 _0407_
rlabel metal2 39698 28730 39698 28730 0 _0408_
rlabel metal1 44712 27642 44712 27642 0 _0409_
rlabel via2 43286 28509 43286 28509 0 _0410_
rlabel metal1 42044 27438 42044 27438 0 _0411_
rlabel metal1 37214 7854 37214 7854 0 _0412_
rlabel metal1 37352 8330 37352 8330 0 _0413_
rlabel metal2 32982 9622 32982 9622 0 _0414_
rlabel metal2 32062 9758 32062 9758 0 _0415_
rlabel metal1 37444 5882 37444 5882 0 _0416_
rlabel metal1 37214 8908 37214 8908 0 _0417_
rlabel metal1 28934 6154 28934 6154 0 _0418_
rlabel metal2 30406 6528 30406 6528 0 _0419_
rlabel metal1 29118 6392 29118 6392 0 _0420_
rlabel metal1 30728 6426 30728 6426 0 _0421_
rlabel metal1 35742 6732 35742 6732 0 _0422_
rlabel metal2 33994 6494 33994 6494 0 _0423_
rlabel metal2 34454 7344 34454 7344 0 _0424_
rlabel metal2 35374 7004 35374 7004 0 _0425_
rlabel metal1 27324 6630 27324 6630 0 _0426_
rlabel metal1 27186 6766 27186 6766 0 _0427_
rlabel metal2 27370 7344 27370 7344 0 _0428_
rlabel metal1 35558 7310 35558 7310 0 _0429_
rlabel metal1 36248 6766 36248 6766 0 _0430_
rlabel metal1 36524 7990 36524 7990 0 _0431_
rlabel metal2 36754 7174 36754 7174 0 _0432_
rlabel metal1 36662 8500 36662 8500 0 _0433_
rlabel metal2 36570 7174 36570 7174 0 _0434_
rlabel metal1 30728 2414 30728 2414 0 _0435_
rlabel metal1 16330 11118 16330 11118 0 _0436_
rlabel metal2 20194 11152 20194 11152 0 _0437_
rlabel metal1 17112 11186 17112 11186 0 _0438_
rlabel metal1 15870 14790 15870 14790 0 _0439_
rlabel metal2 15870 5984 15870 5984 0 _0440_
rlabel metal1 20516 6426 20516 6426 0 _0441_
rlabel metal2 21206 8194 21206 8194 0 _0442_
rlabel metal1 16054 6392 16054 6392 0 _0443_
rlabel metal1 20148 10030 20148 10030 0 _0444_
rlabel metal2 17250 9554 17250 9554 0 _0445_
rlabel metal1 15778 6426 15778 6426 0 _0446_
rlabel metal2 16698 7684 16698 7684 0 _0447_
rlabel metal2 17802 5236 17802 5236 0 _0448_
rlabel metal1 16652 5338 16652 5338 0 _0449_
rlabel metal1 14076 5678 14076 5678 0 _0450_
rlabel metal2 14306 5882 14306 5882 0 _0451_
rlabel metal2 12926 6494 12926 6494 0 _0452_
rlabel metal1 13478 5678 13478 5678 0 _0453_
rlabel metal1 17158 7990 17158 7990 0 _0454_
rlabel metal2 16146 7820 16146 7820 0 _0455_
rlabel metal1 20838 6630 20838 6630 0 _0456_
rlabel metal2 17618 7548 17618 7548 0 _0457_
rlabel metal2 18170 6256 18170 6256 0 _0458_
rlabel metal1 17848 5610 17848 5610 0 _0459_
rlabel metal2 21114 5916 21114 5916 0 _0460_
rlabel metal2 21390 7548 21390 7548 0 _0461_
rlabel metal2 21298 6426 21298 6426 0 _0462_
rlabel metal1 20700 7922 20700 7922 0 _0463_
rlabel metal2 23046 7004 23046 7004 0 _0464_
rlabel metal1 21904 8874 21904 8874 0 _0465_
rlabel metal1 22586 9418 22586 9418 0 _0466_
rlabel metal2 21390 10914 21390 10914 0 _0467_
rlabel via1 22410 9894 22410 9894 0 _0468_
rlabel metal2 21666 10302 21666 10302 0 _0469_
rlabel metal1 18722 11118 18722 11118 0 _0470_
rlabel metal2 16790 9724 16790 9724 0 _0471_
rlabel metal2 18262 10948 18262 10948 0 _0472_
rlabel metal2 18078 10404 18078 10404 0 _0473_
rlabel metal1 14674 10064 14674 10064 0 _0474_
rlabel metal2 13570 10982 13570 10982 0 _0475_
rlabel metal1 16928 10778 16928 10778 0 _0476_
rlabel metal2 14858 11764 14858 11764 0 _0477_
rlabel metal2 15502 11322 15502 11322 0 _0478_
rlabel metal1 15180 12206 15180 12206 0 _0479_
rlabel metal1 19688 12410 19688 12410 0 _0480_
rlabel metal1 17710 12138 17710 12138 0 _0481_
rlabel metal1 18124 12818 18124 12818 0 _0482_
rlabel metal1 18262 12716 18262 12716 0 _0483_
rlabel metal1 16100 13158 16100 13158 0 _0484_
rlabel metal2 12374 14586 12374 14586 0 _0485_
rlabel metal1 12190 14416 12190 14416 0 _0486_
rlabel metal1 15272 13498 15272 13498 0 _0487_
rlabel metal1 24564 31246 24564 31246 0 _0488_
rlabel metal1 18998 31858 18998 31858 0 _0489_
rlabel metal2 19274 32266 19274 32266 0 _0490_
rlabel metal2 23414 31433 23414 31433 0 _0491_
rlabel metal1 24242 32878 24242 32878 0 _0492_
rlabel metal1 25346 34918 25346 34918 0 _0493_
rlabel metal1 26450 33966 26450 33966 0 _0494_
rlabel metal2 25990 33082 25990 33082 0 _0495_
rlabel metal1 23506 32878 23506 32878 0 _0496_
rlabel metal2 25806 34068 25806 34068 0 _0497_
rlabel metal2 28842 29274 28842 29274 0 _0498_
rlabel metal1 28972 29478 28972 29478 0 _0499_
rlabel metal2 30682 28832 30682 28832 0 _0500_
rlabel metal1 32476 29546 32476 29546 0 _0501_
rlabel metal1 32108 28730 32108 28730 0 _0502_
rlabel metal1 34132 32470 34132 32470 0 _0503_
rlabel metal2 32798 28968 32798 28968 0 _0504_
rlabel metal1 34684 29818 34684 29818 0 _0505_
rlabel metal1 34140 29478 34140 29478 0 _0506_
rlabel metal2 33902 32249 33902 32249 0 _0507_
rlabel metal1 33534 31790 33534 31790 0 _0508_
rlabel metal1 33856 31790 33856 31790 0 _0509_
rlabel metal2 33810 32232 33810 32232 0 _0510_
rlabel metal1 33672 32198 33672 32198 0 _0511_
rlabel metal1 32890 32878 32890 32878 0 _0512_
rlabel metal1 33856 30090 33856 30090 0 _0513_
rlabel metal1 32982 30192 32982 30192 0 _0514_
rlabel metal2 37490 29784 37490 29784 0 _0515_
rlabel metal1 37996 31790 37996 31790 0 _0516_
rlabel metal1 37628 31654 37628 31654 0 _0517_
rlabel metal1 36846 32334 36846 32334 0 _0518_
rlabel metal1 37766 33082 37766 33082 0 _0519_
rlabel metal2 36662 32946 36662 32946 0 _0520_
rlabel metal1 34638 32300 34638 32300 0 _0521_
rlabel metal2 36294 32572 36294 32572 0 _0522_
rlabel metal1 30222 32198 30222 32198 0 _0523_
rlabel metal2 29394 32028 29394 32028 0 _0524_
rlabel metal1 33304 32266 33304 32266 0 _0525_
rlabel metal2 32798 33422 32798 33422 0 _0526_
rlabel metal1 30130 32436 30130 32436 0 _0527_
rlabel metal1 34178 33898 34178 33898 0 _0528_
rlabel metal1 32062 33864 32062 33864 0 _0529_
rlabel metal1 31004 33354 31004 33354 0 _0530_
rlabel metal2 31142 33286 31142 33286 0 _0531_
rlabel metal1 33856 31654 33856 31654 0 _0532_
rlabel metal1 33212 33082 33212 33082 0 _0533_
rlabel metal2 36754 8636 36754 8636 0 _0534_
rlabel metal1 36938 9996 36938 9996 0 _0535_
rlabel metal1 36662 9928 36662 9928 0 _0536_
rlabel metal1 37904 7922 37904 7922 0 _0537_
rlabel metal1 32798 8602 32798 8602 0 _0538_
rlabel via2 38778 17187 38778 17187 0 _0539_
rlabel metal2 37306 16439 37306 16439 0 _0540_
rlabel metal1 37030 13294 37030 13294 0 _0541_
rlabel metal1 32522 9520 32522 9520 0 _0542_
rlabel metal1 39054 12852 39054 12852 0 _0543_
rlabel metal1 36662 14960 36662 14960 0 _0544_
rlabel metal1 35742 13498 35742 13498 0 _0545_
rlabel metal1 32154 13260 32154 13260 0 _0546_
rlabel metal1 35420 17170 35420 17170 0 _0547_
rlabel metal1 45678 13226 45678 13226 0 _0548_
rlabel metal2 30590 19108 30590 19108 0 _0549_
rlabel metal2 28382 23086 28382 23086 0 _0550_
rlabel metal1 41446 22644 41446 22644 0 _0551_
rlabel metal1 41630 19788 41630 19788 0 _0552_
rlabel metal2 36938 13770 36938 13770 0 _0553_
rlabel metal2 36938 17204 36938 17204 0 _0554_
rlabel metal1 34270 18768 34270 18768 0 _0555_
rlabel metal1 41262 14416 41262 14416 0 _0556_
rlabel metal1 30728 15470 30728 15470 0 _0557_
rlabel metal1 46460 14042 46460 14042 0 _0558_
rlabel metal1 30958 18326 30958 18326 0 _0559_
rlabel metal1 26082 22644 26082 22644 0 _0560_
rlabel metal1 44574 23052 44574 23052 0 _0561_
rlabel metal2 43102 21012 43102 21012 0 _0562_
rlabel metal1 35006 19890 35006 19890 0 _0563_
rlabel metal1 43286 14586 43286 14586 0 _0564_
rlabel metal2 31786 16524 31786 16524 0 _0565_
rlabel metal1 46552 15130 46552 15130 0 _0566_
rlabel metal2 28290 18428 28290 18428 0 _0567_
rlabel metal1 23322 23834 23322 23834 0 _0568_
rlabel metal1 48622 22644 48622 22644 0 _0569_
rlabel metal2 45218 20026 45218 20026 0 _0570_
rlabel metal1 35512 21114 35512 21114 0 _0571_
rlabel metal2 44574 14620 44574 14620 0 _0572_
rlabel metal1 30038 16762 30038 16762 0 _0573_
rlabel metal1 48622 14586 48622 14586 0 _0574_
rlabel metal1 26174 17680 26174 17680 0 _0575_
rlabel metal1 21758 23154 21758 23154 0 _0576_
rlabel metal1 46276 23834 46276 23834 0 _0577_
rlabel metal1 46230 19482 46230 19482 0 _0578_
rlabel metal1 36570 22678 36570 22678 0 _0579_
rlabel metal1 44344 16218 44344 16218 0 _0580_
rlabel metal1 27830 15878 27830 15878 0 _0581_
rlabel metal2 49174 14076 49174 14076 0 _0582_
rlabel metal1 23184 18394 23184 18394 0 _0583_
rlabel metal1 18814 22032 18814 22032 0 _0584_
rlabel metal2 48254 25840 48254 25840 0 _0585_
rlabel metal1 48898 19346 48898 19346 0 _0586_
rlabel metal1 36248 24174 36248 24174 0 _0587_
rlabel metal1 43056 15674 43056 15674 0 _0588_
rlabel metal1 23184 16218 23184 16218 0 _0589_
rlabel metal1 51750 13940 51750 13940 0 _0590_
rlabel metal1 21896 18394 21896 18394 0 _0591_
rlabel metal1 19826 23834 19826 23834 0 _0592_
rlabel metal2 48346 26452 48346 26452 0 _0593_
rlabel metal1 50462 18700 50462 18700 0 _0594_
rlabel metal1 35650 24820 35650 24820 0 _0595_
rlabel metal1 40618 15674 40618 15674 0 _0596_
rlabel metal1 21620 16082 21620 16082 0 _0597_
rlabel metal1 52302 15504 52302 15504 0 _0598_
rlabel metal2 20286 18428 20286 18428 0 _0599_
rlabel metal2 19826 25364 19826 25364 0 _0600_
rlabel metal1 49496 26554 49496 26554 0 _0601_
rlabel metal2 51842 19210 51842 19210 0 _0602_
rlabel metal2 36478 26401 36478 26401 0 _0603_
rlabel metal1 38088 14994 38088 14994 0 _0604_
rlabel metal1 19274 17170 19274 17170 0 _0605_
rlabel metal1 53774 15504 53774 15504 0 _0606_
rlabel metal1 19090 19380 19090 19380 0 _0607_
rlabel metal1 20286 25194 20286 25194 0 _0608_
rlabel metal2 50830 26758 50830 26758 0 _0609_
rlabel metal1 53912 20026 53912 20026 0 _0610_
rlabel metal1 35190 26384 35190 26384 0 _0611_
rlabel metal1 36018 16116 36018 16116 0 _0612_
rlabel metal1 18722 16592 18722 16592 0 _0613_
rlabel metal2 56258 15572 56258 15572 0 _0614_
rlabel metal1 19274 21522 19274 21522 0 _0615_
rlabel metal2 21206 25466 21206 25466 0 _0616_
rlabel metal1 52440 26010 52440 26010 0 _0617_
rlabel metal1 55292 20026 55292 20026 0 _0618_
rlabel metal1 33074 27030 33074 27030 0 _0619_
rlabel metal2 35190 16490 35190 16490 0 _0620_
rlabel metal1 19458 15436 19458 15436 0 _0621_
rlabel metal1 56948 15470 56948 15470 0 _0622_
rlabel metal1 18814 21012 18814 21012 0 _0623_
rlabel metal2 23322 25670 23322 25670 0 _0624_
rlabel metal2 51842 25466 51842 25466 0 _0625_
rlabel metal1 56442 20434 56442 20434 0 _0626_
rlabel metal1 32384 26554 32384 26554 0 _0627_
rlabel metal1 35466 17306 35466 17306 0 _0628_
rlabel metal1 19918 15130 19918 15130 0 _0629_
rlabel metal1 56764 16762 56764 16762 0 _0630_
rlabel metal1 22034 21046 22034 21046 0 _0631_
rlabel metal2 24886 25976 24886 25976 0 _0632_
rlabel metal1 55890 25262 55890 25262 0 _0633_
rlabel metal1 55522 21488 55522 21488 0 _0634_
rlabel metal2 33350 25466 33350 25466 0 _0635_
rlabel metal1 36386 17646 36386 17646 0 _0636_
rlabel metal2 22218 15300 22218 15300 0 _0637_
rlabel metal1 54326 17306 54326 17306 0 _0638_
rlabel metal2 23874 20876 23874 20876 0 _0639_
rlabel metal1 25438 26418 25438 26418 0 _0640_
rlabel metal2 56350 24378 56350 24378 0 _0641_
rlabel metal2 52486 21318 52486 21318 0 _0642_
rlabel metal1 31694 24752 31694 24752 0 _0643_
rlabel metal1 41538 18292 41538 18292 0 _0644_
rlabel metal1 23138 14586 23138 14586 0 _0645_
rlabel metal1 53176 17306 53176 17306 0 _0646_
rlabel metal1 26358 21114 26358 21114 0 _0647_
rlabel metal2 28014 26180 28014 26180 0 _0648_
rlabel metal1 54326 24140 54326 24140 0 _0649_
rlabel metal1 51106 20978 51106 20978 0 _0650_
rlabel metal2 32706 23290 32706 23290 0 _0651_
rlabel metal1 39330 18224 39330 18224 0 _0652_
rlabel metal1 25668 15130 25668 15130 0 _0653_
rlabel metal2 50922 17612 50922 17612 0 _0654_
rlabel metal1 29348 20570 29348 20570 0 _0655_
rlabel metal1 28888 25466 28888 25466 0 _0656_
rlabel metal1 50876 23290 50876 23290 0 _0657_
rlabel metal1 47886 21862 47886 21862 0 _0658_
rlabel metal1 32614 21658 32614 21658 0 _0659_
rlabel metal1 38226 19414 38226 19414 0 _0660_
rlabel metal2 25806 13260 25806 13260 0 _0661_
rlabel metal1 47886 17136 47886 17136 0 _0662_
rlabel metal2 29302 21046 29302 21046 0 _0663_
rlabel metal1 28290 24140 28290 24140 0 _0664_
rlabel metal2 53774 23052 53774 23052 0 _0665_
rlabel metal2 45310 21386 45310 21386 0 _0666_
rlabel metal1 31878 21488 31878 21488 0 _0667_
rlabel metal1 38778 20468 38778 20468 0 _0668_
rlabel metal1 26404 12342 26404 12342 0 _0669_
rlabel metal1 32200 9554 32200 9554 0 _0670_
rlabel metal1 26772 10098 26772 10098 0 _0671_
rlabel metal2 33534 31212 33534 31212 0 _0672_
rlabel metal2 34178 31025 34178 31025 0 _0673_
rlabel metal1 33212 30566 33212 30566 0 _0674_
rlabel metal1 38410 28730 38410 28730 0 _0675_
rlabel metal1 40802 29274 40802 29274 0 _0676_
rlabel metal1 43378 27506 43378 27506 0 _0677_
rlabel metal1 41170 29172 41170 29172 0 _0678_
rlabel metal2 40618 29138 40618 29138 0 _0679_
rlabel metal1 40802 29002 40802 29002 0 _0680_
rlabel metal1 41147 29546 41147 29546 0 _0681_
rlabel metal2 43930 27302 43930 27302 0 _0682_
rlabel metal2 40802 29444 40802 29444 0 _0683_
rlabel metal1 40894 29104 40894 29104 0 _0684_
rlabel metal1 40480 29138 40480 29138 0 _0685_
rlabel metal1 34187 30906 34187 30906 0 _0686_
rlabel metal1 34592 30702 34592 30702 0 _0687_
rlabel metal1 39514 17646 39514 17646 0 _0688_
rlabel metal2 43102 27846 43102 27846 0 _0689_
rlabel metal2 43654 27744 43654 27744 0 _0690_
rlabel metal1 42090 24786 42090 24786 0 _0691_
rlabel metal1 40802 25194 40802 25194 0 _0692_
rlabel metal1 42780 25670 42780 25670 0 _0693_
rlabel metal2 40986 24956 40986 24956 0 _0694_
rlabel metal1 42688 24242 42688 24242 0 _0695_
rlabel metal2 38962 27302 38962 27302 0 _0696_
rlabel metal2 40986 27710 40986 27710 0 _0697_
rlabel metal1 40388 26894 40388 26894 0 _0698_
rlabel metal1 40572 26962 40572 26962 0 _0699_
rlabel metal2 39974 27200 39974 27200 0 _0700_
rlabel metal1 43102 29818 43102 29818 0 _0701_
rlabel metal1 44712 28730 44712 28730 0 _0702_
rlabel metal2 43470 28730 43470 28730 0 _0703_
rlabel metal1 43884 28050 43884 28050 0 _0704_
rlabel metal1 38433 25330 38433 25330 0 _0705_
rlabel metal1 44252 28050 44252 28050 0 _0706_
rlabel metal1 44896 27914 44896 27914 0 _0707_
rlabel metal1 45954 28730 45954 28730 0 _0708_
rlabel metal2 43470 26146 43470 26146 0 _0709_
rlabel metal1 45724 27302 45724 27302 0 _0710_
rlabel metal2 33810 10642 33810 10642 0 _0711_
rlabel metal1 35328 9622 35328 9622 0 _0712_
rlabel metal1 25898 34646 25898 34646 0 _0713_
rlabel metal1 26496 34442 26496 34442 0 _0714_
rlabel metal1 26818 32368 26818 32368 0 _0715_
rlabel metal1 25806 32912 25806 32912 0 _0716_
rlabel metal2 22034 33728 22034 33728 0 _0717_
rlabel metal1 20286 33864 20286 33864 0 _0718_
rlabel metal1 16744 32334 16744 32334 0 _0719_
rlabel metal1 15916 31994 15916 31994 0 _0720_
rlabel metal2 18354 33422 18354 33422 0 _0721_
rlabel via2 36846 18581 36846 18581 0 clk
rlabel via2 37122 18717 37122 18717 0 clknet_0_clk
rlabel metal1 16560 12954 16560 12954 0 clknet_1_0__leaf_clk
rlabel metal1 40756 19414 40756 19414 0 clknet_1_1__leaf_clk
rlabel metal2 16698 15878 16698 15878 0 clknet_leaf_0_clk
rlabel metal1 36524 32946 36524 32946 0 clknet_leaf_10_clk
rlabel metal1 52762 26860 52762 26860 0 clknet_leaf_11_clk
rlabel metal1 55752 19890 55752 19890 0 clknet_leaf_12_clk
rlabel metal1 44252 21454 44252 21454 0 clknet_leaf_13_clk
rlabel metal1 37536 19890 37536 19890 0 clknet_leaf_14_clk
rlabel metal1 49128 18802 49128 18802 0 clknet_leaf_15_clk
rlabel metal2 53038 14688 53038 14688 0 clknet_leaf_16_clk
rlabel metal2 49818 13634 49818 13634 0 clknet_leaf_17_clk
rlabel metal2 37122 7072 37122 7072 0 clknet_leaf_18_clk
rlabel metal1 36938 14450 36938 14450 0 clknet_leaf_19_clk
rlabel metal1 21252 14382 21252 14382 0 clknet_leaf_1_clk
rlabel metal2 33534 17680 33534 17680 0 clknet_leaf_20_clk
rlabel metal1 31947 7378 31947 7378 0 clknet_leaf_21_clk
rlabel metal2 32798 5168 32798 5168 0 clknet_leaf_22_clk
rlabel metal2 22034 7038 22034 7038 0 clknet_leaf_23_clk
rlabel metal1 12098 6154 12098 6154 0 clknet_leaf_24_clk
rlabel metal2 12190 12002 12190 12002 0 clknet_leaf_25_clk
rlabel metal1 27462 22066 27462 22066 0 clknet_leaf_2_clk
rlabel metal2 19274 23392 19274 23392 0 clknet_leaf_3_clk
rlabel metal1 18538 20468 18538 20468 0 clknet_leaf_4_clk
rlabel metal1 14168 32878 14168 32878 0 clknet_leaf_5_clk
rlabel metal1 20746 32878 20746 32878 0 clknet_leaf_6_clk
rlabel metal2 32338 33150 32338 33150 0 clknet_leaf_7_clk
rlabel metal1 33626 27506 33626 27506 0 clknet_leaf_8_clk
rlabel metal1 37352 26962 37352 26962 0 clknet_leaf_9_clk
rlabel metal2 19366 1520 19366 1520 0 en
rlabel metal1 29394 2346 29394 2346 0 gpio_in[30]
rlabel metal1 28704 2482 28704 2482 0 gpio_in[31]
rlabel metal1 30912 2414 30912 2414 0 gpio_in[32]
rlabel metal1 31142 2346 31142 2346 0 gpio_in[33]
rlabel metal2 45126 1792 45126 1792 0 gpio_oeb[0]
rlabel metal2 43838 1792 43838 1792 0 gpio_oeb[10]
rlabel metal2 43194 1792 43194 1792 0 gpio_oeb[11]
rlabel metal1 38640 2822 38640 2822 0 gpio_oeb[12]
rlabel metal1 40572 2822 40572 2822 0 gpio_oeb[13]
rlabel metal1 47426 36890 47426 36890 0 gpio_oeb[14]
rlabel metal1 24748 36890 24748 36890 0 gpio_oeb[15]
rlabel metal1 34776 36890 34776 36890 0 gpio_oeb[16]
rlabel metal1 46920 36890 46920 36890 0 gpio_oeb[17]
rlabel metal1 32292 36890 32292 36890 0 gpio_oeb[18]
rlabel metal1 40572 36890 40572 36890 0 gpio_oeb[19]
rlabel metal1 41216 2822 41216 2822 0 gpio_oeb[1]
rlabel metal1 36662 36890 36662 36890 0 gpio_oeb[20]
rlabel metal1 28934 36890 28934 36890 0 gpio_oeb[21]
rlabel metal1 27692 36890 27692 36890 0 gpio_oeb[22]
rlabel metal1 25208 36890 25208 36890 0 gpio_oeb[23]
rlabel metal1 41216 36890 41216 36890 0 gpio_oeb[24]
rlabel metal1 38640 36890 38640 36890 0 gpio_oeb[25]
rlabel metal2 35466 38056 35466 38056 0 gpio_oeb[26]
rlabel metal1 37996 36890 37996 36890 0 gpio_oeb[27]
rlabel metal1 41860 36890 41860 36890 0 gpio_oeb[28]
rlabel metal1 27140 36890 27140 36890 0 gpio_oeb[29]
rlabel metal1 37444 2822 37444 2822 0 gpio_oeb[2]
rlabel metal1 36708 2822 36708 2822 0 gpio_oeb[30]
rlabel metal1 39284 2822 39284 2822 0 gpio_oeb[31]
rlabel metal1 39928 2822 39928 2822 0 gpio_oeb[32]
rlabel metal2 35466 1792 35466 1792 0 gpio_oeb[33]
rlabel metal2 41906 1792 41906 1792 0 gpio_oeb[3]
rlabel metal2 42550 1792 42550 1792 0 gpio_oeb[4]
rlabel metal2 44482 1792 44482 1792 0 gpio_oeb[5]
rlabel metal1 37996 2822 37996 2822 0 gpio_oeb[6]
rlabel metal1 36064 2822 36064 2822 0 gpio_oeb[7]
rlabel metal1 34868 2822 34868 2822 0 gpio_oeb[8]
rlabel metal1 34408 2822 34408 2822 0 gpio_oeb[9]
rlabel metal1 42596 36890 42596 36890 0 gpio_out[0]
rlabel metal1 43148 36890 43148 36890 0 gpio_out[10]
rlabel metal1 33488 36890 33488 36890 0 gpio_out[11]
rlabel metal1 30912 36890 30912 36890 0 gpio_out[12]
rlabel metal1 30222 36890 30222 36890 0 gpio_out[13]
rlabel metal2 58466 19737 58466 19737 0 gpio_out[14]
rlabel metal1 22678 37434 22678 37434 0 gpio_out[15]
rlabel metal1 23322 37434 23322 37434 0 gpio_out[16]
rlabel metal1 58190 26486 58190 26486 0 gpio_out[17]
rlabel via2 58466 22491 58466 22491 0 gpio_out[18]
rlabel metal1 28474 37434 28474 37434 0 gpio_out[19]
rlabel metal1 43792 36890 43792 36890 0 gpio_out[1]
rlabel metal1 58006 19686 58006 19686 0 gpio_out[20]
rlabel metal3 751 19788 751 19788 0 gpio_out[21]
rlabel metal2 58466 23341 58466 23341 0 gpio_out[22]
rlabel metal1 39284 36890 39284 36890 0 gpio_out[23]
rlabel metal1 26772 37434 26772 37434 0 gpio_out[24]
rlabel via2 58466 13685 58466 13685 0 gpio_out[25]
rlabel metal2 20654 1520 20654 1520 0 gpio_out[26]
rlabel metal2 21298 1520 21298 1520 0 gpio_out[27]
rlabel metal2 23230 1520 23230 1520 0 gpio_out[28]
rlabel metal2 22586 1656 22586 1656 0 gpio_out[29]
rlabel metal1 44436 36890 44436 36890 0 gpio_out[2]
rlabel metal1 29578 36890 29578 36890 0 gpio_out[30]
rlabel metal1 45080 36890 45080 36890 0 gpio_out[31]
rlabel metal1 25760 36890 25760 36890 0 gpio_out[32]
rlabel metal1 45724 36890 45724 36890 0 gpio_out[33]
rlabel metal1 36018 36890 36018 36890 0 gpio_out[3]
rlabel metal1 39928 36890 39928 36890 0 gpio_out[4]
rlabel metal1 32844 36890 32844 36890 0 gpio_out[5]
rlabel metal1 34132 36890 34132 36890 0 gpio_out[6]
rlabel metal1 31556 36890 31556 36890 0 gpio_out[7]
rlabel metal2 46414 38056 46414 38056 0 gpio_out[8]
rlabel metal1 37444 36890 37444 36890 0 gpio_out[9]
rlabel metal1 26358 7310 26358 7310 0 kp.buffertop.keycode\[0\]
rlabel metal1 26358 7718 26358 7718 0 kp.buffertop.keycode\[1\]
rlabel metal1 28796 5542 28796 5542 0 kp.buffertop.keycode\[2\]
rlabel metal1 27968 5542 27968 5542 0 kp.buffertop.keycode\[3\]
rlabel metal1 32706 8466 32706 8466 0 kp.buffertop.keycode\[4\]
rlabel metal1 32752 6630 32752 6630 0 kp.buffertop.keycode\[5\]
rlabel metal2 31786 7242 31786 7242 0 kp.buffertop.keycode\[6\]
rlabel metal2 33810 4148 33810 4148 0 kp.buffertop.keycode\[7\]
rlabel metal1 27646 7412 27646 7412 0 kp.buffertop.keycode_previous\[0\]
rlabel metal1 27186 8398 27186 8398 0 kp.buffertop.keycode_previous\[1\]
rlabel metal1 29256 6290 29256 6290 0 kp.buffertop.keycode_previous\[2\]
rlabel metal1 27508 6290 27508 6290 0 kp.buffertop.keycode_previous\[3\]
rlabel metal2 31326 7548 31326 7548 0 kp.buffertop.keycode_previous\[4\]
rlabel metal2 33902 7684 33902 7684 0 kp.buffertop.keycode_previous\[5\]
rlabel metal2 31878 6086 31878 6086 0 kp.buffertop.keycode_previous\[6\]
rlabel metal2 34546 6086 34546 6086 0 kp.buffertop.keycode_previous\[7\]
rlabel metal2 20286 13855 20286 13855 0 kp.buffertop.nrst
rlabel metal2 17342 4284 17342 4284 0 kp.clkdivtop.count\[0\]
rlabel metal1 21022 6766 21022 6766 0 kp.clkdivtop.count\[10\]
rlabel metal1 21482 8466 21482 8466 0 kp.clkdivtop.count\[11\]
rlabel metal1 21620 9146 21620 9146 0 kp.clkdivtop.count\[12\]
rlabel metal2 21390 8534 21390 8534 0 kp.clkdivtop.count\[13\]
rlabel metal1 20930 10710 20930 10710 0 kp.clkdivtop.count\[14\]
rlabel metal2 20746 10880 20746 10880 0 kp.clkdivtop.count\[15\]
rlabel metal1 17066 10608 17066 10608 0 kp.clkdivtop.count\[16\]
rlabel metal1 18676 10438 18676 10438 0 kp.clkdivtop.count\[17\]
rlabel metal2 15686 10812 15686 10812 0 kp.clkdivtop.count\[18\]
rlabel metal2 15870 10880 15870 10880 0 kp.clkdivtop.count\[19\]
rlabel metal2 16514 5423 16514 5423 0 kp.clkdivtop.count\[1\]
rlabel metal1 14260 11662 14260 11662 0 kp.clkdivtop.count\[20\]
rlabel metal1 14766 12308 14766 12308 0 kp.clkdivtop.count\[21\]
rlabel metal1 18630 12240 18630 12240 0 kp.clkdivtop.count\[22\]
rlabel metal1 21160 11662 21160 11662 0 kp.clkdivtop.count\[23\]
rlabel metal1 17986 12886 17986 12886 0 kp.clkdivtop.count\[24\]
rlabel metal1 18538 13158 18538 13158 0 kp.clkdivtop.count\[25\]
rlabel metal1 14858 14790 14858 14790 0 kp.clkdivtop.count\[26\]
rlabel metal1 13662 14450 13662 14450 0 kp.clkdivtop.count\[27\]
rlabel metal2 14766 14722 14766 14722 0 kp.clkdivtop.count\[28\]
rlabel metal2 15502 14076 15502 14076 0 kp.clkdivtop.count\[29\]
rlabel metal1 15640 5746 15640 5746 0 kp.clkdivtop.count\[2\]
rlabel metal1 14536 6426 14536 6426 0 kp.clkdivtop.count\[3\]
rlabel metal2 14030 7548 14030 7548 0 kp.clkdivtop.count\[4\]
rlabel metal1 16606 7378 16606 7378 0 kp.clkdivtop.count\[5\]
rlabel metal2 16698 8670 16698 8670 0 kp.clkdivtop.count\[6\]
rlabel metal1 20562 6834 20562 6834 0 kp.clkdivtop.count\[7\]
rlabel metal1 20424 6766 20424 6766 0 kp.clkdivtop.count\[8\]
rlabel metal1 21666 6222 21666 6222 0 kp.clkdivtop.count\[9\]
rlabel metal1 15640 4522 15640 4522 0 kp.clkdivtop.next_count\[0\]
rlabel metal1 23926 6970 23926 6970 0 kp.clkdivtop.next_count\[10\]
rlabel metal1 19642 8058 19642 8058 0 kp.clkdivtop.next_count\[11\]
rlabel metal1 23690 8398 23690 8398 0 kp.clkdivtop.next_count\[12\]
rlabel metal2 23690 9452 23690 9452 0 kp.clkdivtop.next_count\[13\]
rlabel metal1 23184 11186 23184 11186 0 kp.clkdivtop.next_count\[14\]
rlabel metal2 22862 10404 22862 10404 0 kp.clkdivtop.next_count\[15\]
rlabel metal2 16882 9826 16882 9826 0 kp.clkdivtop.next_count\[16\]
rlabel metal1 18400 10710 18400 10710 0 kp.clkdivtop.next_count\[17\]
rlabel metal2 13478 10030 13478 10030 0 kp.clkdivtop.next_count\[18\]
rlabel metal1 13984 10234 13984 10234 0 kp.clkdivtop.next_count\[19\]
rlabel metal2 16238 5406 16238 5406 0 kp.clkdivtop.next_count\[1\]
rlabel metal2 12466 11492 12466 11492 0 kp.clkdivtop.next_count\[20\]
rlabel metal1 12466 12104 12466 12104 0 kp.clkdivtop.next_count\[21\]
rlabel metal1 21344 12274 21344 12274 0 kp.clkdivtop.next_count\[22\]
rlabel metal1 19688 11798 19688 11798 0 kp.clkdivtop.next_count\[23\]
rlabel metal1 16054 13362 16054 13362 0 kp.clkdivtop.next_count\[24\]
rlabel metal1 17618 13192 17618 13192 0 kp.clkdivtop.next_count\[25\]
rlabel metal2 13294 15300 13294 15300 0 kp.clkdivtop.next_count\[26\]
rlabel metal2 12282 13804 12282 13804 0 kp.clkdivtop.next_count\[27\]
rlabel metal2 13202 14212 13202 14212 0 kp.clkdivtop.next_count\[28\]
rlabel metal1 16192 14450 16192 14450 0 kp.clkdivtop.next_count\[29\]
rlabel metal1 13478 5134 13478 5134 0 kp.clkdivtop.next_count\[2\]
rlabel metal2 13018 6052 13018 6052 0 kp.clkdivtop.next_count\[3\]
rlabel metal2 12466 7548 12466 7548 0 kp.clkdivtop.next_count\[4\]
rlabel metal1 15272 7514 15272 7514 0 kp.clkdivtop.next_count\[5\]
rlabel metal1 17802 7514 17802 7514 0 kp.clkdivtop.next_count\[6\]
rlabel metal1 18768 5882 18768 5882 0 kp.clkdivtop.next_count\[7\]
rlabel metal1 19550 5576 19550 5576 0 kp.clkdivtop.next_count\[8\]
rlabel metal2 23322 6052 23322 6052 0 kp.clkdivtop.next_count\[9\]
rlabel metal2 26726 10931 26726 10931 0 kp.controlstop.mode
rlabel metal2 57454 12988 57454 12988 0 kp.controlstop.msg_tx_ctrl
rlabel metal2 36846 13260 36846 13260 0 kp.controlstop.next_msg_tx_ctrl
rlabel metal1 37513 7310 37513 7310 0 kp.controlstop.previous_key_count\[0\]
rlabel metal1 38318 8432 38318 8432 0 kp.controlstop.previous_key_count\[1\]
rlabel metal2 36018 8636 36018 8636 0 kp.controlstop.previous_key_count\[2\]
rlabel metal1 37674 8942 37674 8942 0 kp.controlstop.previous_key_count\[3\]
rlabel metal2 40618 10370 40618 10370 0 kp.controlstop.upper
rlabel metal1 33718 4794 33718 4794 0 kp.debouncertop.keyvalid
rlabel metal2 36294 5814 36294 5814 0 kp.debouncertop.next_receive_ready
rlabel metal2 36202 5712 36202 5712 0 kp.debouncertop.receive_ready
rlabel metal2 48162 14093 48162 14093 0 kp.decodertop.data_received\[0\]
rlabel metal1 50682 20944 50682 20944 0 kp.decodertop.data_received\[100\]
rlabel metal1 33005 24378 33005 24378 0 kp.decodertop.data_received\[101\]
rlabel metal2 38778 17952 38778 17952 0 kp.decodertop.data_received\[102\]
rlabel metal2 25898 15572 25898 15572 0 kp.decodertop.data_received\[103\]
rlabel via1 50277 17170 50277 17170 0 kp.decodertop.data_received\[104\]
rlabel viali 23965 21522 23965 21522 0 kp.decodertop.data_received\[105\]
rlabel metal2 26358 25636 26358 25636 0 kp.decodertop.data_received\[106\]
rlabel metal1 50646 23188 50646 23188 0 kp.decodertop.data_received\[107\]
rlabel metal1 49358 22066 49358 22066 0 kp.decodertop.data_received\[108\]
rlabel metal1 32338 21624 32338 21624 0 kp.decodertop.data_received\[109\]
rlabel metal1 28474 10744 28474 10744 0 kp.decodertop.data_received\[10\]
rlabel metal1 39468 18938 39468 18938 0 kp.decodertop.data_received\[110\]
rlabel metal1 24748 15538 24748 15538 0 kp.decodertop.data_received\[111\]
rlabel metal1 46874 17068 46874 17068 0 kp.decodertop.data_received\[112\]
rlabel metal1 28382 20366 28382 20366 0 kp.decodertop.data_received\[113\]
rlabel metal2 30222 26486 30222 26486 0 kp.decodertop.data_received\[114\]
rlabel metal2 52210 24004 52210 24004 0 kp.decodertop.data_received\[115\]
rlabel metal1 44758 21998 44758 21998 0 kp.decodertop.data_received\[116\]
rlabel metal1 32706 22644 32706 22644 0 kp.decodertop.data_received\[117\]
rlabel metal1 38364 18258 38364 18258 0 kp.decodertop.data_received\[118\]
rlabel metal1 30314 14892 30314 14892 0 kp.decodertop.data_received\[119\]
rlabel metal2 41538 19516 41538 19516 0 kp.decodertop.data_received\[11\]
rlabel metal1 49266 17646 49266 17646 0 kp.decodertop.data_received\[120\]
rlabel metal1 27692 20774 27692 20774 0 kp.decodertop.data_received\[121\]
rlabel metal2 28382 24990 28382 24990 0 kp.decodertop.data_received\[122\]
rlabel metal2 51934 22780 51934 22780 0 kp.decodertop.data_received\[123\]
rlabel metal1 48622 21998 48622 21998 0 kp.decodertop.data_received\[124\]
rlabel metal1 33603 21114 33603 21114 0 kp.decodertop.data_received\[125\]
rlabel via1 40066 20978 40066 20978 0 kp.decodertop.data_received\[126\]
rlabel via1 24426 13906 24426 13906 0 kp.decodertop.data_received\[127\]
rlabel metal1 41561 11050 41561 11050 0 kp.decodertop.data_received\[12\]
rlabel metal1 36179 19346 36179 19346 0 kp.decodertop.data_received\[13\]
rlabel metal1 40572 13838 40572 13838 0 kp.decodertop.data_received\[14\]
rlabel metal2 32154 16388 32154 16388 0 kp.decodertop.data_received\[15\]
rlabel metal1 46782 14960 46782 14960 0 kp.decodertop.data_received\[16\]
rlabel metal1 30912 18598 30912 18598 0 kp.decodertop.data_received\[17\]
rlabel metal1 24794 22610 24794 22610 0 kp.decodertop.data_received\[18\]
rlabel metal1 48530 23800 48530 23800 0 kp.decodertop.data_received\[19\]
rlabel metal2 30314 19074 30314 19074 0 kp.decodertop.data_received\[1\]
rlabel metal2 44942 20672 44942 20672 0 kp.decodertop.data_received\[20\]
rlabel metal1 35282 20910 35282 20910 0 kp.decodertop.data_received\[21\]
rlabel metal1 40480 14382 40480 14382 0 kp.decodertop.data_received\[22\]
rlabel metal1 31004 16626 31004 16626 0 kp.decodertop.data_received\[23\]
rlabel metal2 47426 14654 47426 14654 0 kp.decodertop.data_received\[24\]
rlabel metal2 26358 19176 26358 19176 0 kp.decodertop.data_received\[25\]
rlabel metal1 23184 23290 23184 23290 0 kp.decodertop.data_received\[26\]
rlabel metal1 47472 23766 47472 23766 0 kp.decodertop.data_received\[27\]
rlabel metal2 46690 19618 46690 19618 0 kp.decodertop.data_received\[28\]
rlabel metal1 36363 21318 36363 21318 0 kp.decodertop.data_received\[29\]
rlabel metal2 27830 23647 27830 23647 0 kp.decodertop.data_received\[2\]
rlabel metal1 42780 14858 42780 14858 0 kp.decodertop.data_received\[30\]
rlabel metal2 31142 16389 31142 16389 0 kp.decodertop.data_received\[31\]
rlabel metal1 47058 14960 47058 14960 0 kp.decodertop.data_received\[32\]
rlabel metal1 24288 18190 24288 18190 0 kp.decodertop.data_received\[33\]
rlabel metal1 21206 23086 21206 23086 0 kp.decodertop.data_received\[34\]
rlabel metal2 47794 24055 47794 24055 0 kp.decodertop.data_received\[35\]
rlabel metal1 46598 20502 46598 20502 0 kp.decodertop.data_received\[36\]
rlabel metal1 36386 22610 36386 22610 0 kp.decodertop.data_received\[37\]
rlabel metal1 43562 15436 43562 15436 0 kp.decodertop.data_received\[38\]
rlabel viali 29670 16558 29670 16558 0 kp.decodertop.data_received\[39\]
rlabel metal1 37168 14858 37168 14858 0 kp.decodertop.data_received\[3\]
rlabel metal2 48990 14909 48990 14909 0 kp.decodertop.data_received\[40\]
rlabel metal1 23368 19346 23368 19346 0 kp.decodertop.data_received\[41\]
rlabel metal1 22770 24208 22770 24208 0 kp.decodertop.data_received\[42\]
rlabel viali 47518 24174 47518 24174 0 kp.decodertop.data_received\[43\]
rlabel metal1 49358 18666 49358 18666 0 kp.decodertop.data_received\[44\]
rlabel metal1 36478 24208 36478 24208 0 kp.decodertop.data_received\[45\]
rlabel metal2 40250 16320 40250 16320 0 kp.decodertop.data_received\[46\]
rlabel metal1 23230 17102 23230 17102 0 kp.decodertop.data_received\[47\]
rlabel metal2 49496 14382 49496 14382 0 kp.decodertop.data_received\[48\]
rlabel metal1 20240 18666 20240 18666 0 kp.decodertop.data_received\[49\]
rlabel metal1 42826 20434 42826 20434 0 kp.decodertop.data_received\[4\]
rlabel metal1 22264 23494 22264 23494 0 kp.decodertop.data_received\[50\]
rlabel metal1 48530 26554 48530 26554 0 kp.decodertop.data_received\[51\]
rlabel metal1 51796 19278 51796 19278 0 kp.decodertop.data_received\[52\]
rlabel metal1 36409 25466 36409 25466 0 kp.decodertop.data_received\[53\]
rlabel metal1 38410 16048 38410 16048 0 kp.decodertop.data_received\[54\]
rlabel metal2 21666 16626 21666 16626 0 kp.decodertop.data_received\[55\]
rlabel metal2 52578 15198 52578 15198 0 kp.decodertop.data_received\[56\]
rlabel metal1 19826 19414 19826 19414 0 kp.decodertop.data_received\[57\]
rlabel metal1 21068 23698 21068 23698 0 kp.decodertop.data_received\[58\]
rlabel metal2 50646 27710 50646 27710 0 kp.decodertop.data_received\[59\]
rlabel metal2 36294 19618 36294 19618 0 kp.decodertop.data_received\[5\]
rlabel metal1 52118 18666 52118 18666 0 kp.decodertop.data_received\[60\]
rlabel metal1 36984 26350 36984 26350 0 kp.decodertop.data_received\[61\]
rlabel metal1 39330 16116 39330 16116 0 kp.decodertop.data_received\[62\]
rlabel metal1 19067 17034 19067 17034 0 kp.decodertop.data_received\[63\]
rlabel metal2 51382 15776 51382 15776 0 kp.decodertop.data_received\[64\]
rlabel metal1 19458 19346 19458 19346 0 kp.decodertop.data_received\[65\]
rlabel metal1 22218 25840 22218 25840 0 kp.decodertop.data_received\[66\]
rlabel metal1 52256 27506 52256 27506 0 kp.decodertop.data_received\[67\]
rlabel metal2 54878 20060 54878 20060 0 kp.decodertop.data_received\[68\]
rlabel metal2 39054 25874 39054 25874 0 kp.decodertop.data_received\[69\]
rlabel metal1 40526 14450 40526 14450 0 kp.decodertop.data_received\[6\]
rlabel metal2 38686 16252 38686 16252 0 kp.decodertop.data_received\[70\]
rlabel metal1 19642 16048 19642 16048 0 kp.decodertop.data_received\[71\]
rlabel metal2 48070 16218 48070 16218 0 kp.decodertop.data_received\[72\]
rlabel metal2 20516 21522 20516 21522 0 kp.decodertop.data_received\[73\]
rlabel metal2 20930 25092 20930 25092 0 kp.decodertop.data_received\[74\]
rlabel metal1 50279 26316 50279 26316 0 kp.decodertop.data_received\[75\]
rlabel via1 53406 19822 53406 19822 0 kp.decodertop.data_received\[76\]
rlabel metal1 34546 27030 34546 27030 0 kp.decodertop.data_received\[77\]
rlabel metal1 37444 16082 37444 16082 0 kp.decodertop.data_received\[78\]
rlabel metal1 19734 15572 19734 15572 0 kp.decodertop.data_received\[79\]
rlabel metal1 30314 15572 30314 15572 0 kp.decodertop.data_received\[7\]
rlabel metal1 55108 15470 55108 15470 0 kp.decodertop.data_received\[80\]
rlabel metal1 19090 20978 19090 20978 0 kp.decodertop.data_received\[81\]
rlabel metal1 25162 25874 25162 25874 0 kp.decodertop.data_received\[82\]
rlabel via1 51658 25874 51658 25874 0 kp.decodertop.data_received\[83\]
rlabel via1 54602 19822 54602 19822 0 kp.decodertop.data_received\[84\]
rlabel metal1 32798 26962 32798 26962 0 kp.decodertop.data_received\[85\]
rlabel metal1 36938 17680 36938 17680 0 kp.decodertop.data_received\[86\]
rlabel metal2 19826 15164 19826 15164 0 kp.decodertop.data_received\[87\]
rlabel metal1 53724 17170 53724 17170 0 kp.decodertop.data_received\[88\]
rlabel metal2 22402 21216 22402 21216 0 kp.decodertop.data_received\[89\]
rlabel metal2 45954 12784 45954 12784 0 kp.decodertop.data_received\[8\]
rlabel metal1 24932 26350 24932 26350 0 kp.decodertop.data_received\[90\]
rlabel metal1 53240 25874 53240 25874 0 kp.decodertop.data_received\[91\]
rlabel via2 52210 20893 52210 20893 0 kp.decodertop.data_received\[92\]
rlabel metal1 33626 25228 33626 25228 0 kp.decodertop.data_received\[93\]
rlabel metal2 37122 18496 37122 18496 0 kp.decodertop.data_received\[94\]
rlabel metal2 20286 14790 20286 14790 0 kp.decodertop.data_received\[95\]
rlabel metal2 53038 17051 53038 17051 0 kp.decodertop.data_received\[96\]
rlabel metal1 24610 20978 24610 20978 0 kp.decodertop.data_received\[97\]
rlabel viali 26173 25262 26173 25262 0 kp.decodertop.data_received\[98\]
rlabel metal1 53498 24072 53498 24072 0 kp.decodertop.data_received\[99\]
rlabel metal1 32430 17510 32430 17510 0 kp.decodertop.data_received\[9\]
rlabel metal1 23874 4794 23874 4794 0 kp.keypadtop.next_keycode\[0\]
rlabel metal1 24058 3706 24058 3706 0 kp.keypadtop.next_keycode\[1\]
rlabel metal1 27140 4182 27140 4182 0 kp.keypadtop.next_keycode\[2\]
rlabel metal1 26220 3434 26220 3434 0 kp.keypadtop.next_keycode\[3\]
rlabel metal2 28382 3230 28382 3230 0 kp.keypadtop.next_keycode\[4\]
rlabel metal1 28980 2618 28980 2618 0 kp.keypadtop.next_keycode\[5\]
rlabel metal1 30084 2550 30084 2550 0 kp.keypadtop.next_keycode\[6\]
rlabel metal2 32430 3230 32430 3230 0 kp.keypadtop.next_keycode\[7\]
rlabel metal1 31372 4522 31372 4522 0 kp.keypadtop.next_keyvalid
rlabel metal1 19412 2618 19412 2618 0 net1
rlabel metal1 58374 25806 58374 25806 0 net10
rlabel metal1 19780 13702 19780 13702 0 net100
rlabel metal1 28297 3434 28297 3434 0 net101
rlabel metal2 32890 5066 32890 5066 0 net102
rlabel metal1 35243 16150 35243 16150 0 net103
rlabel metal2 34270 17000 34270 17000 0 net104
rlabel metal1 20010 13838 20010 13838 0 net105
rlabel metal1 19589 23698 19589 23698 0 net106
rlabel metal1 15923 32810 15923 32810 0 net107
rlabel metal1 20838 20502 20838 20502 0 net108
rlabel metal2 28658 20570 28658 20570 0 net109
rlabel metal1 58374 21862 58374 21862 0 net11
rlabel metal1 31878 21896 31878 21896 0 net110
rlabel metal1 27929 35734 27929 35734 0 net111
rlabel metal1 33074 34680 33074 34680 0 net112
rlabel via2 19918 21981 19918 21981 0 net113
rlabel metal1 39015 15402 39015 15402 0 net114
rlabel metal1 43095 11798 43095 11798 0 net115
rlabel metal2 41538 9282 41538 9282 0 net116
rlabel metal2 53774 14688 53774 14688 0 net117
rlabel metal1 46736 12410 46736 12410 0 net118
rlabel metal2 39330 21250 39330 21250 0 net119
rlabel metal2 29762 36618 29762 36618 0 net12
rlabel metal2 42734 20298 42734 20298 0 net120
rlabel metal1 36708 21114 36708 21114 0 net121
rlabel metal2 56718 20366 56718 20366 0 net122
rlabel metal1 47617 25942 47617 25942 0 net123
rlabel metal1 47288 29478 47288 29478 0 net124
rlabel metal1 46506 12206 46506 12206 0 net125
rlabel metal1 47610 36754 47610 36754 0 net126
rlabel metal1 24748 36754 24748 36754 0 net127
rlabel metal1 34960 36754 34960 36754 0 net128
rlabel metal1 47288 36686 47288 36686 0 net129
rlabel metal1 58328 18258 58328 18258 0 net13
rlabel metal2 32246 36550 32246 36550 0 net130
rlabel metal1 40756 36754 40756 36754 0 net131
rlabel metal1 36800 36754 36800 36754 0 net132
rlabel metal1 29072 36754 29072 36754 0 net133
rlabel metal1 27876 36754 27876 36754 0 net134
rlabel metal2 25346 36550 25346 36550 0 net135
rlabel metal1 41400 36754 41400 36754 0 net136
rlabel metal1 38824 36754 38824 36754 0 net137
rlabel metal1 35328 36346 35328 36346 0 net138
rlabel metal1 38180 36754 38180 36754 0 net139
rlabel metal1 15134 19482 15134 19482 0 net14
rlabel metal1 42044 36754 42044 36754 0 net140
rlabel metal1 26910 36754 26910 36754 0 net141
rlabel metal2 42550 36550 42550 36550 0 net142
rlabel metal1 43976 36754 43976 36754 0 net143
rlabel metal1 44620 36754 44620 36754 0 net144
rlabel metal1 36156 36754 36156 36754 0 net145
rlabel metal1 40112 36754 40112 36754 0 net146
rlabel metal1 33028 36754 33028 36754 0 net147
rlabel metal1 34316 36754 34316 36754 0 net148
rlabel metal1 31740 36754 31740 36754 0 net149
rlabel metal2 58282 23868 58282 23868 0 net15
rlabel metal2 46230 36550 46230 36550 0 net150
rlabel metal2 37398 36550 37398 36550 0 net151
rlabel metal1 43332 36754 43332 36754 0 net152
rlabel metal1 33672 36754 33672 36754 0 net153
rlabel metal1 31096 36754 31096 36754 0 net154
rlabel metal1 30360 36754 30360 36754 0 net155
rlabel metal1 39468 36754 39468 36754 0 net156
rlabel metal1 29716 36754 29716 36754 0 net157
rlabel metal1 45264 36754 45264 36754 0 net158
rlabel metal1 25944 36754 25944 36754 0 net159
rlabel metal2 31694 36244 31694 36244 0 net16
rlabel metal1 45908 36754 45908 36754 0 net160
rlabel metal1 44942 3026 44942 3026 0 net161
rlabel metal1 41400 3026 41400 3026 0 net162
rlabel metal2 37306 2754 37306 2754 0 net163
rlabel metal1 42044 3026 42044 3026 0 net164
rlabel metal2 42458 2754 42458 2754 0 net165
rlabel metal1 44390 2992 44390 2992 0 net166
rlabel metal1 38180 3026 38180 3026 0 net167
rlabel metal1 36248 3026 36248 3026 0 net168
rlabel metal1 35098 2992 35098 2992 0 net169
rlabel metal2 57638 13430 57638 13430 0 net17
rlabel metal1 34408 3026 34408 3026 0 net170
rlabel metal2 43654 2754 43654 2754 0 net171
rlabel metal1 43332 3026 43332 3026 0 net172
rlabel metal1 38824 3026 38824 3026 0 net173
rlabel metal1 40756 3026 40756 3026 0 net174
rlabel metal1 36892 3026 36892 3026 0 net175
rlabel metal1 39468 3026 39468 3026 0 net176
rlabel metal1 40112 3026 40112 3026 0 net177
rlabel metal1 35328 3026 35328 3026 0 net178
rlabel metal1 34914 4658 34914 4658 0 net179
rlabel metal1 21712 2346 21712 2346 0 net18
rlabel metal2 15318 14212 15318 14212 0 net180
rlabel metal1 36524 5542 36524 5542 0 net181
rlabel metal1 36861 5270 36861 5270 0 net182
rlabel metal2 25530 30906 25530 30906 0 net183
rlabel metal1 56672 23698 56672 23698 0 net184
rlabel metal1 39330 10064 39330 10064 0 net185
rlabel metal1 57592 21522 57592 21522 0 net186
rlabel metal1 57546 19346 57546 19346 0 net187
rlabel metal1 57592 25874 57592 25874 0 net188
rlabel metal1 57546 18258 57546 18258 0 net189
rlabel metal1 22310 2448 22310 2448 0 net19
rlabel metal1 12650 14348 12650 14348 0 net190
rlabel metal2 23230 4352 23230 4352 0 net191
rlabel metal2 23598 35870 23598 35870 0 net192
rlabel metal1 22218 35088 22218 35088 0 net193
rlabel metal1 20424 7854 20424 7854 0 net194
rlabel metal1 23138 3502 23138 3502 0 net195
rlabel viali 24701 33490 24701 33490 0 net196
rlabel metal1 13340 11118 13340 11118 0 net197
rlabel metal2 25990 3706 25990 3706 0 net198
rlabel metal1 22402 33422 22402 33422 0 net199
rlabel metal2 30130 2516 30130 2516 0 net2
rlabel metal1 23506 2414 23506 2414 0 net20
rlabel metal1 23782 30702 23782 30702 0 net200
rlabel metal2 16882 13124 16882 13124 0 net201
rlabel metal1 20562 31314 20562 31314 0 net202
rlabel metal2 16698 4284 16698 4284 0 net203
rlabel metal1 23690 29614 23690 29614 0 net204
rlabel metal2 25346 3910 25346 3910 0 net205
rlabel metal2 16146 31484 16146 31484 0 net206
rlabel metal1 26726 7854 26726 7854 0 net207
rlabel metal1 32936 6766 32936 6766 0 net208
rlabel metal1 20056 12206 20056 12206 0 net209
rlabel metal1 22586 2346 22586 2346 0 net21
rlabel metal1 30314 7378 30314 7378 0 net210
rlabel metal1 26680 7378 26680 7378 0 net211
rlabel metal2 16330 32572 16330 32572 0 net212
rlabel metal1 34224 5338 34224 5338 0 net213
rlabel metal2 14122 6460 14122 6460 0 net214
rlabel metal1 28980 5678 28980 5678 0 net215
rlabel metal2 27922 5882 27922 5882 0 net216
rlabel metal2 31970 5440 31970 5440 0 net217
rlabel metal1 25024 31314 25024 31314 0 net218
rlabel metal1 26358 31858 26358 31858 0 net219
rlabel metal1 34546 18734 34546 18734 0 net22
rlabel metal1 16146 31450 16146 31450 0 net220
rlabel metal1 18124 31790 18124 31790 0 net221
rlabel viali 18728 31314 18728 31314 0 net222
rlabel metal1 18952 12886 18952 12886 0 net223
rlabel metal1 17434 12954 17434 12954 0 net224
rlabel metal2 26542 13056 26542 13056 0 net225
rlabel metal2 29394 24412 29394 24412 0 net226
rlabel metal1 26726 33898 26726 33898 0 net227
rlabel metal1 39146 20434 39146 20434 0 net228
rlabel metal1 20102 12614 20102 12614 0 net229
rlabel via1 36110 24157 36110 24157 0 net23
rlabel metal1 13340 15470 13340 15470 0 net230
rlabel metal2 18170 8330 18170 8330 0 net231
rlabel metal2 22494 8908 22494 8908 0 net232
rlabel metal1 48254 17170 48254 17170 0 net233
rlabel metal2 22034 11322 22034 11322 0 net234
rlabel metal1 26542 34544 26542 34544 0 net235
rlabel metal2 14122 11594 14122 11594 0 net236
rlabel metal1 45862 20910 45862 20910 0 net237
rlabel metal1 13156 7378 13156 7378 0 net238
rlabel metal2 14858 6086 14858 6086 0 net239
rlabel metal1 18446 20842 18446 20842 0 net24
rlabel metal1 53452 22610 53452 22610 0 net240
rlabel metal1 29532 21522 29532 21522 0 net241
rlabel metal2 16882 34748 16882 34748 0 net242
rlabel metal1 39928 13362 39928 13362 0 net243
rlabel metal1 16238 18734 16238 18734 0 net244
rlabel metal1 18630 5644 18630 5644 0 net245
rlabel metal1 22172 9554 22172 9554 0 net246
rlabel metal1 38732 19346 38732 19346 0 net247
rlabel metal1 51382 24174 51382 24174 0 net248
rlabel metal2 21298 34374 21298 34374 0 net249
rlabel metal1 18998 19414 18998 19414 0 net25
rlabel metal1 37030 7446 37030 7446 0 net250
rlabel metal2 38778 7548 38778 7548 0 net251
rlabel metal1 46460 24786 46460 24786 0 net252
rlabel metal1 19090 11050 19090 11050 0 net253
rlabel metal1 43240 12818 43240 12818 0 net254
rlabel metal1 30314 13294 30314 13294 0 net255
rlabel metal2 39606 18462 39606 18462 0 net256
rlabel metal1 51612 26962 51612 26962 0 net257
rlabel metal1 47380 26010 47380 26010 0 net258
rlabel metal1 13570 10642 13570 10642 0 net259
rlabel metal1 34730 17646 34730 17646 0 net26
rlabel metal1 13110 14586 13110 14586 0 net260
rlabel metal2 52854 25058 52854 25058 0 net261
rlabel metal2 24150 20638 24150 20638 0 net262
rlabel metal1 45218 19482 45218 19482 0 net263
rlabel metal2 31234 16252 31234 16252 0 net264
rlabel metal1 48070 20944 48070 20944 0 net265
rlabel metal1 29394 26350 29394 26350 0 net266
rlabel metal1 52118 21590 52118 21590 0 net267
rlabel metal1 47794 26962 47794 26962 0 net268
rlabel metal1 48300 22610 48300 22610 0 net269
rlabel metal2 38134 18326 38134 18326 0 net27
rlabel metal1 49450 13940 49450 13940 0 net270
rlabel metal1 47242 16014 47242 16014 0 net271
rlabel metal2 51382 21420 51382 21420 0 net272
rlabel metal1 38502 14994 38502 14994 0 net273
rlabel metal2 49910 28220 49910 28220 0 net274
rlabel metal1 49634 15470 49634 15470 0 net275
rlabel metal1 44850 16558 44850 16558 0 net276
rlabel metal1 51382 17170 51382 17170 0 net277
rlabel metal1 30958 15538 30958 15538 0 net278
rlabel metal1 48668 19346 48668 19346 0 net279
rlabel metal2 41078 18462 41078 18462 0 net28
rlabel metal1 41262 16558 41262 16558 0 net280
rlabel metal2 51566 18938 51566 18938 0 net281
rlabel metal1 23184 25806 23184 25806 0 net282
rlabel metal1 30314 20910 30314 20910 0 net283
rlabel metal1 54234 15470 54234 15470 0 net284
rlabel metal1 25714 26384 25714 26384 0 net285
rlabel metal1 45310 23154 45310 23154 0 net286
rlabel metal1 56534 25228 56534 25228 0 net287
rlabel metal1 53268 26350 53268 26350 0 net288
rlabel metal2 47610 14212 47610 14212 0 net289
rlabel metal1 49082 19380 49082 19380 0 net29
rlabel metal1 45540 18394 45540 18394 0 net290
rlabel metal1 32154 18190 32154 18190 0 net291
rlabel metal1 53544 18258 53544 18258 0 net292
rlabel metal2 22954 30906 22954 30906 0 net293
rlabel metal1 21436 2958 21436 2958 0 net294
rlabel metal1 29256 2278 29256 2278 0 net3
rlabel metal1 56626 20332 56626 20332 0 net30
rlabel metal1 39882 16694 39882 16694 0 net31
rlabel metal1 33212 12954 33212 12954 0 net32
rlabel metal2 36478 11356 36478 11356 0 net33
rlabel metal1 39238 23086 39238 23086 0 net34
rlabel metal1 19274 16150 19274 16150 0 net35
rlabel metal2 20470 22304 20470 22304 0 net36
rlabel metal2 20930 21794 20930 21794 0 net37
rlabel metal1 47058 23630 47058 23630 0 net38
rlabel metal2 53314 20026 53314 20026 0 net39
rlabel metal1 30498 2448 30498 2448 0 net4
rlabel metal1 33534 15062 33534 15062 0 net40
rlabel metal1 19274 15674 19274 15674 0 net41
rlabel metal2 19274 18054 19274 18054 0 net42
rlabel metal1 18998 21964 18998 21964 0 net43
rlabel metal1 24702 21998 24702 21998 0 net44
rlabel metal2 36846 14450 36846 14450 0 net45
rlabel metal1 32936 21658 32936 21658 0 net46
rlabel metal1 31832 24582 31832 24582 0 net47
rlabel metal1 36386 20434 36386 20434 0 net48
rlabel metal1 41170 16626 41170 16626 0 net49
rlabel metal1 30682 2618 30682 2618 0 net5
rlabel metal1 44850 16762 44850 16762 0 net50
rlabel metal2 39514 15368 39514 15368 0 net51
rlabel metal1 55982 17714 55982 17714 0 net52
rlabel metal1 56580 15538 56580 15538 0 net53
rlabel metal1 52900 21318 52900 21318 0 net54
rlabel metal2 55338 20808 55338 20808 0 net55
rlabel via2 39698 15147 39698 15147 0 net56
rlabel metal2 32982 29682 32982 29682 0 net57
rlabel metal2 33442 33796 33442 33796 0 net58
rlabel metal1 47334 28186 47334 28186 0 net59
rlabel metal1 1610 14280 1610 14280 0 net6
rlabel metal2 19642 16847 19642 16847 0 net60
rlabel metal1 26266 18632 26266 18632 0 net61
rlabel metal1 25162 21318 25162 21318 0 net62
rlabel metal1 20654 23766 20654 23766 0 net63
rlabel metal1 33350 21930 33350 21930 0 net64
rlabel metal1 36432 19754 36432 19754 0 net65
rlabel metal1 35834 20502 35834 20502 0 net66
rlabel metal1 37260 17306 37260 17306 0 net67
rlabel metal1 38548 16082 38548 16082 0 net68
rlabel metal1 43516 20434 43516 20434 0 net69
rlabel metal1 58374 19278 58374 19278 0 net7
rlabel metal1 54786 19720 54786 19720 0 net70
rlabel metal1 55660 15402 55660 15402 0 net71
rlabel metal2 47794 23494 47794 23494 0 net72
rlabel metal1 54740 21590 54740 21590 0 net73
rlabel metal1 56028 21318 56028 21318 0 net74
rlabel metal1 16514 18768 16514 18768 0 net75
rlabel via1 40344 12206 40344 12206 0 net76
rlabel viali 22114 18258 22114 18258 0 net77
rlabel viali 20104 18734 20104 18734 0 net78
rlabel metal1 20332 21522 20332 21522 0 net79
rlabel metal1 23138 35802 23138 35802 0 net8
rlabel metal1 23411 25262 23411 25262 0 net80
rlabel metal1 26910 13362 26910 13362 0 net81
rlabel metal1 36478 19686 36478 19686 0 net82
rlabel metal1 34132 21998 34132 21998 0 net83
rlabel metal2 35926 17068 35926 17068 0 net84
rlabel metal1 38272 16082 38272 16082 0 net85
rlabel metal1 44666 16048 44666 16048 0 net86
rlabel metal1 39284 17306 39284 17306 0 net87
rlabel viali 51200 19822 51200 19822 0 net88
rlabel via1 53776 19822 53776 19822 0 net89
rlabel metal2 24242 36754 24242 36754 0 net9
rlabel metal1 48070 21998 48070 21998 0 net90
rlabel metal1 52417 20910 52417 20910 0 net91
rlabel metal1 39744 17170 39744 17170 0 net92
rlabel metal1 27140 12070 27140 12070 0 net93
rlabel metal1 39376 12818 39376 12818 0 net94
rlabel metal1 20707 8466 20707 8466 0 net95
rlabel metal1 18269 9962 18269 9962 0 net96
rlabel metal1 18722 13335 18722 13335 0 net97
rlabel metal1 19304 14994 19304 14994 0 net98
rlabel metal1 18216 14042 18216 14042 0 net99
rlabel metal1 1334 14382 1334 14382 0 nrst
rlabel metal2 24886 34884 24886 34884 0 sending.cnt_20ms\[0\]
rlabel metal1 17986 31110 17986 31110 0 sending.cnt_20ms\[10\]
rlabel metal2 17250 31076 17250 31076 0 sending.cnt_20ms\[11\]
rlabel metal2 19826 30804 19826 30804 0 sending.cnt_20ms\[12\]
rlabel metal2 21482 31484 21482 31484 0 sending.cnt_20ms\[13\]
rlabel metal1 24426 31858 24426 31858 0 sending.cnt_20ms\[14\]
rlabel metal1 24656 31450 24656 31450 0 sending.cnt_20ms\[15\]
rlabel metal1 26128 31314 26128 31314 0 sending.cnt_20ms\[16\]
rlabel metal2 26358 31076 26358 31076 0 sending.cnt_20ms\[17\]
rlabel metal2 26818 34782 26818 34782 0 sending.cnt_20ms\[1\]
rlabel metal2 27094 34782 27094 34782 0 sending.cnt_20ms\[2\]
rlabel metal1 26910 33830 26910 33830 0 sending.cnt_20ms\[3\]
rlabel metal2 27186 33626 27186 33626 0 sending.cnt_20ms\[4\]
rlabel metal2 22586 33490 22586 33490 0 sending.cnt_20ms\[5\]
rlabel metal1 20240 34034 20240 34034 0 sending.cnt_20ms\[6\]
rlabel metal1 18814 32878 18814 32878 0 sending.cnt_20ms\[7\]
rlabel metal1 18354 32742 18354 32742 0 sending.cnt_20ms\[8\]
rlabel metal1 18032 32878 18032 32878 0 sending.cnt_20ms\[9\]
rlabel metal1 26956 28730 26956 28730 0 sending.cnt_500hz\[0\]
rlabel metal1 30406 31110 30406 31110 0 sending.cnt_500hz\[10\]
rlabel metal2 31326 32164 31326 32164 0 sending.cnt_500hz\[11\]
rlabel metal2 34454 34272 34454 34272 0 sending.cnt_500hz\[12\]
rlabel metal2 32154 34170 32154 34170 0 sending.cnt_500hz\[13\]
rlabel metal1 32798 33456 32798 33456 0 sending.cnt_500hz\[14\]
rlabel metal1 30176 28390 30176 28390 0 sending.cnt_500hz\[1\]
rlabel metal2 30498 29410 30498 29410 0 sending.cnt_500hz\[2\]
rlabel metal2 33166 28730 33166 28730 0 sending.cnt_500hz\[3\]
rlabel metal1 33764 31926 33764 31926 0 sending.cnt_500hz\[4\]
rlabel metal1 34086 31790 34086 31790 0 sending.cnt_500hz\[5\]
rlabel metal1 38778 30566 38778 30566 0 sending.cnt_500hz\[6\]
rlabel metal1 34500 31790 34500 31790 0 sending.cnt_500hz\[7\]
rlabel metal2 39054 33048 39054 33048 0 sending.cnt_500hz\[8\]
rlabel metal1 36570 32436 36570 32436 0 sending.cnt_500hz\[9\]
rlabel metal1 39882 29138 39882 29138 0 sending.currentState\[0\]
rlabel metal1 40465 28526 40465 28526 0 sending.currentState\[1\]
rlabel via1 40235 29138 40235 29138 0 sending.currentState\[2\]
rlabel metal1 43654 29580 43654 29580 0 sending.currentState\[3\]
rlabel metal1 44022 29104 44022 29104 0 sending.currentState\[4\]
rlabel metal1 44114 29172 44114 29172 0 sending.currentState\[5\]
rlabel metal2 31878 34612 31878 34612 0 sending.lcd_en
rlabel metal1 57500 23630 57500 23630 0 sending.lcd_rs
<< properties >>
string FIXED_BBOX 0 0 60000 40000
<< end >>
